��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�k�۸�m�i(b[�{�㇌�]�i�5'�`;Etg
<������H�W޵α���N-�`��6����ݾ�FF��eF4��_}<�ےA�[,�|{�?r+-��5K�z��!��[��S}Σ{$Gx^����c��ƀPfƆ���FD����q6�OQRryE����>��֚9ʾ�i�gL�'uj�⍍�Ϊ�ot��?�{��Ʀwa��M!`��ic;�Ϗ��Zeh� ��,c���|�u��P��4�5�ލ�"
FB�}�>�s�g7�Z�rبDt�����k�ۣ�Z���̵�J�"��Ϫ�m��Ѧ*q�f��ӭ�Q*h�oOTʟ�����D��xPt����Oj�yc��	��U��U����qB&	t�.��,�$e�4�d"��Y�+�6ڋq!��-�,�Ĝߓ�4���O�R�O��[y6�gN��fX�s�y;^ܷE<`��X��<�K�����vg�������Um}�J��9�H�N+$��=M��H:^Fp�8��Ou�;lAZ�FpM��_�q�-�H[tzL/&�B�	]�!�����XJ���#�d�#�S*Lڟ�|�!�H�jN��X/�W��K
��Ww�e�\"V��̒?�n�f#f�Z[o'�);�Հ��$���!V5���=U;�^1a5Zz��;N�>�|���ǋم@>F.�.�vnAY�_p]�jC�'D��� �&;`[��Q��;� �´��pMl��4��y�"��$	��})H^�]�`W���i�UfF(`n
���/�����0)]�K0�@صs�-TZ�[��y��� �bJVdAJ� ��A�u�uơQ�:Wgqҏ�O��MM��7.fp���y��;�|�&i<�'�^����$��TBc��[�L�$�(��&7�ռ˒g�<fA&Z�Mˠs䘊&���(���˃\װ���	xȉ(�aB{���w�=l貰�t9��tv�3{����9�Ww ����첏��=88xw1��Ӳ��h�b���;q��%���{Jh8�J|f
�7�.-�ր.ֻ��V��bM�5*T�$"��Bg�C�T �0B���-�_uk�|�bG��?Ug=��^N�g��Yb��}�u��ok��i���������6���P��P؜��F����א��8�������z�&�1����B%O٧�۰����nZ�=�:�����$����rC.�("�B�p�"t�G`�s�-�ll�p�������N��H���b_-�w����h}�	�0�t��F!��_sܪ���hj�h��/��z���\E�'�?��wz[�T�7�5� 9X�]x-�Y:�bP�5b�=�q�#}�+�Wß_�)���������K�:�[��/��3o��q4���ӓ?�|KyX�b��r�ܽҴo<ئ���g(�v:�����km�����������ڦl	/vo����'qƩxu%�K��'��*Qex
��)ǧ#�l#Im� �9q6���9��!T�uI���3zW�s�NK�^pl'��p{����o�|Т������2
�BO�ﴚHp@w���@2,�f��{��|�� �_k����;Q=a�jq"ۥUa�
��*N��+W�ok����d�1-�>-r%���"�F/�z��#����C�2a*a���bh�^V�*�ٰ`;���+��J�,B�����- ��cL�	�-Y�U:�s�s��lf� ��x�TJ#���[�^#~����c����k"�/�$�Pk3o��;�h&�+��Մ�T�Y j��p[�����> G��k�v�d��.�[�Q�0�O�
��z�:mN�P;(w������=hP����߭�	�\5����HXe�U����)�N�Ŷ��ܓSpj�g��I��/T[O9�a���-���P�q��zV(�8��р�:�����&�k��b�/`���Y/1%�!'�x��=]�ǌ�8E(\�w0�:g��9 ��^�^c#Ѹ�����af��mΩMCu[{�<� z�Z��	3u�t?�s�'����Y��؞Э�E��L4̿E���0�ޔ?��;S�x���;�9�JI=|�05 PA�A���Z�Ц7��n�RzX�@΀��4?�Z�B�*�����o2¹��4#e�	c��@�!C����=�����fX~A3S�P��7�B��{c�@_0oWu���t��\��y��Eu5�6ɿ��(1Ka)`k�y��g9rnMe�I3�o�R��gP�*�Qf������ٙ{�]�7��o�Z
	�]:�.t
/)@�U���aBr��)� ӀWbj?-.!0v�o��Ǖ��*�p�Z-μ��*^���V�`P<�%|�.a��D�>���Ҷ�p��v��]�!���7J��
�d�g�K�azQ�б��4
;*Z^�k�����'�P|5���Q� ��=(��8G���$�:�ۜ��JYC��y_������.<�p�9��&�K-��!���u	}�GZ���������g���o���l��~av�/��b^��i(i��I��>���nl�A�����$[4��,�o�TY2�=����_�F�ҟ[���.@z�1����I�Ex����Q�-�Ё�l0V�;�މ���G9�{��^�L��!ߟEQ��H�?�{R��PT�侌a�E�!?��r͊7���g l?=�f��J�� �U]�ZŌ�x�3�%���@~��s�� Q���T�(S��"B���xTHv�4���������Rk�]��L��=����o�E,�3�|7إWU7Npa[u�Xl�YO#1�'�e��"��o��~7�肊�>��W�F�X#"��#R�M_ ��h_��#�}�8�l�#"����꘍M�O��{�A�\��g3X�(����2��p>Vmg�0��v�*��p?2O�ب�e���n��)<#.���b1�c��:΢�LE0�z��yY6��e���(v�uu0HQ+�-���v�C=�