��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jåا{�\�u�?߷�dn@6�zf��r������;$VF�w��>�h�hB��4jJ:ѧ����}��;�À����8�ݣ��,l o���Tl�)Ї1�����eyJ$��o�pj���be/���a�!�7�u�O�����b���7/��B"h^0 ��x�\��<!�.��N~�|?z�>n�u�$�1.�_�лOY�R�����+/�l���e����c�ti��Y��2�w�:�)Ύ&H/(:��*��l��<D��~���r3���CK�-�'Z�c��D�,N�w�F����~q�\b�O�.~��*=����Kϣ'��x
��g.9�ZԈ�Bs���yD��߈�s���|->!��d�h_v�wRY���7۱-�g��b;����I��z��φ~@����a�q\IΞ��t��Q�J���v�<�,�PE����([��}i��WQ��D"�R�?#|�I�����G�Z�"��f�.�p��B��7��V��i6A��_�Зs��A$�@��L���`�ߜ��c�Q��I4�򪓞�$��Y��Q?�vޯ �o�3͏dN##0�_�ܪ>��q�� ߠl�jf�%�W�� ��0"��}(��+���>��iI�{�$�6&{0� � 5k�ÆU&5�q���y�lh%KA2Fb(���F)���A�D2����k�V���JZ��!2�P��]ӊm�BwԥZ5j�9�Q72��o��?��*�X.e����F��#��G��}oq�f:=P�,2smɯ�^D�B�ŀ�'JR����Y��&�'_:�Pu# x�-��WM��ĩ� �?S}�՞Gb&h���1�nA���lM6�!4�Y���P�A�������kZ�n�P�p�Ȯ;d%fl�������5}T��K�s]l�)���Y;���U+/��i6 cH�0�����M��gJ���îW*8���s�sf��>����_V��ӣ�r@�l�,͘�A�q��t���,ZԷlZ	�|�y��|(��I��3/�溭�a�B���r������?���cQn`�G����	��`��De���g�o5ؘ��T��	ݭԮ�GI���s�۟P�9K���i��pYR�@�J���v�&Gc9�$#r3�e�85���d�3��1a�/MaNs�1�K�,�+`�
�O�� yK-�\;I���X�M�V�?St��o��A�G�s��?�uN|�t�A�/W�js�Is��c�`a�0�1��(f.^����q�(D�K�ӹ�۞\���h�Ei⺕����bkr������`o����� p �?���`��kʱ�v�ʕ^K��n>��N=Ξ�r���eH{�D��#�j�y�����b�Ð��$V��\�3{�Xv~����.AU)�g&��KWt�r6�J5̈$7�o�1E���A�V14�@�z�橂����с�	+���i���9�9.+��@�uZm�?qBk-$�ݶ��X��5�ݟ�NORA�WE-E^��ȸ�Kry�U�p�;��^�l:����0d&�S�'�&;����D�JR���Q�>v������#,;��][7��|��)�