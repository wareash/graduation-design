��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jåا{�\�u�?߷�dn@6�zf��r������;��[����t�K,�h[���B���zT)[-�j���u�_�/��x����	����c3������8,�6�|M���\��v|s1�&%�DPd�u�>���ꆈ�˿�(���G5D�v\͑Sƕ2����d����J�R���c��8 m��gFR��a9s��RH�NI���a��x���X2�g�F<r�}-~+`6�U��d*0����i�&0��d˛�nt��>�ive)Y��e�ҊK(i��%#:�L��t�<W+;7Oem%Y'i��k�����+�R�{�����F�P)<��`��)�p}_�	��9�t�Xvl�~Ԗ�p��_�>�5�Z���S�5D�0�x�-��G�'�A���a	]pR��=d�uPK"�#yxɢ�Qy�%y�FA5�K)����in8툫+�ejܤ��Pb�}WQ�L�f�s�)j�[���/���z���u��Hi$B�7�Z������:�4�!r���r /#��$Ge�O�$1P�d?"R��?�Q
Nd��Z�B���$"#^޻m#����4-e٧/���k/�K{��&�����.{	��?,Nl�(��\�4߄����>�xrHJRI��aՆ��t�����'��
@ܞ�	�k�@h1E�qߧ	lRI���V�����){A����P�f�-~�qX�b=�Q�;�$��_�,v�c�R&�����ח�״�X[�ӝx[�[���v鎚k��~�=�莙��;@���٣U#m�?���	��'�j�L8˼�sԣ��Ju��fJ���>_/�����gM���)�^�^��8��W�Rb��V�6WPw۔��Qr�qN�!6���2�b�S��f�W*)��),�K�$��-��jE���͚ͺ��2�/o�r%�O�sM�ՙwB�l�?Ǌ|�N�Y�ld�}@�q��Z,}�����-����\Q� �=�H��<�U9��9�iҷ	�ao�9eE�~c�^ݭ;�����m{����'�w�\�3���z���4�������ڌ:�4<l.�:l�_�Mܼ�c5�Ώ�L���	���^^�!֋�}���TM3������;UZ��}��Ϟ�WG͏kw u0����k�P?�ɟb9N�Bq>�5S3�����kC��	�"���p���¨�>b�·�
~�X�QG�Ԧ��Ɲ7us&�{P��|��I�V�xu���a�1��'�Q���kP2\.�-�-8�8�lXA7��t���ш6���2� !�p��>���te��3]���=�E����w��f�<���ʀؽR��3�GT ����
d�\�Bio�`�T^bONP�"Sʩ�}o�_N�z�O-���ƥx�vn�Y��ˑ��\x����v^'����M� z�A�T�'���1�0�7 *V�;~�{Uq���`Σf�DT������g�3���k���ttuS��ll��"���1Q��6����!1�e�<���E\�V������W���2�l���E���r���Cs_�\�"!�h��#"W����1Mֹ��^�} ������Nu��ɡ�ӭ%#�$D*��n�˒�����Q���I�D��^.��*���P�ᘤ���Uvb���%����(�(6���4���I��z[D*6"N̬���t~�.��u�׮�pK�S��U7E,K(����4%x��
"�P�6M�o�z��|���߾v-�%>0�St�����t�C07������&�����-��̦�}?}X.B#�P�������!�/�S����y"��z�DT~S-�ij]�G�a/�!���5���6B`<��҄1���Z�uWd
)�0�[��)B��[����MP+��@�?V�ޗ�p��
#"��E�<�T#p���dw�~�F����^Խ�Yk��F��m�q%@ͬΐCvN�ni��y��D��(�qݣr���)����q�=/���?�W�:����@q�g��x ��<  , :2�$���C����ԋ
G- 1>5��z7;����`�AsŴ��R�M]�C��ʰ0�5���񠉀TϪ��Xb�qlQ�y���0�8 ��E�v��TD,ܠ(\����)�	�%��"K:^��	��e�Ԓ�<C��Q����n�׻�1���s*�g���Ht�v�����a��C��tJ�?~ZӪTr@!Gc�h*(��S1�?�� ���:�)�ga�\?�mO�_���"��ENxp}���_��H������*݋��v=�m��L\�3��\�7�C�(u���'�C�ʽ��fT�gk�)����}H?70-Z�W��$����M���lI3)��n�
�����;���(N�D���S����;�#s���3�����5Zz�Z}V챨��t�ٰC�n~�@6�Jo��l%=F{6��Ґ��	���.+F�7�댂T���V�ĥ����#��mٟ��7��j���g^��P��/���n���i��o �A�Ҧ�Fշ��@E��E�4��B��҃+9k�l"�p��qB(��i��Y�{\ja�G��x���@�f��x����-7Q�RD`r�z��~G�_R���Ze\`\~���+@.��6p.�D�=�,�_��� o���*�Cۂ�(�ဖ}���H���:Q)p
k�eϯ[Ki���'�F^�l�hmG�r}^1�V~_9U����:/
6o��������Ҏx�=g�+h����gB�Xb��BQ��kN��ah@Ld�7��2�\f�.��uA�5��f�e�U��?��ݩ^���3y�c�؃����K���u�{L�߰�.��P�?�"���x�" N��)��689���;?Զu+�-wRC��O/�aQ�������հ��v�I��Q#�6df_4��܊���o�f��/�*�`b���;Za�ei��r�w���w�X�)�=�G�h�ݫ0� MØ�F��u��j"��"�e)g�S�v
?������f���� l��%D���O��f�i
4�����oqo�`Q�H���U��]��z,��@/�y|��xZ������g?IbT�UJh.������^�䱔,��Xv8��9u7�pj��r<�1�*����ܪZ��N������7����;����2�K�OJݩ���=�`��c�aAH�l\&��'?�/\F�u�Vue��u��"?�\o|����)$"Y!j$Q��G�O���@A2:'�֩�u��!p��ŁQ�^;*�k���I.M/2ϳs�9�u(�j���hT��筐F+�ҥd�E�V��.���vY�h;���RF �ptŀ#Ej~�E��$lC�N=�S����d��wP����]��⚾��\`̂���fKձ�������w��˂����.B �i�B i�9�����Y+]4�Ŀ�#1�⛕�P;��˷D���~*�wKy��&���P�%%�i�u������z�w�]Uy�oR��]G��h��ޒ�E��Of�o7�=�
x˅�۹f�:#W=ޓ�w�j��Ě�+a^g��wA��P$���n��޶�Sdb^D�MA�����E��H�xm,�V<g��&��#"�z���yT���z9�jJ��/��3��f1�g C��W�Q�F*��3�x����0p�r�Mi�������aP���7QOը��@/"�����5�7LƂVC<>�x ���9\1�x�@�cf�X��o�?*�.�4�+u%�0��`�y���4�qXG)�)QL��abH�����0\c�&}��?��/&��Q��<u�%Z�y0����ܴ�(�$�E��g�2�R}��0���sAbffY�H�upI8O�.UZ:�����9I>�Yy�	�*E���gؠ��Ra�>�UO���z�_U\�l�z�(m��E��Z0�fE����@O/:1w	�+�9�����iC��>��;\|fh�w���4]nN@d��b�xF����]��;�������ԧs-q9m�Rc�K�d��lH�bL���^�a�?[���z�Ha�GĿ����S�o�����fx30�����cǶ�_C�^1<E3���;f�_�)�e t���E���Q����@���-����"��
^%8��e��?״�h�w��n��w�@��O�Z5v���ڡ!4t/���Ě���F�
��2�6��t�����ug���+�h��=a���!nF8؏�]�s�iH�3S�ߛS��BV��0�2f&���sS�C?Hm�7f��i�&(�Uem��ƴ��i����Q�8���!z:#��_��[���b(�\�f�>�4��-�sŃ�S��6��)���/>���CA.R�x�4vq�r��h��ݚ%`-�FΥ�~.S�o�O���9j�ӎ��3��G����������:I>��L�|�'Ø�7R0��["����V��X�!n��g_O�B�.j? �k�f���̅V��"ծ�� @T����u��뱤�j,�#/����Nm���EXxՀ�f)0�%���v���Lڶ�bI7;p�*qI6�TQ����^��s)~��� O�L}���+�F;��@yCĳ��j8�q���vz�n~��CSQŬB��p�27�n4��t`��$"�]a����n"�2P��+�nI[5�.E���8�E,�釬6)�,�9�E%��O�v��,H�
��A�,��Ahx�$a�7>�5�ܼ����"5��BM_�N횖o�N%�|�h�x<=p��œc�M����pH�� �2wO�X�% �)�B1}�0��[��W�g���sб7���CL�R�޼�����ωV�ʋ~���x�7�W��s��La��v7?��eV����T)���jXn�~�Usx���Pq�y�=�����͸Nd��|l�C�I�^Z��&C]y=S�5 4���l�� ��������,�ٹZ�#��{ty��Hؠ�O�i`
a��p�0t,��~�zZ&�`���ZJ����[WB}0P[D�,��`��6�DƤII�Z�x�!����м<��]��@ξ	�0`݆﫽b�9���S���4���'�?LVJB�#���)̷p	!��?M�O+��n�;���-�����k� <�i�Mr&�#�uO��w�3��X]c�x%��WX���ż��5P��
�-����a���f���
�M2)e_zh{��H��-s� Qd-U楖���6��`H��50�*h����.L�2��OƝ��p&d�������螩��,�rBoD@��G�bg�Uŕ�W%hKR�]\�FV���4���b{�~�C62�M�2*�f5Nb����XD��`
�o����&��<�qx�B�cerb~��'i/X_��+���@�`�F���Rn|&�=g.�fr�N��T���d���h{���"�F��5[��j���G���fK��K|]����<ky�R�Ũ#�+Ʀ$��.Un˟Hg5=�tS1�	��WZ��X'�<�#���t��[�����=B҂��⿓�1�������F�k*��6��;Uܽ>��~@�s7�\���>��@B�wTѤo6�>]�ޯ)n	vq����Cj�\P|�y�-gZ�%���LP�b�z��"B{�����ȡ��K�̪D������t�a��	0���)"N��V�h��a��c���[{	�J<�r"w\a��J����0��2 -R�fW��W鞖�g8�Oʟ:�)d��zc��R@���LA��.����I��{ �|�B�Z?��D����&҃�8��=�/�0�_��r�uޡt�0��f���R$�Ʉ
��"���ZKȺ:���q!�of��8�X�
�2����R]vD�JD)H�k�s��`寸�E�] ӳ�����r/���^wy6uּ%
d�9�$�OA�b��+�qy���2�L�c�r
Q��$�<&u/�l�F�׷��gu���ǆ��H���{�"Pk�N
�tL �[��XX<��G��3�����/#�ǖT-�I��~5�|N/B�ɁCB�m�3�G.�n<n�j�K	�������>2�*渎o���d���p}�J��D�9��~�y0#=�;�p
l�\VrDSJ�i�]N��0��VY�~2�UYk���{��<ބ�M��;���
�ؑ����x�\�� Y^宝�pL�~�K�W5P]"K�؟��I����OU.�4�˝��A��8Z�I$L�gL«�Uu(�՘�J	w�{@��n��6��M�}	�$��ۨ�Ex�{�aF���&|� �5��~w���w."�E6V:O%��/.��fOq�L5���+�3> �ç�
f[lz�J��S��d޹}")1�2�aּ;��[d�R6r�tJ.fKLe1.Z���n�a������@H��_q~!A�W�w	�g�jgqhg �M��/����O�c�e�>���ȩ⑹0=�Y���5��������=�p�ǕV�^k�g�EQ�2�Bo��'0C�`��@���t4¸`�#ԋ�N�=�Le:J�HD��TG��-�+ܻ0'�A0Np�A�u���SgAȕ�'��W���X�cR��V�
{rQfY&�ָt	 _��b}��eCT�������#-u>�Q�J����ڢ�h���U��Ӧr^��;�������]N�;B�������@u��u_�|�G�t� gsfjvD>I�����|\uHN�p�lNN���������K�*�^�l���H]�!���4���w���'�� �$j�x�C���!~�l����� �֯�/�������UL���� AO�BoH^��&�ޡ��`�Zs9��Ua������O����(��ͥ�93j�4~K��ʄ�a�ª-K��ϗ�.�ԇ/��"[� oð���[U
7�u�(Y��?x����c� PT垭	V}��`n#L� ���t��lə�H�ɂ&f�ϫa&��+�_���XK�.��`�^��'vR�����B������<��<웹�ډ$wB,�L��X8-�Y8�1{$��ˬi0Ut%�Rz�X~��-�c����~�|J���K�%~���{7P��pW�S@���9�L�+�&�V%��ޒ��K"l?�I�e��h/:�{�9����=F�����|<�,�D�q�Y�L��|���N���d�vY��t����u>�p����%�Gt����*t ���-��B�t�5������%y��@S��?��d�~� 75��!M��2�����>�:�AF��~�^i���
���~��{�`ĺ�s �t8��j?[���X�M�y�L�ʺ#A�Y�{��J��+�nE�|?��� > ^��Nd*�;9FOk�-�g�@���9��C	�"�N��y3��]MD�X����P��c�1VMbgQ�9�B��#���t�����7�iݼ!�XQ'�p)�5�4��=?> ��#D{ �CQ�S�7�/����_��E6^*�`*�,J�����K� Qt%,�M*�m������g �>����PY5�H�~.��o8�������9�9<��I�K���ͱleM��Y"��q�pSIN;ozH�KǱ�!�˽�t�X���'�9�8uwd���~�9��y�>M���D�=�,;�i���2i�@q.��tw|�Jvu�m��j��3��D��^
���MufY��U䆑�8�%���]&ܟ+80l��LN���%y�Ӽ���П�7h�6�#D^��>�� %�oi��sEN�s � 7�p8QOH���R(�g >��=H�F%��ѼvU�T`��n>9�P�N-���l��Zp�"l��%qtw��D��zy{,�$�M���`����qCɩ�+p�z���,��~;t��iP+kR�$��J]c���N�4�y���M:�ۤ�q���#��d3L��l�l���4��<q:+���!�u]��6q]}�j��q%퓼e��8�����?���=eޏ�W��p[��mΧx�/��e�0;�$q�p^�Ú��&�GS c����x[��t�ñ5�5�����B��|}u���De���z��x��G�0�t�ov{��MQ)a�����``�'ᝨ7Y�e��$vNkrW�TE*�it�<0��`����WӀ�