��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jåا{�\�u�?߷�dn@6�zf��r������;,��o+�[���1��,)gO��J��&�fx��ė���}'�w�g3�Gv>��C��5�U�+P��m<
��1V6w30ԗhMc!�ԢFq0�́�o95��kӁ���=���v�%��h��Y��]30ycIy�7��wK���(�U�_�`9�"u�B����@�<�c@97w����K๷���z+:�!x'ei���a���[����dR9f����%��Wt�(�Q���h�_�y6!Ѕ:��]u��$\snA}	�ufk=,Z��(�u�iF"�� @HNy(*�?[���C/˺�8�Ml�M���t�u����:�jhP紟�@�..]��Eѕ5����H�"�N�x���Z.����=Ago��&{
M�1�\o��tm�_�3�qA7/v��p<?�1
y�<k�S�"��VQ�ք��RCK`�s��� +��_�c�n�]d�M�U���HVLz�a�<8�#5,�w8�;�{�c��Qu([��$g�$P�<�" �2�}���vh���q��ӫ��������nɘb��^R���/t/�M/�]d�.N��J@=��5]�-�`��8��mq�@������r�������R�
�}p˭�HEn'sX��i�N��׻@XjK�=�J�RX�b��,L����2u[b �n���1VI{ٿx��_A��bE�8�T�+��2#�	�i��&HgĩׯA�\�V�����65�LE4�,#Dn<x�'�B�y�hw������ 5�RK��?��t8Ɛ3�fe-�$�Mӷ$~�o��#�%{'���4�]-��֭�6@�5"��tR��Z�yҞ �96��E��+/&y�Ct|�2�#�kpE݄V](kި�Xh�}e�?|7V?ee.� ܡ*:�x��y���M���A������G�N�Ɍ�%�9��7�ԳZ'���I5�Hh�hG�`���5��72&�����Z�5�:L}jb�K����q@8��^w�+�W�*�%](⫸�|a��l(���[��d9/>��Q��9<A��%���<� ^�lAZ�/�l�r�eXn�#�xLypr;'�iɫb:Y�0ܶ�޶��_{�(#P�u�e��<�k��h�WI�s8gT�K��%!����-�V���>
���ު��'���z;��;#WkzB�"�yǣ�a�|A����/��_�Ad�[��j3⌒)�@:���i�ۃ���+I)T#�z9V�t�a��sm���0� ��پw��?���-�_�Ĳ��Ȝ���e��4��/ZJl=��x�+	�Z���I�4|4O��9�'u���G_�ac�������]�B��j�D��?G��.��q5�R�'���<�з?�ej.N�~���x��1�A�6�"+��>2*�v辛�,� V׉)�=&�a?�m��.��봯��I\y���G}%?� �1U����F��Cy%�xܹD�Ѐ�N���{����a��$5��6�i���2�JԊǪ<;SRI�����=��������w<���hOUȫ�)��e���$Bo�n8��[����P#{�u���qQ$�g^� H9���+}��o��o��^v��M�$�q��Te�Q(^�[�st_ī�'�y*��5nj<*��r)Ҿ.p+~�u�9�f�#󓡉�3�[ݫ��\̃��&Hq]�S�/��Qp*L�r��\���2�G.lE��b��
s�i�Jv,������~b���[��~Vr�.��ު;u�W$IzfH�vL�e�o�Q�{8)��*Fbfj"a?8u���a�'c~:�E�����P�P�̒Y���w~�l���|���70��-�4u8�ʉ�*��CV�w��`���= @*`v�b���F\�y��&�s�'���(�t4���|�&����'B�ǂ�xQop3oc���.�y��"i����a��5��y�5���9NBo�(�c�/�耑��9=#���講��MIa�_������L�)�*H%9���������
����5
�y�s���5��Jj������2W�ħ!����1�Qbv��4����.���X��=�ͤ��(�>-����X��)c��HR�3MW�e���u�Rl5L�(�&~�܆����F65�!�ovz�F�����$��&���_��;M�h}�����Ɓn��LEPRU{
�X���ʳ5��+��r2M�y����4N^Z�}�xG�^I� &�*��4w��:��}��AP���w�!��_�n�ˁp����z��;�@?�8,�٥��rP�A�}M�U��Yں���)1��7��ϰJw�0^���:�������pN���&2�,B��Q�@��C)�BJ�y}�G1tO���w��Q2�	�̰�^�]�g i�%4�k>�8���ꁛ��!nTM�uN�ʩ'�#'&&�#�;��D��I^���`3BO~�ÅP&��"����� 0 ��y������qlpB�flC�i*g�y�[�����������	�&�1��cy���%�7�3�`�Ua��ٯ�>���f���>>j�S�bBn��&�*��s�xw�l햅���t0y^x�,O���.`[ƙ��R	���%�fmǇ'ĥ���}=����������;�A�)��Pl���m�
�c�`�P�%�	�t��e��K�A�}Px�o�5 ����G\�#�D���KE{�|�!5y�ߔ�!V��R��~u

&�*1��1c�eT4G�=�a�'�7]����.� X?�w��@��S�/-*('��=<�0�BŗJ;���C��l�--TI���J��/�g�X"?WJL��&�q4�Y��j�K|�s�����#�t:��qE���:���,Ǝq+}1�At;�MP
h�"=��a����}���������N��+��Gy\�w<��'DvEE������g%���r�#H��Č�������(�*w#���Hḯ�#��h�.�[+M/�E���`\���df6���~����w|b�;���.������M�
1�Y�Vx��s9�m�O@k�ӷ&��vӀ�ܽ��aW�׎��֫�"�+bLRt5���6B�;3�.k4PF�9�|ज़��.ڹ�2!��z� �;gQN�WaM��ߞv�F])˜�ڨ ;�!b�RS~��I%���4�!�ut���e>��=�����Ӡ/�zL�J�A}$εܕ+��
�"IR�
-�������2���zR���LA��-bV/��'3��'�2�=S����fh�&]Xd�kYHT^�!4��<c=�j��x$��_��4!���mO�:��j��U�@�� 
���Za��:�{��?��Z�Z���$[~foL,�鰍)���?eҤ�B��*rQKq�ᕿ��h� <������	����,��� ��N����K��
U��e��۩�Zj,X�Zz���L�6�������/m3W���p�x�?D5^�..��Eͅ���n���L�R���6�A�Y��c��2�Ur̺�q�Vre���9�����p����]
7u�ڪ �O5<��]`{��)x�V^���f��H�9�+��*����o{�� ](�vW��>�mη�&C������:���C\��X���\�������`_F~Y� �E��1ר�pј��i�uW���M�Ù������v�@qg��~�n#!F��_~�
I��!�~4F;F�jr�a����u�`}e��D
hc�;B��h�q��'���)R���l!�u�3y���FzNa �Wơ�
	�V��#k�:{�I������9��d)�Z�*�����Z����y?�=�i�ň�3�E� k���n�G��UA����W6�uB�K7m���e�X�a���^Pd^�B)?��g��l^y�[�Z^3�p�?�2슺i�Ѣ������Y��`!#l8�&�E[|����SF�r���<j��Um����{Y�*�X�rW36+��}^3�xw3���ƛU;���~;��5V�z���	��y&L_��J���L#Q��B����e�]S�$�gG���у`�Zc[B��
��X�P&�z�M"�$���&�]!��l�icD��`m�PJ���[q�����\J�}�w[�|h'����dB �� (ės�p�N=���~�1j�1PAaʡ��(������ܟB٫J�"}��va��U��.��8�͍�����?�Gz>0�@��,��ApfO���cY{Co*��sʁ;��J!Y��r@!��HP���e,��^�8��{4��o�
���_)���B{�̪:]�� ��0N�����w��/��J��������]L�9�fλ�AB�t�]d�h��p��c��}p���D��F�¦��ɉ� �7)�;𔂼�R�
g=X�۠�L�4J<;�銹�{���V����C�l֮\�y/�d=�7%�bx^�5�Wj�@F}����4��`!X���aN�<� ���Ȉf~	�K���B�I
�F+��E$��;@�����`?�1� ΐi�(�6p���~���0�h�����?�\Z�KEI���ST�����1T�9o����KB��e��u,��3S��2���i0v'b��*����,���N����_��g������J�*͟����5Y���;fg�ޗ�,dh���u�X���w

��CzyV*�`�%U@ۖ�Q������;���P���9�Â�����4%������/(Ф^<���_�K�ѹ2��P���A\�S�E����٧iJp%q˯9�,�-q_�p
�m~�m��P��kg(���YR&�;�|sY��4�k_W1'uCH�X������l� �@��0s¾�6�'Ր�.g������W�]�m@�v3�6��(H�IMU"�E�v�wC�N�;�R����n���rZ�u�h��c�;ӝܱUm�Ķ��4���Ѐ�k1�`�Ω.Q�\H�p1�`�p�3�4ػ���nbE�|%	q���v9㐌"�P���8��6
�v"l]ǰ���X%<s�9p�Kue_�"��+[�#���(ְ͙�����3��N�Y��&RC��o��7=�^��O�/�����fVb�g?��_����3@{�<�������u1���-��Xm}`� �~�P�-$��pU�A2'�O��cu>�������$��G��c,C�g;ڏ2T�e�"������N�m��<}Ԅ	��b]��:NN6.�4�!5��.Fy�;l��gn���^>]�������W-4��t�%�!tp?E�J�c�����@7�(�L/)="z�n�H��Ů����V*#tB�P�J2���B��[��+�0�\��ɿT��k�嵰��miQ�5�i���;���.�s��/�B�T�,�
�-S�Xh9
n҄~�Y���<Rڛ3R�Jڥ+#�w�A�5.Qy���J_9���(#m+B����`k�a�p�A��7`�g�z�/���S��8ۇg����	�{o�ݖN1T�Az�8Ј��t\*ܼ+%kd��HA
��@/V3���]ᓆ}�"BQ����?*���d2���~s�G����А��"Y��|'?�X�bu��\ܫ�Wx]U��f3M<N
8�j��_�nT�X��fj��L3洃e8]�>���*�yt�e~�b�*�ϕ������=�5 ?�����0v<��L��Q798���	�*�΁��C�zx��I&�)�{'�3w�� Ѐ�5a�>��k6/�����jWB�١�O�M�q�?�u�>ފ!���������۸�-���A�^�%��	?� x��2�A�m�{�>UL䖞C�8J�n��Hj�;��C�2}!MK�oup��-BKdb��_�JO���؝Bz����}�c��=�%H��$��8���Aui������^zP���$�	Aa�r-���kBgiM	��a�ǎ��	�x�e��B�A��O�� ���>���y�P�>3��-�Z@*�8O3���6�>	�f�Q��ƈ��a5+�Y��0I9f;�L�V�T�~�)������[X��Q�����@Kv�Ne��|��8!igR�a˜���s͑ ��;��w8n���q5����Z�f���C��{�N�m�STA�����'wQȅ�uf�|f��xMƙ5�ᘦ>�!�ߡބx�΄� qy$�0r�̀1���H%���nɶ>>�t6L��6��Ĕ��~����Z�=�����Z��N�k��y�.֒7�k�k���rH�.���fS�*\W9�3q;�O�����Y�}BjG��nֹ�Y�����ʑ�R�v{�?_�r\:�EP��|���l*z�6"�e͑q��1��ߺ9��g���p}š�5u�ҕ��;Đ�7q��R�Yِn8HQ`dØ�n��QrW�U��z� ���nUq���>�n]ܚ)�`?Y�����^E�f�����LQ;c��8�A-�Lb��J n��|D�
��ƭ)��-��E�2�� �B90_m��r�]��_�_�J'j���rD�͎�}M�{%�s�a��T�n���� pw���m�sS�3	'A{�wi�};��x:��-����Q��2=��<J27v���6�׎�z�����_;rZev���k��f�y����y��Z/��3.�_O������mB��A�x����H��Z�K��9���r+M�)s���c�2\�|��CY��{q1Q�g]� �Ķ���ݵ��apXj}���߷dB��%o���*AH.���I��;��K>�-_{0�aa���Q�$�{����.�Ϋ%�N�\p���!sx����"���k�����F������-&�q�����#{6eu���j�9 N�u�v��l���C�(��`�B&o�T9��7#��z�ߣ��9�Gy��~5�^X�b�FN� XL�����
F�녆�>ǝʂy�4�����d>%�yP'�����x�E�8�h���6i��,�'�����9���/�2�y�u�����+�Q�����[���	c���X�8�G
.Z4b! �d.�F#�G�@��i����#p��{d�9԰��eu�ݏ�?	wv����W�,�f<���|0�]��ę��hM�N������|Y��3s��:����~��xR�-k]%��D���rg��L΄��A�D��H�"��d�>k�U�_�|AvذCn�x&���l��؀����>����v��JZ�٦�;<��?y�W�*�����jI��H�������r���,R]]Qk~i��5�F�wZG�e������#�ԉ5{�:u·��r-=�J����srl���~>�lC�� E�8��wg?���&�AsP[��#T����[�B\ND�ͼ��x�}Z�?:��CS�''��ozU����z����a���ϝ�:5���7���P ��a��.� @�<��F6
����bn����s[���g��O�j���G�*N�����-_-㣨l���3�u5H�Q >�K�,��8���j,�E�D�Z�H2�N;���AeyJ����rV�\�4���w��[�S "������<�l�4&�1U��n6@e>E�h�Ӛ����Pͼ5��i��<���5q@�׍��D5�%Hgy�q�u��];�X��B��8Hj�=Û�P�ۥ������S��,qU��K�B���P ?Hθ��eь�B�ZQ���9	hH��9U��,�=�%֨T�p��2�q��j�d�e,�%��h�~���\������Y���s����5�,`�U��PQF���ĝnS\�(5� T�������h���v���}�
�����Hގ��oBnO{�{�RF������e�n������8������� xt�3�V��>A��������*{IU[Lnp&��(I)u?5��Nn�0l��=�H���h���SwI�8�l�S�oI�nl�-�i1�o�&�%�c���W-��]��/u�?��GL�et�/%s��6p��L�-���/����\Ж��&�rr�$���WtH#䧌��Qc�u͇��6$�mGr��86L�7��:�[�K���\[`��R�-p��Z�P�5��2G�e����mg�%�Kxc:�v�j��}RV}�v;�����I,�$מB��J���گ���hH�, ������`^�HĔ��4����"��S�aʚ��(��M��R���`�2���j�6/��[�̛FHy���B���!!c��P��l�Om�g�8������KacX��ѽ�����_..�w�0����r����(*�B�$�ף��H`ˢ�Pn�����W]�hJ�<���R��,�@����)so�/�DLk��w|g����|�;?��Bi�/ox�ٲ��9i����7�;�ܜ~�J���5����n-���2�7��4X�D��-vyO��]3���~�g�p�(t�&�p�����7w5���˝H���͆j^c���g��s&F�q��󞜜х���\[�������}`E�hƨ���\��dTKݮ����R�ۧ�c���CS��a˾�.���!z�5���9�r�k>�3���g�?}����\��8��Z���5��/��w�R ��2���KyT$@�������� Xgn}7��7��h捊�aF�O݁9
Z����M�z�5c��od���4nE�8�����Ϛf���}B��^�hF����]�E~�`������>v�0�Q�������M�_�WkI"dvV�&S��T}K?��
��t��{��#R)��Xd {F6���$2�ޙ�|%$>&��ξ�����[�^
+3�!�X/��O���U�����c����u�%a�B��X�p8�ĔH�]:�,Q��4��ٶ
�d�z�e�M�C�Op&9���պ����.gvWs��}KU|������!b����mвh�G<��������T�.=��'����"� e�m�v( ��j!�	��+����ŝ�/y���W�s�C���i��ѽ ��?V�ޕ�U�xH��6\�c`����?	��[��Hn�z���UP�|��v��iL�#��z�r��YFJ憖�{�Jp5 �㴒f;ߪ([7�c����М�@8`��O\z���z�W��~�[�]�G����gl���+�x��y���_/�7�"vLŉqv�|VLR����b�Ø��m����A\qn�춄��$v���{�.在2�F|�Dz�_����:v��I6N���	R���� F'���<�E�t��-���ԩ��	��ң����<#�	��J��G�H��m��:k$�'���¼)ؔY���������]hK��?:sO��BfxW30bDI�n�3�@�g����r�� ���������)�W�_{َ-��Y����=ܹ�9�BT�r�?���+T���C��k�1ZWI���K�b�wDk��\�0v��J72�V���t����wս8�M?�J��k���s=tn�m0#�-n=k��Y����#鹇?����N�7�(��(R��s��=WsxI��� �I��ƴ�WR���}Ή%��@�;�o�C����0�i���db�+4n�b#��o��Q��^lCq�0����7=��lO��H��6�\�\��!�%����e.�]5P6C�%��+��m�v�tݍV ���
�Eh�Dd�Yѽc��Y�`,N�^O�M��;+�}b�b�天��^�1+�䤧'?L�0�d����A�2^Cv�oO\��S��MPw>�C��g�4�A`G�_kN�gc"9� �4@	�Q��
��<�_��$G��޶J�i��^�����}�Z�AM@�7m���f�.;����oxk' �
�%���Ӿ~
\�(F�)�y�����B��E�n�I?|���%C��	5 �W��%zJ6������і縑/!e��[�Cy�����h�}�3�9�'�S�A���������|�+����Z}-�]P#����>�� �$'��-_��Px�5���[�r���΍$a)��m�>�4�ȐtF��)�W�ɡ8�)�:ŗ_�h�Qe1�-��O�c����N�m-(e�-�%EA�U9p5��*�k��� K��b�����R��Q���
b>E��`�\k�u��#�I%�޻֚�$�X���[�>@�r4"űZ��P-��~�^r�\0���Om@��"�)GO�}s�03&~`�NAG����GϾ�|Pk���d���K��S��s�
�ĸFF��}�LW[�O�=����
罧�+�:y�ZPZ#Ln�pw~�3�w����0�ʞ?�U��|3����i�|=��3���(���'�fx=Y%�CD	7bE:^�K�X�!�yy�CD��0l����ɴ��6,/{]>"@n :yO޸y��8��k0�f�I��aEvV�Ao�J�緛��Pd!��8�\��8QY_����F���QugpO-XZ��&��H�$$��|^G�$�^�l���c�#��nnDkG�M�Ş������<N�fAM�렰�'��}�Ė~d4�pk����V=0�������P�qfP���8I��r�o�V�6 U��Zf2�K�#��Y�#������7�S	NJ�}�5�j���}n���kM]}���Ct���~���"���0oN\�)�t�w�ͥ�D�DX�A��O�]�����( �!����'�K�õe��Y��U'%\��bZ���H>����F��E�ۜrF����fQc#D��I���z�u��rq��Hrء��m�x_��>u8F<d�"�ڵ���~��]�#o������#����>?��֣��|�=��pv���?oT��B~ؗ��M�ď�D?ZQ�CU%:q����k˰*�6+�_	c�$�ɸ[��이"��	o�:�+��T&�'��A5�fiժ�O |1�_���S;K�em��cOo��i����y�$��v��1�ƹ��oy})ʭ�9���;�����딴����ؼ�]PZo�o�(�T�L��-��K�nJn�\)Gv���tg�ʎ�����u�v�T睂��F�r�ql�^?D��*�BO:I�L�'�TiW�\��Z{����@���E♔��K�Lk�f���H��}�J�0���-��@�o1��љM�W�J�<�"��Q�us)~Z��L���ny����FR��b���Z�v��=���v8�D���,��������2��w2��� ���Ӝ�]�m�3�\Ԕ-�s�n4�tG�3� eZ�~u�?倱Q���&���Z��kw8�^w�skrgK���_�b؊@�8�����k���b��J�s��NN+K��!]��`*�xW3[�M�>��lvc���$��$a ^ 
��Y���B����J)�����L�ߔ^�%��-���AO9���e�#���L���wH��MЙ�H��������L(C�޽�Fv���D�݁t�?�h�1b��� �J�@N���ߋQ����E$�/VЊ�V��Q�~���i�����t3��j24M�K��e
E�&��L�S�?#ȡ�޹Cb��(��Z����I�K�nѽ�YO筒\I9q�OY@���ꆶ��Jy�s|ٓ9�4�z@77Ur�!�W�_ň˰x��pC�� ���E��#9��WnX��_N��ň{�f���%y@G�{�[�%0ITl�@_�m,��� ͉r3�ה�3�׍����B��A]za�5��Q���T5 ��oW2��EuR�`���:�y��~�EN�}9`���6�K�]�y��?��v�?��O�P��+���SSqw��WA����CV���WX�+q��{�H��9m$��h���y�"b=¿ly�H��}k��_�>�~=�Ȣ�<��}��R�ײ\�yK��	�e�Nz���!\�����d�h�#�cp��=u�;���&[��6\2��۴5���a�J����A���OZ��~q�e���Tb<�ё]0�EW�����P��`/o����s5��U&��;�����b`�=�%S����|���]=�9>P@ �>��_��"5o��d�\5%
���w��(l�iT�]&�1� r���w�YM�h��x��hXRE2!n ��}%	?ܘGV��
 2Ȋ����e��ߣ(FW�a|nfYW�Ey!Սе���"_�J%m�&d{O�>����Z�,i_���Һl�����b rAS���`OZҮa��9.D:�p�	�f��r�lR�|81:��V���Lrv�f)z�v?N�n�6��W�|�2�);�V�zg�whb&;���E�Q{��o���Z23���^�i���a���0|�j�ݣ�dͦ�'C@T����⯇b[i#�0���ޗn���-vԻAD�K[�;��a#󰔒oÂU@�n��(.���;��H"%�D�H{;{��`Ӄ���{v�1������N�~J��1������}�n�)͉�$�_�B^T0�S�zRJ�\�3gw ���l� ��Њ�^#���P��}�tq�rʋѰ��=m�m��]*�Gp��B�랶���!(F&��Uзk��푃�_U�%���XO�)̀�\T�.>��D����,��N�p  �9��>�^ӲءqH���
 ,:�z�����G���&��{�^�QvJ��z�'
G�������'Ɉ|y��:[&/y�2A�R0��3��pkI�`�H��ʞv\e=zf!s�1��i�b3It��K�R�aZ5l`JJ�89� �[�1���(�b�4�0�oo�1��n���jG0o%�,��}x�p�kԆ|�-8���p2wa�R�&[(.�j�za��G��D�Hqo�y��I�4�Ť������.��z�o�����VU���된�כh#u?����n�k����A.QQ>WG*��*P�=͎Ica��Q�XOw��s����v�CHM�9]���(Q�9LԨ�2�Aö_�h���B]p�8
s��!�\e졭?�+�7�B��dFF���93�k�?��r���Jg�#���#A@���������YV;�_Q�������v6D�/Y1Hh�3���3�Kw�]�H(7�bZ�Y�$�z���L�c�����1BB�UT-݊]nuU)�vՌKŁ�CMo�'�F�X�*��}����q�1��&�l6�a���I ���-�����n��m�2u�S͔�o+�`��u����S7�{��?.fS�)r�	�� �H<u�o�Ө�.�8J'�wf�켻Lv������7�$�W��ٸG�u�����[ݯQ��]ܶ/n�K�����B�?W��}��d��?}����(�	�!Z������aG��J%M��̤Ԑ��rرˆ0X3��e��(,��c�O6Ӓ�.47_PI���*�r�cTJp����^���A��tP�Tj��#�I�R8�=�y��:uY�E�Q2��>

'�����L� �^C����b��4%E�n�ȵ�a���}�I}u��"��%��o� �ا�wW��������:��Ѭ4���7��� g�M�-�/���}����rj咩`·2��㝈�(�/��ē�	۰�0K�3xU�����0�����ٌaH�~ c'u�9��Q[-QEPtF�=r�e�[U��uY���K�r�(�V�Fx�ӝF���[�%y��TM��m5���$.�ю%��y���Q�U���/N�x�/}�N���sIb���(A�vP�xOA*R���p�ຜ��=x����/)��O�|�c㲜���OBn��T��Cݩ6U�
�M@�MYNiԩsI۶ė�ȗR��/+��}o� Z^�{C��#�3w��P��t�JD|,�z}� =� G� ����6!~��Bd8�&2_o��͒Tr�Ӯ���k�>"��u��'�`���v�)qaֽ業N��Q<k4bg�H,�#!X�����OOzQ�\�$Y( \Y�)���/؋`i�V��;N
���!�*t�#N-�ƅ�߿�hUE]�?�n��K9(�^Hw����yS���T�D���$i�u&L�~�Ū��d!~s!F��F�(�Z�LIԲVs��G�I�,Y�"�h�,<�-� ��;*T^. �N]��"����C��4֤�!���{2>�j�3� S��u)g뻢�����ݣX�[*n�v}������P�S<�T������,�
Ǐ_�0�}aq�gy��p��w�Vc5w�2�Ҏ3�c�Y2���X��S���fD�h§�Q�ۉ_�-`)�N[��������OCL��K7��7��'o1	&G����¥���.�>����o�مC#�@�>6KX���9p���NC��d�j����r-���c��\@@�Itr.�J��!7�x;iI"p>LLy�V��ғb@u�1���������B�?'t����S9SJ#ַ�%)���]e�ʌ��
ü��-��O��6��h0"��Ҿ�$��4t���̃K|�_�֩���[�|;(BE5�K�	���Ӱ�f��ep�=���=8��M]����*��7�;X8 �f�E���"$�R�U�������z=��#!���*��}������~-�mѢ���{"��?���#��ո�?fY-��u�ҳ,��L���ǘ��lV)�eg&�y��eb�[�y�;^�v-$��DW����f��D��ʶ^���O�.4�c�p=���!�fR�cX:��V>�$[c\NBt�_���V��P�Jd�C�^;R�k?�q+Y�h(�;r�1���H#gc�p�_rw4�M���܇���0>醡�M铭x�c���l,D-�x�VU�rJ�h���AL�Q��H����,'K!�o�so������Bm����)���.3&��i��v�?�sO�׭[�h�x���3��?��1���q�d�H�=��O,���+1�#��~�kH�۝�G��4�����bfD$��uq��6Y���
hS�\��(\'���1��3���;��6�[G��Uq1��gU��	"�Nt����"���{p��m�(�'k�қ�Tfr�5#C<	��Ί� ��j)I�o#*��On#��|S)t��ؚz�Q��(Ka4��S�������~� GkP�%W�ra���#b���K0R�g�6�z?ݐAF�dt�Y��*sv��|�N�^y�?�A�1Dj�\��TX�>����u�����3��N&�����o��;��T��Ƹ��RA�}�P�PҮ��Uo���A��ÞF�"��g����[��3v�+{��x�=U���!�g��B@=��*G
��btm5pў��^�)M�jCynl<��c�ٚLj"���L�$a`���U\S�2K��#�'B?��@�mȜh*j��^�?B}�h�_��H��~�ڤ�;ua�w�m��ݙ*��Q~ݟ�՞�!(WW�S�Ȕ�\�0N�M�{oH��x�̓���;�-"J�먛Т��ԉ^g��OJ9����j��|P��v����1���)���d潂�JV`��׋1��Qb �����~J;E��#�*��Q�ғϏ?��4&$���~U之̼��(���Ȥ��"���M�!-���"3�`4K�$�ե���5�l��~�,�<AE=:އP�7/��^��"@�`�� �QFO��=��/�i��q�u(��K�����oeH��P���3�[�����Y�\�bA}]&8$�!4�,�(,�Rn�Y�n����m؍a�����-ѝ����x�R���G_M�(�ܥ[�P���攉�����k�O}ֻ��F�e��K��Q�NtBX,�|72��!$��µ���-���f����	A��P0:�Ȼ	��Kd#t��U���B0�荹���$R��gB۸z�bO����T����lK��M�!e��U���Y�%܁[r릮P�;���$4�(�D�=P�UW��YyB�d��0�'�1O�ɋ�r�%�����$���$�%�9jd���|e�WEa�4������>�@-�����IJg,�.���Ee��3$$K�Ze��F,�i�;�;_yt0g��:���n�����S��� ��pJ�{�H��Lj�V�� �I���q�}��F` y�j�\Ƨ�Lq)�i��-�h>�3'g��L||60�&�p�9�w��\ k�XiC��r-���e]]�!�;�����T"n*�����f�f�eP'�Ed�zS�Ϩ��L�?�+��n��1F��zX���"~�a�Qܢ��x�R*D'Z���V�^�~����_h;fX���H�Q�R}ǝP���9��d�m����C:(����ޖHG���5�E֨c�;��9��g�����^!�r<��(�.,؎ꗭ@}],��Pp8a���(4"��^�҈���w,~�&��='��Tq#�`���|�kbp�e6��H��L�ei%"wzA!��oZjж���Z��)��\��yv��%���1�dE8��qf=eͻ�Lɰ��qʗ��0�
8-�w�Kir�ջf�V�<H�bõ�M�R�?���)F���l@�bl��pB@L���t��P�Ah��!l��(�N`FB9�D�N��	����j]�"��eK����Y�D�KZG��j�$��%����1K,�E�����kg��w�65 }�WN�������u�8���I�!ƪQ!�P��]�Uǔ���E���ZɈ9�gW=Iم�ctt��!�ط�ζ�흛���e��G��P�-D��9m�T
V�K�>��G�q0����(�Er��/5������}�� �Y�W���;��)��F���0����;����gB^;��y0'ږ��>�4Vț_H��K��p~��T��lF�Y�Mܤ����Q����q]t|�M�7�F�"L�b* t�WG=�;S��F0��(c37X!s��>��a�+�{�Q� �ZL3�r쮎h H�u@n~_���89W�Ͼ= �� �V�ՠ2��D�hU�� V��Cv�#����-�x���>Y�b����DpTx�3A-J��1t�ނfv�m��m�����#������
��	O����8�*\�z�i�W���o8�ī�?�@�)���k��d�w`���n��y����
[�
� �a��Oc1&��K֊H}4�%yDC�,K��7�j[&+7y�X�~1Ai�b��Ⱥ��*�ۊڰ�?/XBn�;s������r}�ڜ��]�4U�Y�O���"�d�zNB��MM �0N%9��逮p��9L��ݍ�i���P���in� �R}Lڎ�+ �.�
E5z�
�x�c����nN'��W�V+�tb~�L�Ang~v~1}t�b,r�c�c��Ğ��V� ��t��>:65����;f������S�ɘ�v~���s	��`�!�z�Sux�ʤT��p:��i�Xn�u�Y��j.�L�6�J(J2�Xq�7OS{nlY�S#���*O915����b�~:�JC�[ĶH�@�jI�A�W��n@�k���.�1�w<A,&�@��:�3[���jif#�yu��<uЁE���o�>4RM�ŰY��T�o��6�/��w�h��Z;�}as�٩�-���� U0������n�>�Y��(� �����Rظ�)6=m7���⒑1�TL�|ĵKm��D�]��ʧ���'�S��w	rt-u�n��~���H*�A`��f�4�n_q��ܞc&,<��3�+���i}�'�	��mY]�*������G�!���$h�?�T��Q�8��xUkDQIB�@6޲������C�_m�4>Lp�i��4O�8�%iӓ�[8����+�����4�h=%�,(�Oyq�=.��n�����}��ƞ���mM��塚�T�y'���#=�	�����LSBp]����SJ��{�`-U�۠�T�@[�4�y���T�&�ψ���A�e!"J����RA"]�ֺ\a^�6�  z�yCs
Ev�Xi�j�����Fv��w��`���K0�t���>���oa�><<U�1KM��Ϭ^9�����%G���{;&�8��+'� 4�u����h5�"���b	o�Nq�����  t�|O�;��X��P���������S�8�~���Q�r�Æ�N����s¢2aPV�ϋ{΀#!���P�֟>}SH�
/��� | D!!�KJ[�Y���d�B�Qp
N�"�<!��A �b�X�b�������N�t�VbODt���H��^R)��E�0{
��B�Ksg������ȱ|n�>P�׎�,C��I	%w�ҘN^����V-��B��>��0Y�*_i�̨��ކi%zU`�1�������������C=+)�,��>9�}����&5+`��}�dK����$�E�>}w�#+~�N���d}�Y�v7W����C39 �3
ݠ�a��_%o&EAft-��$�J�����
Y����ʧ�^�N{4Ž��J���N�1��{����1�lZ�n�IV��o�7%��a�m��Ξ�=.���Q��WN�y�^m�\�(h%��H�<sL��- ��,��[�d�\&�s3+*�Vw��� �\^va�V�[�|�va�衣���l��$;\g�������7�;��ĴE�Y��Q��>׉N!���j���d���$0���t�2,urg��x˙�,�dy�F�s*R�0�a@1j��=�L����D�qL����(�8��Q�M>����l�h9���	��;W��?*WSjZ������L��H��S�c����0�T�-Gz�c=��������X�-��4�]b��0ҟꢬCtZQ_;o
#ܨy�1]a�f�H����eX�[��F2܁��7AmR��G~�'��X�7L$Sྱ����jy]
�bt�W�kz	��PWe�U���x��)��"�xc�-�^Ml���r�+Yl0����&j|2`6l���3V���$by-`��5��n�#����ZS=,�6�p�R����^Y��g��ͬ��D7e�N=���C4c��
s�� 9hj+w�tK����i���|A�����psEМ�G�ic��i�#c�bŮ�Z��@��J�E�� xɍǼ�}(�2��DJ;ܡ����2�=5L�W�)3�RҖЌ�p�B]�'��h<���;��2WI!7�}�J���r`��g�_`Nik�Z
��Qdb!���:(�:\��@aYh�o�K"gk(�!���Tf(�r�cQ��e\�b��ph'��u��V^y���!�D� ��.ƻ5��g�i��v�9��\s�5����%H.���R$��4cAٌ�k�I�r?�Ɇ�LU���� ��@�<�:S���s�Z�@SN��ц��>wkܸ%�9#y��E
x:�ݨ��m����pܽFXZ��a�+jw
�n�9��I��!�p9�n�nKJ@��? Ч��OI*�x�xL�q�g�����%�+0�'_@  <ԙ���7��8}Ut%�#�у, ������+�(����1��_�lmf|�EJ�`� ��H�x���GphWjJ�k��A�C�SL��{�Q�-���O���~�e�s j�z:��2�h{U~���#�I.&9��> ���X��~Ar��y���l�P#r` ����)N)����Db��K6-�f�;����KY��c��8�[� �˵P�nᗵ��Uߵۛl�~Ѻ��{{z���}L�=V@���?Ϫ�M�/Y�H��9��>�`M@������D�.�§`�����!z��vi�^+)�w�èw,bW�ߔT�%[���p���`q�}��G���nʽF�Z#�vg}L�I�&,l�zSX���:gqD�����eɨ��� SU�4ՠ	����{���H�#�����r��G��p��[>|V��q���!�sR��B�PS�� ���c�U�jbt�h�^�ݏ���r�i�,T�� ��0iRt������&�_5r||+n�S��=��P�dl�kD�K��/�^%$�\��U4�Rd��F���P+dv&��YmP�.���_x�*�ǉ��597�kS�-7��=�����*��õђ��
���<B:�ٵ�ґt�ą"��'����I���d`C���b��@�V�E���L�q�7�Q��o���q���-aN������5+���RA~^g�1���F��9��C �P�
�.O ����scd]���,��� ����'��)Xǿ��JN?+��!�'5b`��P���!B�'yh�)�2�~���A2����=�`)��H�@)�y���`|�ʺ8��)8C�Y���8<`��)��E�e��#���'-Hk%)E��m����
B�̑}[!��ۘ<����V���8�z��(�Q�� ��}�;q�<�� +n!(f��� ~����t�t_{98KD(��^5A�^"�:h��ײl|oO�C(�V�R=���~'�e����k���hh���>r1��@��e�J~��O��><�N��IΝXRf4��Jq�[�B�*���C�V?�)��ы�h�N��ԮU������j@��H�a=k	S���u'\�H�1e�no�#	ô���Nl�	;�144D�9����sTw+��2��xl��hu^�Ox�Ԑ��խ6�r�s�y�F�tUx:�i4���JٕM�֦r�R�~E��-iI�l�[O���E�A!Wǫn��P�&��l��Z�������Y�h��u�	�ۗ��y���� R�)�PH�ms�y�K��nI�sI�3��A$�;��U���;�G=_�<,3)�C2�we1���:C�t۫\F�nS�)�]Y.�!�I��ί�5���2�f�h��B(e,a~�k���l�����r�@/4��
��w~Hfx�J�>BN$
�|�1���ե���j�1G�+H����Θ`Z�=t񙺄[BY�N�oCm����N�9ɋ�k�MXp��o	�,��p�*���A{����}w��G���A�l�d�g���ѪN,)��cz�4i�[7�ΏR��W�����0�
��̠��'ӣ�RF��10o����V�< &�����PHl@`1
N3�r��S
#T�h��h��/�"ق����8'2Xf\�v��kS�4_�9ɟ�LP�t��fo��a��Nt�ZP^�����Q$b���į%l�tR�@Q�8j������sT'~�Wz����QF�y�j�Zx�o�H�*�ϴ ϑ'��LʺI5�	$?��?ݣ����s�Ë����g���'��A�;b��^msM�����[>�՗�d�Ĥ�BE������}-�v/ˮ�7jf����F��iQ��T�����p"ǹ�}��c�T�A����^cc�[�>��4��Yi�kq�0��3}W�=�G�$?x��ֿ�`>����^d���Z~@6���ȃAiG��D!�-�J᭶�~�!�/3
q����^p�SHo/NG2wiPu6�q�uw���Cl���1csA�@ ������a���q4�le�@�������u5M�@��҅.,e/��{<��6��;��\����V]4e����\H����{/�b��\~��hiu�PR���O�*�҇�6��>�e\���_sD���[�":���a�93���p���|�f-C��hٟ_��o�-v�E�į�E��;TQ�\^n^N��r�ڽ,5$���{���>ܵ)���y�Hlw0Y���@Y��0��a(w�4z�y$s�;9f��<�N�;Z^��-n�*Ew�b �D�*��%���9(ZV@D˯3� Ss�ip&O{�I���#��ս�7�PY5,�%��u��?C��Ji�(��.���~q� �GVOˎ�͇p������_�)�K:0�2��\2�Kkp�(6����6�����accE4[j��#C�E���C�p�aP��?C�1+��ڣ����e�"��~�?������SOTT�$bu��=;x/�8Y̛���#�>�S���x�߂.M��<ib�h��nLc��+3�c���)D(�Z�)kY�3�m�P�=T%5��0@�g`��3��X��s�s��T�f
�Bc�Qg)˾� F��I�@�g�Eq��p�g~��{1}p��Og�:8�n��bq��4����9_�[ձ^U\o1BM���S��` $�)o�����Z9�9�W�����9R�\���p{K��4Nݲ�)ʫ]���a6L�
�O$�ݹ�8O4��@��nq�i!r�u�I��2n���+�:@�_z�^1b����\3r��_���%X �����AjI���K�)0N��
�jѫF`�'�gh�B l�]w�˳��Ґ�H����̈���\&q�;��;K�0���W��?���+&���պT�E��5f�-e�~��f4KUxFB� �Z�s�·�����h���QOҧ%�ۃ戸N��DD;�u3񲦻�{d�ۿ,����XP���8���9t���e��,�,�w���eY�V������8)s'h��s���H�1g�n�1�5O����@��;�A��8��὞����r���j���{%�4���'���lA�
.��mF|,RKTl�����;*�!�
�����M��]�o���&�64���x3V�����^I04{���%����,�����<�@���	��3�A!��5>�a��&�\�OC_�

�Qw;�&aPK�����On�P��u_,���Çş ӳI��4A�~�ڄ�E{�'� ̉?�2N�T��1��ULy�����c��]5�f��Ƽ�O�H�k�K����&��U�`�+�:��1��Z�����]����ah�����3�XB.ō�x�դ^^`����E�m��/��:�γ<yj�޼��6sA#� 7v��=��F˵�)�Il;;�r �^�e�B�>q��x,8Ɵp��p�.K4:õ�4�h��Bk��W�һ�X7
�
�����`�d�q4�1�y72ƄP�t�̣~�ua��ư�&]���*���N^Pv�Q����v��$W�r�Ŷ`��~I�'>���t;f��Ң{#�X�m�Ro��X�pz ���>���{P͸%�D j�#J�[��T*���w~�L�@-E~������UsS�Z�4[��Xf�H}o�q}�i;2a����R�����bu��j%�M�풁M��uig��j��4���#��L㢇�4/��O����z֣��/�7����|�4�=3��Jq$�Bt����e8��g6�at(����FȒ�#L �F)P
:��0Ѵ�C �,�dM�=���
�����,r�9�>���+36!?~4�_�v�����F� �d��y&�]�F*��kVĶS�y-�I_��c��1j �9�/U(�Qb@�ԕ�*f�����q�N-P,�v�M�߀���t��I����Ω�U�
���te��]���ݕL���˸+=]��g�	���bE/����PԳ���u]>5ԟ�٠������l^���Ei֍�w7�:�E�_���Tq�;<�!
�lv�>m�������֊�&�#}��qͺ��/��0��wF����<b�[JWQqJB�O�L�Ǐ�!�7�m1�l]M�)��$�i����.l9|&=/����]b��#�f-H����</{�d�L`޸��,���c?�V9Ѡ��K1S�s���}{����SLv�����J�]�a�@ÁH�J)�"��[�!��M��ӡ�Ҝ����U\�+�%t�9H~�/ZL�_��̜�M����d!d�$�Q*�F�V�&���	���v*��'�B�y0<�n1+����}բ���F`��"�gk�����8^� �b���ˠ�J�b�`�s�gE�X7��ȣ����0�z}��L��;�5Z�6��@	]y��yWUD
R���:@ �9B~SLZ�r�`I���:���9�oG�b u��z��V�!%s���G-���4���?����[�"��ڗJ���IQċH��!�ڱ���<����F�۠Q9�0o����S#�'2�80h<��SL܉�g����Y�f~��<v#�����Փ�
nJ����åтŝ�x��ɧ{-�x3��gq�*<'^;}�z�f����{��W�%v�Bx01Y��� u�u#�$�GoR[�܋0���hrWn�
��$�^'��
�H[KC�(M>�[��$⛮m�)�ǅ�Vg�H���I���JP< �,*��s7:ť����S�oS��/�{p�ćνg����g� {kjk�I�\F��C5ʺik\�=��^�hT1�<�\�q"��7�=�1���׏~w�_���{����U�q��{��T{�Zj��/��#><%�BtGm���f݊� 1m�R�L�Wq��l��D�(F�;0�su���ELA�^p��\�im�pP(@�B�+���š��:t��aRy��e��6��k�3b�Pȗ&�$Z�y��R�x�:_�'�}�#��,D�1�P��"�#��e�������8F�^7�o�͙;
n��(���`�vۓ$�2�`��AQ-$<,�p�Ԁ���"ø+�}�@㙆��Y��s��)�<%
����w�v�4m�~���C߿�j�Z��+�