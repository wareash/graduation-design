��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� ;l�Fv1�Lژ�O���3��������F����Q?���b�V����Ţ� K��Q�G�D��i�o�Yʫ�|�F�V{:�� �{��LBB���Z��^sӽy/��[����I����k���'_hx\�Ƥ�?���ƫC8�r��j���?�[�b��Gk����s��$E�C���Iv{��Ϗ.��R+!9u@Gf6�e+~�7k>�_3�T�@�@����58fW�o$�T�h,|���z.yhb+�[��>���W��Oѹ/t7y����8�A?X�Xw��J~���k.W�$�'��(��ꉑ'[J��TF�S���o�z󷬓�I�UW���{�|�M�a���@�F�J�Q�tx�tEV��Z��i��lzt����#��I ������T0�=C��'1#"V,���)�r����4p1����Ɠ��LS�d�,BbD�י��)�@/
X����0�9�C�'�8�5��I��*���ŀ�К�;R�g2�9B}������Qj����F�5#,VF5~z�wY@�g�ږ���jbY'��&W���Q��p�>��@牣@N�#���Up��]���ߏ����\c0�4i���jK�tƩ�H-c�����d�@+�FRxY�,��~F��(��y���^�)P݈�k4<�w���Z���?4���E�}��_�á��š�0ޜz/B��Ѽ��#f�݌$��3��z#G �W�fĨ��H+hnؐ�&�,�Ɍ��9�ċ1�(ֱ�{��v�RF�T5r�����F6�}6��2l����Ɯ-pw@���
�O1���3��~1��І6	��v�A���@�e!����� S-����193��n���2aD��T�=��@�j���ksrK�g������Qq�M!?N[Qa��R(��e�����t�xAEƝ�r	��&�J��Zh���dDB�����-�<�Iπa���@���+{\������!F��^�JA��d��0��*�u��|��``:	 �%�&��7�8��Nex6f���r-����"�2��4�C*�tتp�v7��$�j'�փ�&�t/��K"�5�@V���ŝ��(�\v*2O��ϸ�Y�, c�:�j2� io����y�L��H:�a3����4;�
�+(Y�),Ml�Z�}�@Uס���=�Y�y�/f��-��`�@n�7��u�F��A�>�A��T""���~]-=�G��IEW]�߆}�K���eJx�B4Ҥ] �f|�p����[�����X�o�i��_=r���H���kY�N���u*|G�5���" �v���3�UK�6��
��wO*#'�Ǐ���q�H�-��u���0+U���b[W<V�5�K�A,.��D�3�+����aFu1D��ѽ������g���2TL�)���+�o��{���%�~ �"d#	���L!� �d3�q�5oP���j8�Yw
��q!�ű~���L{�sf��fB6�����oxN�mP�[󮡰��+�y�2<;�� ��O��t�u-�BNcH%~7�k�Tk&�DM�|���gySėb��hO�9���d~�=�Y"��܍�l��=����U�;f�)�p|�8gMe{��W�#^~���_n���9$Z�zӄ0X?�v3��9�`ᏣV/�g��c���!-�id�"�ۓ�u�(~0#�`�����N�$�޻��얏p�w��Ԝl�q_�K�s#��3�~�C�h�L$�||��i��'������e���>3�p]d�QY!q��gjT�ۨ�;��`[�ˑ�'����%blqs59�C���f���:�e�#�a��`���k�V*ܟ��Z^@4�ɮ3�� +�'Bux���@i�������D�H�c=K����R��w��%��N�:�SB��5�_��{�R�����k��Hf�p��Tz�n�e�eٶ #��
�7T,��L�@FR{M8��SZ,;^�J���7�af\�y��]��>tϠ��Ky2��Q�w�w�'+"��� anG ��������i:6�|���U�|�nI�W�8k���|����?jwL+Y��:��YJ"T�Q�a�O�ƣs�i�xs់�3ԎL�Fq���