��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����Mڨ��˳0]��?l
�4�!�ߦ����"�p8"	~��kB�J)��NbM�L��\jO��#y��r�3wA�y�}�S�{�����X�.m�lM(��R�g������B�*�NV�X-?����$��$�3�s�`;��y�@�u�ߗA�R�|�Ԝ�+�)]f��������҅i[^�"[��t��00��6�ĔR�*[�]�V�t���9�c%kz�Q��*N�| ea�z ��@������mU���h�$}���~�k��'C ��� Z���>J����ׯ,�'��3@akCc�U�U��?��a	6S��K󊀧uh���Z��&���9�+�)�b�В���ɀ�t�]z[��z�/`� !g�!*��P�����I�<V�� /o"�����@�g柅˳���.���5����9�i��)�!Ҏ���f8�vh�3�Z��ZC�:3Ϲ@�+��&�Ư���	��������Ϋ< �����"�����!b�'G����Z�!�R�l��Ã���3�����y���H�>����/{���?R%|��n6���gJ�2!b/ΧW�}�/FM��%����� ǜBk{�.�-�ّWz�*J`����'29�05�J�NYŪԚ��N�F2���������q��y�-Y�	����D�0���7��%��,�-.�O,P�y�w	�	�JT6'�Z�Ҟ���4��\��י����Ə��g��y��E��q�"�ӊ��N���H��`����=l�r�Ed�tP\��� �c�G�����/�('�'˷5����+��3]ʸ�:xõ|D,"���V�d�@��^Nm�D�dK�+l����E�ȟ��_��O�՟	����ȢM�6��������U�²��;偐&r�+����q���_j/�/3Ew�?'�Y���7ϓ,4���W�X�`]���eop�B����nIN�_K�����+�-�J��^��8��c�.)��+eR\_�-�/��?���}��@�|�VBp�zq�4���tsT������wPφ�(�,/��3�3~����]4�_x}����M��t,�Wv,�,�t����#���ιXz�^U��#|n���q��LlW�'_�@aQ�Ѽ��Սu�7�q��"�u$��NɌS3&rCL ��#��$���&x���Z�����h�!�(	���/_X	ṱ��
)_�� ����T��)7[�{8�v����w!�$�]�����qo)��N��1�K����ޙ���Ju�ɰ$`�9jy*rv�!��9@:� ���ɂ+&a�"+�U�������1E�����V�]����[�Xr�؝e������{O#.6�|�����8fK��a�FZtK���[sx4�/���J$�IxG��oԍٷs�H�Tio�w3���Ē2j�����2|O��6���a)G�7>��J�����k�΄Y5~R���hH)��cX�������Aa�%��BA�>ՠ+��g>��T�\�@�`�Q�*=Up�o�V�M&=�ї<h��%�R<+jhV[E�k.�2ku����B~����̋:������}z�FD����RAmڴ��������b{IJ �MXN;,c��,yf��{�@��lg�hhQ��Vư��F���%k��[�e��A�w�@��N,�P�����{ٹk~�� �J2{e\~�������"QUXa�$���Ԍ�x������UrAJ�:�PN��|<Ƃw�j���Ǫ\#&�yT5w�x��]��G���u�"Ϸ7(18LT�݁�Hz�����^�w��-�ی�C�\���G�'Uga(��� CN8�YW[�&.�m�tҶF �?���K�X����NǦ���rH8�	�!e����WV�E��jk�;ҫ������R�m#jK#����x�/-��r!��ҵ�Zv)8����S�����:�B��˔�r|y_zb9@���B�/������ɣQRB@��a49���I��Ô+���{����2g�E�.�'Z��.˺�=gY�Pm@�g��L��A��8�8�R!���oH��!�t܋�����O�1���M�W��~�LN�n�i��;�v�T3���k�<����)�Ӎ!ӯkx3��/�e��Bm�s��/�ޗ&,~��|,�=Φ ��t���|�
$�����|��Y��{������M����C���gX��	�$�Tށ��M�hb��6����' ���H��P3��Xn���酄7��5�v��p*�O������zl�w��DHK�̯�Gp$5�8�'�8t���R���/�@�a�U�Ւ����\Эu�MJ@�*G�B�¸���ɸ�</�铆ћ2֡1�0�l�=�����. �)�<s��-34��Q�{�m�[q�.�|��M4Ǿ�y֪| ��L����C@�������