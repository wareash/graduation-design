��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|��&���i} Ĳ?��\0����굶�%v�@S�8Y��,|��$�ѥ#��/�z)՝�����jq��|�&C=u�c�b�J�Q����1[O0VZ���@-����[�?���E2=UpuX,-gS��6\M��L�8ʉDA�̼/ԓ��*2ְ]�y��)��_Ѥ1zbd�rlx�N ߾=���*�D�*>�=F��k�=��j8'-G����Y�'�O��g�<ʚ�t��J�Z��bC뭃��������������>f�d���X�����mK�f[�^n8���;bN6|�>� -���Hܬ-���q���c!%?N8_�a�d�������>S�O��( �Hw5��~�u{��4Gvr�/b�� ��9
��ҁe~�+{�AM~��Ʀ��iٵ^͵g�A��eg��>A�tҹ,Z����j������a��[�A#�sqP�^��%���&���@ ��ho�=�\�a�$d�7��!wg�q���<�Ӎ
���݇K`g�k�ގ4����\b��`�j���v����F���8*�� �%f��h�K��������nw��Q��w�� W�W8H�3¹8��w�]D[G��|l0�A���ҷٚ#go����uo�(�b�u�z�%�~柫�o����A����}עN��2�o�TFd��br-l�m���6�N��'��&�7��;��+KA�u ��ַpW���^l�
?Z���~1��� �����62��\��}��UN��J�K���?���R.c=9�.�x�e&po���� M�?|���Y�oH@��Q���MW!�7���H�Ơl�g=��0ܓ�w�#��z��t����_\s��sf֢a��c��*�6Bf3ůh
l�h6"υr���(��� �����Ū?^4
SR�d	�;������H����yP3�w���\��K�Ʒ�B�Y��o�<ka��|VE~�-fk��SX��a��|(E�� � ǘ�����kHNZ6M����<R�Y�i)uV�ߍ��~5;
�q���5fmi�����\4�K���+����Q4VP���N�P����s��ſ��h�s�l��2�b���+ĸɺ�c�睱�9�\�[��Hr`Ĥ�%[�Oc^�Eڍ	�[E��!����#T�Æ�J�gEM7;gM���TDH���d ����Wl�/G:rl��am�=�ʀ��Ȕ�SO���ިtf4���\�Jѥ��~K��=�H�:��0[�H�YK��K�#�]$|oa�w�=V;�h�+��.$
{0!��7��#�_��	O�J{�Ul81��I�R]TN�����9v}�7��kl��uR�X��a(�js5Um1DW�,�n��6 �����}rt�p�F�	Xk���Gr �&N�ƺW�2i�et���`D���l���0�t���K�A��L�b����~g�Yn�� ,XW`�w�0�6)7��SVS�R����t'A�o�H����K�Kb`N�Ȝה?�L���M�[*����Ae�Β���hJ�cv�jP-�F�x���V����ە�\��Fo�`��G�z�A��w�S�&��h$O=�_X��G<��"
��y� z����4��fG	uk+�֙�$���U���[L�!��E7��H|t��������Ü�~�.(N��Z~W��9�C���Vj��2G)�p����rd��X�	b3g���w���j8��Yv�E��R�a��HN�?�5�6ɨ�5��^%Ł�i~��4�"�n_�B�T�j�A��l��=	���2��K�����b����͟�X��NI*|U�+6�њ�=ˑ�L�͝���yΡ�8�-x�A�R��N�O�x�揼y���6|!�A@�o}�R�X{�ۈ�P���x��L�:j�)��^�[�^��ϭBNxw�����f�_��n&���)�m��"�����ү�4��3�C�_$�2q��j��TAwH_����^����{�V���|�O���p�n�~+��#S�	~�L� �f�<fk���`_���.9�ٺE~�c�>��U^����r�л�.�9�:{�E7�3\�	>�F�y-y�4�Y�e�^�,�x��+VJ�D���(� ��~
�5���G�Ч�|PK�1��Ym+�3�T���z��H�[�ŏ/(�Ο��9F�Ue���K����X�n�&w������
�Ki@d(~5!x�u��F���̘6���]}"Áu��Ox�c$�	ˏ������y��#R�n�������Bs�#fSW�.ٺ_���Լ�Wd���^(d�K٧����뢷�()�%���>�d��=���9���g�q���	W �<�ۇ�[)F��Ac���#4"Q�x�1�@�G�-�.��Bv{;���y��J�TH�eVy1�<]�����v���k����iX0�o��Y6�Oݼ�?/ GVg��t��((րK`�ZvsXt���%*��z�Eީ�(1�-���lwY��;{?6��
���
K��dP��	��輴�*�r���!T�=���� �x�Nу��޵R�Ld�؇��L�T+%��,�|ƱJ���`j��b/�2<1R�<P����*�����p_� ]_��5q�`����q�c��g�:�C�o	��W��V�>��~9� �Oh�ٷW�#�m��~4�`�2x����a�	��|�%!�$w���*�=�X �y��$N���F�'(h�5L#��!$~yh����wkoӻb��L�y��wPK�Mea��\%��w-��З(Wȉ��57i�k��GMЋ�yIv���˩� F���r�x�8�yo�Et�>���n& >���nJ��"D�K�4�~��}�n��m�T�����H@[h�:� 	�z���¯��]/�)6H	�x�l!ro`ԕ�):�5�ޤ�2�����i���A�5�����M��yĻ���:CCy��q�UP����I2K�U2�>�l��TFV~��� ����+ї�������_�G�)���Y�����İ����{Ylm�\�م������:2(<6P������^�#��Ts���8��Qҽ�!�Fn��yf��ndҜ>�0�/S�;5����O6�N��oO�a�Gh3r�����U��p�z��-a����x�$M���)4v_@x��T�������x�7#iM��ｧ�YX���n�XS�DY��QF1ڴ�ʘsS�= ��i:T2��f�WW�N =�v #���#_z�����:�{ٹ�����E�gFu:���s�Bt`j�=�� �+�%��O�@�(è����/@��_�o1���L��̎�onW���������6���}�N��B�kB�R�r&�L�Wf� |g0��Ņ� �E�/y�7l�C�U�2�X����{y���f���~3k��J�!�䘞"���� ��ǧ���Ea�[���N�9�<����{�̛
��	5���$#�■�D����T �������=oFv)�S�ҧO��s�)-����η����	��^�ޑ�z�wZ�1�n�o�8$#'�s��H?��bNkj�<���6~*����כ�I^��@�sW�[��[G�"e~=�Gi���c�X�����bG��ɡ�)�{�������s�0md4��k�jZa��Q��ŶK��X������w�8��R��.��_��Gڵ����rFͯ
�\V>�-���{�k�ݖ��Tɻ�������d�����IkʐW�kτ��[��*�85D�q�4Ch®���V�/�?W�O���4�zc�����_���P>��sv�]E��e����C����r��v��R!޲�d�P��_��ץ�A�_W%����@�~��`�x�����i�fe��� ]M9���Qj�|b���j�LX���I4�n꽽��'��q^m��:z?�|�G�i���s��q��W@Qݪ��q����(%�¸&ƌ=���k� 4^�l�i�U:l����l�u���Ύ�{�������wP
�:@&���`I`�lU
1��7�T���������v'I�� �ξ���(�hh#O����rv�A��}��(��6���K���
������>�#�o��N�h�Ռ9��'����B��!���V�+*@P#����h9��؅f<�u  O�����R�8۠��J��ls��d���^�@�Q����M��F�S!����b��]��KD�d�	*�P�K�D��o�)�P��Q�K�L�ѯ6���@G��h�ȼ��j~p��	�0X��gZ�D!��L��<�?����]���8�䔚-�p�Q��Ò�U�ŝ�( ~wt�pr�4�% �������W���<���3���J1w0Ȧ�k��=�5����q}��#ָ��-9��Z�%ԟ����aX�M��"����[m�����ɠ���3�V^��;B�w�h�'^��8�z�k�h|�>1Pt�W��j�^9?����bۢ5�ȚhE�(���F��I	
�9�q�F���{F����q���������A���;ʐZ�S�.0��y��5���2�F�l�p�5���7t�8�ڰ÷��+.�{�Q��u�I
%�5�1��� �{9W�3�� �y9�;��5��ƞ-�{x�l3B�����M��pSAǑ	y3ll���9�:�.oD�=�P����}�<�U�GTփ����������[��{>$*�(>J#��L��<�
ѓj�_R�v#`\���z�Ў�@�9v�����"xK�<q+��!����	�k� �X�eI\D�WO7r1<�YO�?�G��I���Vj��:���f̭��ڕ5���Q�{yr�3���#Wt٫u.��;�o� <{%��i��ӎ�8"��&�
Jݶ�������ֵ\�$ʥ(��'��|���B��{x���~��q�ކ&m,��4�-��L �3?���p�ֽSƧ���<社%�Z	]��Ŗ�=ʹS,n�>��f�����m!-��B�GԳ�Q�ٳ��x�]�I
� [(�+�'e�b��B������U�H�.X�4�����⡅��P�|8��3l��X���5�;�a^p����N	f�1Q��H����8S��� ə��R<�K�+�H���"��:�}*��{F�"�MQ׿VQ$5��)�����3�Q�Q��aa,�$��_��!��u��FHN����^���?yQ��?�_�O��� )ζ�Mׅ�t�[��3����	��:����gL�z6��/�1�lɻ�!�!����5��S�+Hgr�C.�Y]X��}P.WΣ�kx�c��v"�%���&����%�J6�%�����j���70���t2�  4��Ȇ ��U�f4�L�F�ڿ��3q/�p�˴�Z�zoF�.f��W�X�^&�Ę+���:sE3Ol��i����ʧ��pj����:�NU�ܳ�_��7�u�Z��l%��nA��R_�Q7R����U��5WD���lv�Uj����ש��$���7?6²22 9>�e,�ֆ�G�+���:�&���IB$x�(�v�^`]�x�!7#�+��^$<��(ș�|��Z��ƕ}ϽTDE��W����F˃<3ͩ��d�(��HLzO'S�"���d�0��{<1#9��1��/n�d��>�	ۮA#H;�g��Ο�\_\���0X�e�T�����b0��Ƚ��l��4|J.Cش��%�B=�/\��3��+���`��J�2��eԡ�N/�y0��*��Z/b�W��
%�s��r����g�l��m�j��C��{c�8�e7�vA��i��`Qb^��ܩ���ؔ�Q�~������r1�n��}^�9r�8�'�YY�V��ԅ褚 VuK�C:��z�z4�#sI���K[�V_S	r˓:&	�l��Xݥ�S���]Q.�������UC��8t�R��h5�L���cW�wc��x�Q=R��x�$��Y�2��D�o� ����u_�Z�H�"��V�r{WH<N
�$b.�k�U7b��e	MB��͈�j~w�ԳW�a�-%k�����
�����؏�%��@ܺ�]�QG�O�t5�=�G�
WǬ8��"@��V=�}ϸ�ǡ�`|��6B�V<u�'13����}5���Ib!��Vt�6��F��C���C +,q6%�s������f��>��s_T��'�/a�ʼ�h��^O��6������(�[(�&��sUu��ea�q����{�z���-i���=f���z+�G-B�Ϫo�U�O�>�K�fx�r�"RĎ�Ox7ϴ��K�4D���q����z���r�JT�֊�7=�ʼ3�Ň5����΂�PY3�>��D��ҡ
�x�:e�3pG�ܓ���)�~��D�W녀w��\�Ĕ�Ǡ� Qs;Vǲ��������Yb���\X�4�{�C���q#r��	P���٤���$Vd��x�����:2�#��`�e���=�q��a���q���K	/Y�W|��D�����`����oO�6�U�%�/_n�>�69����Q
bq�aҷ��5��в�mKU�����g�A+��p>�-IG����qe��)r�`]8:+�`d6��B$rC4�	>J�ft�@^m�N�F �����aR�c@+,���+k2X�jX9���\����iӜ ���\��\�$���e���]�,)��3`g�&_���}D�O1.��Qr�C-Zd����I��r&�P��PT��=`?W�	��^��]N�E��-w�[%W��;�M�N���N��Gl�`���� �]�`�(�	�k�f;Տෳ���dt����v{�t���1�����G*Fg�X[V��OO��~"x�w��+�D�{?�2Y-y'�5{���a<���s��Ť�07A�T.�Q�A��ȵ�(Ȋ�g�d5D��vK�I���o�n�ԨX�f��]�r�^�����8�UsMI�{(�����0fS��3!)�eV{k�l	��Dh��aZ$���}���e>��j�8O�,��Tdb���|�$Af��t�C��f�XJ*�t�����Tcs�(�KA	���w%)�S{�c���*�{��5=9��@]v�5�QW垕�"�$/t������?�rl�I��Ȑ�o���-~6�Ձ�E�&s�a�G�4�1@����7��in���bi���"��HOds�)���-�p��@���]N���ê#k�[�V^#f���WG�V��1�)�����;��(q���-�������Pёi�Bsg"��y���J��8Z�^�:T�{��40h��P��#�#�9P���뙭k� vg��Żw�M	�����ӷ�#��vM��f�B�~Ofβ ��hO`�e��g��`��~��=�X�2���A�����Xt�Y�gUx�Ǣ_(���@`���K6��mI:6�I����6�S��˶O�Nŝ��]?i��6+p��iSE#���s�q(}�3�JYrK��u#��
O����]�8���!�w�7W�w�c"Y9�(Q1)�foA�;�����4�D���_��|���;G+��U�d̒x�9;,C�� ���S��������|����3'4�G��I���y�xb�A�>�}�����x�<Y(���X4�$K9z�1�p����. ;pv^*�D鿋�bS% ���q��ıC���]T�S�f��G\��;1�������)}��̞��Զ���Yq����E��S|���W_��0Q���i�dki^���"��|��V��zIJ�K��O3�;$%C
[l����+>
��� mGC]}���"�) ^�a4UީO���q�~㻛3� ٟR�BWK q�f��h�|�;+*�d;�=1��h"�^
�\G�醀u!����t6vG��8;�	H2tyƔ���Q_�pW`�:�cVr}�m<�.�?���<7x7��rw�����e�*[�S��*���,|�Dm�±��І"�T�S1�K1ѹ/��u?j��!�f�P��W��{�.��9�y�4������l�c6Ҵ/p���s�(�Yx�!�p�O�ŏs��W�^���\�poߠ�o�Mc���_	�Tn�Z �b^-f�:���0M?s�A�����'��կROj5$6��3��E�E�Ը��4��?��΂�ϑ��x\8�Y��\Ü[d�N3rv�RSf~dn,�go.*蔨:�������Z�S��H���z	���	߰z7.�D�r�����e(���$0�D�|̹���ͅ�'��I�
)�1��|�"`R���nE�M̓�`���Eh������c��:exo�g��;k�T4(E���{���8�NxeH���<���,͝�(3�E�Jt{ס&̒9����1Ы�j�Ϥ��\v��E����"3���iPm���ݺ��	�\UÓ����J\��t�H�Zp��lP�����t����4�wٱ�y�q����I��N���"�#��RԚ��km����o�U���܁]i ������/nDM�mO��w4�I�u�5 C�EIPt"��Q�T��A(&5��/���j� q��'��Hr#:Y	��E~��a��B�Z����!'U֡�ZF3W�؍U�� ��3w�	W	��q)UZ=H�[g��{����N�A�:�v�� XC��Q�Y�P��2�;>�+@ɦ��hY6��f{k�vr}S���\�<Η�/�#�!̵����2�Ũ��#BcW�; �k�����=9uo^
��S`|�Gܢ�/6�D}b���'A��+�<dۚ@�V��Yk5������v�"�}���b�uf�
���Pm��^�(ia�M�/mԤ@��~]��qVZ0�)'&��"�+jGR�������~�M9ƅ�˯��'l晷G�s�N&��"?Ԥ�4  ���4�=���2��?&W��{����(��l8M���7�Us>!"�w�N��JE���gF��B�k�a[�E\ے;U���
@����,f� ���M��{O�f�&�;��6;~N��:���^��ê����t0����� y�%�ԉoD1��B9X�~��Jد�"���|<�#���5.?��weF
m�L���5<�ld�j��Y�����y$v.����xPg�!��^�yU�QҢy�-&�N�hW,�$]@XV���SC$�'�S��{��/-��d�h�MƖ���m.��Y����X���B���� �^*$9d� ��#5	`Յ^��@.�U>��1��|Yf��G~�1<YI��d�PG}�M�k���x_ڠ�eOcQ6ࡺ��+���=]�Z�\Y
��#�d���aޤ���w�S�L@�RC���RF'�ǿ��+A�^w�u���|���'kZx�k	x!^m֍mCу�^��~��So)�mx襤\P�u�_`��҉�K��\�u�$a�>�x�q��шq��-��~��d@۱�6�F�5�����](�����tv��N��H��֚0���@T=9M��ċѢ�Ɗ�K�&JZ�ݼ�d��rK���_%�&��=��+(�£[)�Z��WX9vW(߹$��)�f���/5���і6s�^��0@�u�b�R�I��Q3t���-�N�v��?�a`����<�p^I�1��(�$�"�*��N��},=vö�S�	o��m�-�]����:^��\�W�
H��t}����_���Jo��o[	"��v����ݜ��ʅ��yק@�.���gm�ÊVX��g| D�2U���#��B��XF��ܱ�D%������1�Y����i;2[�t�XP�<QA�cN��<��!���5Yલ�lxU�ºXJQc�n&y\$��s6(M�,/O׺�Jhwq /}sU�a�yJ����1����0hr�T�\jt�m��M��/�&�d ���prW���Y��Y��oi�x�a0�V��
��5ϖ�lF�^3�w7�2VWƏ��9�<�\��L12��a�(V�GXwcB���Z�7���n��L�: �)�BpF��5]w@��lɪi�=ρ>W0@��)ʊ���G����p�lɆ��0w_���\���^dZ���G`-���<{�B"x�8��%��*m��S�܊�A+��U@ه�k�f�-�z��魚u)�n_b�
 ��V���Mmin��+����7F(� �Ѩr��gd�e3[<U��C�t	�q0i~��//����OJ���S]i-��4�f�
K^��&.� \2� ��Tc�G�~��+�>���c#i���e�Fh7��:M�h��H���$!�+�H�`ɜ�~pz}ؔJ��@�ٻ���!���$���X��Z��O���ƢR�£)��wV��{�Ly���b����d��� Ͼj��'D��%�#���3Qb�ޒ%bt�����s��w���Ϯg�uco�9_"�n��sB���걘}�djt'��@d�Bf�ލ�=�N���3�Fj�8ȋ��"�h�y�$GB��:l�44�%Y�1'�&��`R�� [�+-�Lv�S6�s���������v�<�'�5�<>��X����sK�v���*��$�шw>鿩�4D��T�v�d����Mﾛ�5����C FQ�?Y"Y<�q�8b��压���ܿk��#5Gߌ��4��Ta4��?k-�G��^Kxq�%��)�И��� �?���z;0S`,%H��#⺛��SɅwՙ�@q;��V���9�̥=��\�FS����[Z.֖Oڂ5�1]�T�~������K�3�l���u䂃-;��2 T7�k(��!��ꐱ+2�l����K�xfkfrL�ל�u��[B�:����w����*~���)~�������R��JG�(��a�J��)z蒣�Lixpt�z|�ċ�3����Ar4� �U7)2�w�����f$]�����#�Ά�WF���g����*�'���D�X ���GxP<��L�7!1:��X�n����7��҅5{SEa�cנ�~��Z��z+XV̧4S[kc�=���^f.�O��(�(�M.��*��p��[�ZjX�qs�bV���|w\].(����v{����+!�`���s���N�i@b(���;�VeE�D�����LI���hz$���}��\.�`l��1�VJ$����^/E{�ш�P�)}�Z������_D��NVpY��-ȥM �U�b���x!U�a"l�f}��!�@~~��YqK,/��BC���4��r���]��&2����4�,�Nȿ��k�rY��e��<y�.q	m�u�]�����|���h�v#!stT���U?&S�@����An��?&S�f`覣|Uo�z5l�=5,��Ś;�x-dJ��J���4v>�ͅ|G�N�� ��0I��Ф&�&�h5����=��n�����F)�Vp���R.�q_�zJt*�����&�P���a��1�ه�ͭS��+\`���8���֕@��&�o�������r Zk�+��:�:&}P���]�f����I�o5x�g=��� �g�2�J ����̲Wy{���E@¿ʘc�$@J!'	6��jʳ� ϑd �:=��{�Kr��>���q���~���4��8�g���	k.�s�^��ILp�^�D��McD���cIuH[��?�]4�h�l�-���y3q�z%��������I��]S��թ^�u+��D{}��"���5��P#�<Bb��W*��g��n���7�N��� �.ع��u��+e��G[,��	T�~��y��v�Qc�W�r �@&���<��N��DzL8њ(�XKV��0rg���{���>>�H�{�lMI���%�t/\a�>�uz���*�"
�qh�6���Źf��iÂr>Q������:�����J�J���jP9�h��'G���� Ru�p��(�L}�$餎ȄN����?Hc�����O��6=^��/�؁��4^������}R��c,��ӂ�������!��w�z9Q:��u��3sE� �ȡj_*��WW`2G��H�*nH1��7ˮD�*Gˌ�ٞ
�7��5���U�C*��Q��h�C(��	m��5-�KP�	����`�Q�5���D<1N �(����pf��K�$�D�a�u�M�}�r�]���tFy�'7,r5^`�7�0	,{u ��~�P����g�E�W��#�a���G3p+�vO�5��y��Ԋ�	�S6D٢2Lo>�*K�{e'�e�-�������!�z�̾dyyK�2��hl���y l�a�ׁ�$Li/OkȚu��9�l�������WD�9jd��G�S�����ikg�i�qC]h�C:ϳ*� ���k�C�ߟ����xH=E4݇�K�߁�P_��#&9�RJk���64�Nc�z�^��f���u#KJ�@��&P��#��E����I�zu�N	��VNdt�wn-|�:�Ĥ�}L<�7o�n���iw�w9��t͞S<e[>�
��mI�ct 5p
qhd(�VQ��4J6�曏RŽ	�� ��$ހY&6�;a�6����-��=�zw՗�:��D���GI'�.���=rA@���)�Xu�ʻ���6ʽ����|%��,�Y5��1()df����)�	��PՏki� � S�E ���l iF!u��(-��(Y��|W{y��ֹ]T�����
�T�r3}�ܨ	y�d��c4f]e^ö�i �+Q���~?p�������Z�Uz�_���W)�/|i���(qOn���ƾ�aD�;��
 �5��P�;��0|�GF �H�1L;���|E�ER����+Õ��Bq�g�r��r4��ŉ�g@����dSY�uJ�^��U8��/�d:��3M}�)9,R$U�j�,8���/�s\�{�a!�s]�2��򸪽7dFj��ӄ�r��#.Wt��f�[����IXQ�b�Q�+6��g��617���	����xo�E�6 �~��~]\��,�.uI��C�TjL��c�yi�p�ĵ_W�����)�I�1�{A {��`�jR��Xݻh���!x���	�>��׆n��S�<�$7�uY���Zn4¹pz"���d��o3�Y��⃉f����[t�n�� *�'/�7�h-����o���Lג���I�p�#7Ʉ�T�ʥ�%>�M���)�� ��C�Y�K ��V�O'դĝ�v�̏�$!־�X�H�M�d(uC�0#�o��$���$=:�����_I�z�)i��D�T.��됿Yx�j�iXHn�4�����;+��F��_%�rK�S8�N݋��#�2�����_Й��2i S��r��o����MS1U���J�,�7��O�H�v���J�4teM�⡢�q��dfn�2�'���D�ۙ��
U�հ����E�|�&��Y��wݮ���z}�6Q����(h�,J>6h �Gd	%Ca)�?뾺�����yV>��22��~@R��b1�sx��qu�_�~a�4�Y qȦ�'߹;\ܞ�B��g�N* �C�ʐBy;Ã�؉�C\8�i<��b��m�$���z:����� ���^���]�����,����L��?k�\'��R욬���+L����B]�� ��;B��p�kA,�*/�j�N!V�Cr>Uw��׏�T���h��󮺙F�^�{�WR:�C�ZS���2M���M������:�����{�T�d&��d�9Ɔj����"�Na��s�d>�����a��b���'DX��Fd�.�+~�G�>������d��9��z!�u���=�4y�9����nKHK�^w���{ů�Y�����aSh,��7�!1��g�	xHY������ȝ�VNc�yw�t��V����J��\s�;Nb>�G}��D��A<�f֒�m��a�Cǀ�Ǽi"7�o~5Ҟ��/�1�߶���@q�ђJb*gjX����)=cX��H>�O󵈐0�,(���X�i��Ow�8t�E�GQc�x������f���ϸx���U��^F7G�F�l�*|J���&�	"�C��0כ�o�w-�Jr��
�t�v��caM;���U�<q79C�g )���͵fSЙ����%��׺��S�KH��/U����m&F�"�ba�Y������/��8��Sɘ=�H��T�߬߇Ѣ�o�M3��LLܾ;'�j+8�1�%�u	>�Q�Qw�z2�A�����?p���Y\t�[r�D�ΔS��!u���u�\ ����Z��o�_b�^Ų�H=���˨e4�km����)�5$nm�sg�`5��Hw�f'��4���ZoH��!8�.���4�� %	/�S▷��8��N㌁�4Z���%�2��Z 
�����,u|���?%�g����������@1fe\h���!�//�/�6�#ۓ�Ar߉s�1cŌ1��k%����0x�:�ı~����$����G���IU�seȺjK������hW#��\�����]f ��]�t@��"w��m����Z�����͕��@=.Y(µ��Lf�¼E[N9�æ�j���~�/�	�O.����i=Tn8�YM��얠�����݋�NP��E(n&�0c������u>�����&Z����Na%�0Ũ�����!b�H5�ѪS�nW^���֍������N>�_$z^�4Ԙ�Rd���Ă�S~z��>	��O�7�I����.�A=N��;�����R�&��{l����"�D��[�/[&3�l�����Dc�V�����w��#
{ߨY˳潹�E�����2-k\TƑ��P8~��Z��ZzHXJ�~�*{)w��T��A���y����rN}q�����(Q"��ާMyx���q��1�0Ҟt���8��fj[{�zV��(�8��#4XhF����z��9f��y����8��M��k���+=1R��ɓQIU2��B]�326_}젂�`u����è�[`,�-�Wd|��0$�'G�Y�����D|,q��Q 0{ԭ�pTސ҅��'u��H��=���=.�4}��-�~�Ƀ�>�6Q�Ϟ�:��YPlFp6�Ly��ƼVUKn���o:[�3�j/�~D^��07�id M�����[�ѭ@Q�H)���]��p�Q���G���I��V�������;$����E���yurIlM �V]�]����R��RQ�M�`�/�X2�o������n��:o��p5 ����'V���,��u�$�!�l��@? #cgo�sX�ˉ~�Tt=~�S[�+<�J�sP��dT����gL'FgI�������E�1h@W��*@����!�����~��ґ��A�|xp���z	�&�w܂3psPP��\�u��X��(��6�;�9� wT�E�Z��L��zF�}^����pmQ=\G�'�)['��m� 'ώ�h�K�ߎ!�6�,��m�IUF�oA�����T@[��cA�/3��O^?���Vب���5��{!n�!��M�M��E��&��^��@�<���W��fKgL% �;(�.���W�<�/�1��&�� �V��+�!��8��u�QA���YL�nt���C�^]dJH�g0�V�F�cj�����m�y�,���H��q�������J�����n�nK�8A�n:F0��C���K&���d˲�z�3�P
�Gy_�h��(<;&Tz~;���޵!m�1l�������z<=r���y�ئE�w�<���K{�(0��.Ѥ�t��ҾBj�}{�i7# ��p�^2���J�@!���=���犍I$�H1	�C��u6���hHC�j�>3i�=�c�8C�=�LX�K�u�*B�Ì'<���TF�6El���
e��[��n?�5���4��'�<��"Q��U��5��e�5%>���J��}f��[E�|O.��b&��c������4~�8�g�Ǽhi�#W���W����$D�96��WJGbD��+�ke��������W[X�[��n͒IC_΅�����m��Ǣ��o���Eߪ�{�M�L伨�?�n/���A�F�sT����U�;�b�:�fɳ�#Y�rLO��H1C��$�[
ͬ���R�����|�jVK�nlǄ�i��/�։��-w^$Z��BA�z�N���������M\�)�pbՄ��c1C*$��BY6������L�ٵ!�`
r���J�T�G��}����4C�o�ϱ�e��3j�9MUL��-G�Y��|xQz�:e��'��%4�=դ�A�6��V
�\��`9����/5m�5�nk���w����RϾX�8���A�yg���:6�rrѮ���2ZU8.� ߓ0�Qc%?>�?� g��[���I-C�Ic��~h3J(W(M$�O|���M�]�'ء蠵�/	�϶J
�3n
�J�o���zp�yS�0na'RUf��8ӽ�a�ǀ���p�N��>G���1�FH8�󱽥���d�k�o�fת���&�}o(�X���x�ېS�I?c�2�4�nV�
cw<a.̓$��?(����|�M�.)���8n�7<gd�(��7&����ϭ��ݳP��@�JXd)�ji�wv|��(�<Q���#��2��a�^�>�=!�I�n�}�����KsXW*�;k�Sc�XP'���D�G�,�l��<��/Q�ik��R��-�
���mT�S�p8΀��;u-����A3'׶`3���j���Oo���t�rd�
�b�ƾ[���hb|=鳆*��Pmz����Br�����WN���Π@al>-�����:{[n����G���E��f͕���8��2�@$@7�|(�R�PA�ڮ
J��Am�"�,'���2	M�H�!�'�Q�{ҖH�ЋR����I~�m\��"��a�]-�g[Yؠ��2Լt�ƦFH�(�C����A�k�l�?&�k�i�읫1������w�:vv4X<~uЕ���
��^o
b�]Q�ꯛ�;����a|�%x="�����/�}**�3$��P��*�HEǴ,���ҝ��)ސU깗��E�+J�;oXd�P�V�)����Gng^D��p�E)O���_�R1W��(�~YơK^�s��t���塥���%�b�����PqF5�$GI� �1&&��]P�$G	'��voГ�@��ʍ��Q�d�Zjy�����j3��ۏ�w�������	�p<���BR�$�
{c��[\Q"t����5$&�݇��
A\ְ����n�I}���l��O���C08:㲀=���R�����75GnZ�[8��4z[�"G���~��>���e��]x츟�Ņ��){'�?Qn������i�6)��I	�Z���y2�Lޘ�ȭۿ��[��+�
g�zN!��zrJ{�D�ѣ���������rU���q1
���pO޷jTC�z"��{��	?&jp�5kՂ&�����^�c���	6�B�k1� ��4�HA뚬���%b3SGa2��"�}\�"����R��K@���S���DG,���ў'�lK��|`�h���#�'����a�'���9��u��O�8�w8�:&X���xQ �V^�OSI4û��kwNq��]��j�:�Ԙ�G̵o�I6ئ��'#8��ٷ��\��)�:�K?�S�[��Ei��TX�ȅRţȪH
k87�w(sE1B��
m���x�oa��|ԅ���5�Ww[��,AB���lN$���eX3��!²BN����T�6��#�����cN�k^����!g�Ƅ�	S��|tj��*��/o�]��F�a��Qşw��@��ّ�C�N��B{��r��iKm�Dgd�vs�"	S(Q0���-Wf�v_L%���/�)��	B����7�{ ���̰Zu�m��|���Ȧv��tϓ���������b��vb�SC�0������i>�G�)�Y*���ӊ��.�L�F)ؙP�!swm���w8��Ϫ���aㄫrU5���C|�u��������3
��ʐ`MЛ�4�v1�3Cjncm8���l�N/�S��ŧ_kߋXG	�?�XL�����h���`�a��M�ϧ�(7��X�ꨦ���c��j�s���]��0�%Q$-����G�]� 
(�%������c�mt���B�4ϫ���Lq��� ���62�&S!��֙���.�~���T�4��E3��_����,�eA���s��VY����?R�3�Q`�L��C�܇�^M����u]�g%f^ݝA2�mo3'O%}8��KR�a�1�	�Z���(��^�b���w�j��/U��Y�C�W�1�E[�g ���|Bs�7�&�݅R�-D�3�a���:�8ÈV��"Έ[qy^ǡ�zC���5�%sy%��Hk�y+r��'O�����,��_�$��  �>]�EC�@�0h��s1��I�0����72;㧮��*`n��d�d��+NPd�/{T;y%<��Ɯ�T�X!�>Y֣9C�J���u�ٱ_r��&�WS��Oq�N��"ˍ|������=�JD��y.��!�S��G}����\F�9HD�n@	|������r����vv���G�e�Ai�͟Xm	Q��˒M�`އb�3L������ �-`/�H�z�Ĳ��k��ZT㪧��D\3R)<��ְ�̂k��?��}������9\I\*�h�f"a�d�&��ڷO�i�&��ld[� ��68\�����(IC�sI)lG+2�.�Sp�z����!�tƑ'V�5���1��d0}�0ǯbL~���o�6˕�[�,�V�u-��y<f�}4=�~�-/J{�9�l��۞^I�#��n�'/���x��''$�5˒�>)O�� U�4�q��O��)Y*�sX�,+x�5���H�)`��堊�Q��&���Y_����1BZ N~y�LѦ�lJ�j�T-ɻ���@���
����;�>�j�&t����u����<#~�4
���?���W�ZP�W�^.y�nU@~�l|�yP�'؋���O�e�)��D3�^��T�B0�y�)#`���*����Q
���Ooh3�Z�kO�.�А��)�&Q�l���
D����W#%N�\L�N��~�u�2C�?�J5{�$U l/�Z;���<�z<  ��Q�խ�b��$(~�t�����#���d]$P�]T�OqEmy����Ԧ�s+�9m����Ρ{46[�����B)�T�%���xb@Xo���&`�1�*Χ��Ȫ'�+�8���\.�KW��5�t�ܾ��IW�SгE��?~�Fkΰ��|��·��z&2x �]G\�i��������v�uL{�x���!�)[�,8-|�^�%� E[e����軳H�D��M=y����6�"	�fx��\�s�ի�O̾��3rX����PlX�w��
^����n�����9�<�h�@1��ҘI��D�у�O�OHr���Wr����}�qUS%a��pT����OD����PXB���9�|t��m��-;�d��W�e2��@�@v�,׌�S��U������,��ow�Ԃ=��J ���s�B���Kͨ,�f�co3���r������ɿi��- c=�>��x�����z=�S1M���L|i=4��$�$��3I�[�G����{�N�7n�83�zt8�*r�;r+�W�[�0<��}e!���)Z����� }삣�����p��F�z(f `a�%��uFK�l}�<�q	�j���絰h�p�� ��D��7Oge��b;u�Xc�V�<b�E}�A�Bn�����|&�}�T/?vo�}w���(NT�����Pf�b������)0�D[}`���\�w6D����yF�D��U�:��q�rs<��B�js��d7i�K�!E�c˰6�Y���	����v	I�B�?3�ʸ9��@��*�P��Kek�߼�*%Y
as�d��I�a��C�i-5��=˨~�#�N+u'���@�!G�%�g�"LR�"6?ߪKy�nύKB��~qL�[_��[�j�Y;�ӫ��HIR� ������4��A��2O2Q6��Y��l���76Y�~OQ���u��N�k�{�+�Z�4�����9�g��Կ�:��.���9��'�&h�5�4i֫�~�����^��Kԏk�h��|.�`�8�_��?ע�M-�T�ӓπ,�n֔������8y]]�Kr��#�z6�W���V�=VuhQ�(��o�jUh��M��ר������x,�oc���k��O��77p>�T� 'X�w���"i��>w+�����o����i�(�L�����$l�������mc,�@@Eu��?B�x���0 ����b�v�E��3��}�ͯ �f��EDˀ����p��k;�M��+��B�u!\�L�;���<���������#7��z��/�M,x5����a]�C�=���4�Q؁3�s���($!�����%�;�J����L0�:���%�ʟk��]k��l��x�?�/N8u�̏����[�ć*و/5�Dη)�k1ʄ��۝�]�ë���.�ie�}4T�6ٮ�:��p�������K��kX���"G��J���e�����S0D�~�WN����.��Qgk�t�w���HxC-���������?�5�^۟$ES{1��?�o����0��@������� �̶04i���A��<���>�PMm}��u���C<j�����G��a{�/�&��Ң�n��_�(-]��hoF�=���>��f��9�ֆ$�/�U�C��F�p�9Q������_��hE����U��W�\A�f�jZ�bb������Ӓ�d�����/9��t���1]��I?���Wi��i���3GIL������\j[o�"��V�z.?�Q�ʊ,��Mc��Q3�u�ʎ��X`�Ap(a�iC�Z ���OC�����o���&��p{dB�:��:�pf/Y��5��ܨ�8�n;)m02`��S�7�Sf���W/i��m��ygth-�.�)�TjYZ`C��u��`���LQ�mlO��X�ׇ�U�u�����Q���3�(�l�N9V�����@T�g��k��ዝӽ���{u�#Ɨ�����gWs� 1�-�B�/\S֢Q��A�I�s|ǌ��"��:(Y���[�`��_�t�Hii�<m�DAx�W�B�o-SeV��ܵ�q���������p��qʼ��U�'X���Kd�+HDg|�D��� ��63υ!�|,N�=>d��ֹ5S���_eڇ悱e�.gD$���͇�Чt�"�j��>|����NAʣ��� �D_��<���ʛCH�-M���H��k���p���X0��m;��!0%S�x9
�&�j
���A�bݐ(�@;��ԩ�rH�W*s� ��8�z���G���?����Y�j��gC�1�~��Hmՙ��J��ftw�)Ӽ���3�C�g�I���CyR���z9����9��w��Y�߃�9[6cʧx]<)P�yt��c�<(�R�3�a��-B��0��)Lb�@�"��� ��fK����8�En��ٲz6����['̮��>����������_^3K����@��'���~EK`H�4wR��q���Q���\��u+��8�$*`�����VG4~b��(.X����Э���bxy����:F�K�۴�����l��~��CE 	P��^�Kz�)W_[_yy�E	�O��כy[x����M2��s(*�c�N{�\����2(��	�ڞ��Vϝط=Y�o�xy��	�t�G¸��Pv�E%w턜j0���c��p%*`�P���2~7���J��q�(Ψ(��d��	�ވAr>�^�[sE��a�����|O)ӑ�mV#p7̽Ҝ]v�@�둨{&GD���E4��.`!{���=!���,�Ո_��3 ]��@5�>�Y��.�TC%��LT���
=X�a�jf��x{�y�Q�Dqb�����׮�͜ ��~v�i��Q���,�����qv��yi��WI�Tý�+�T���ĥ��()z�=���R�e�N�a�iSU����8zǚڋlHt)g%�s�s�.ͨFH8���yk�`�/�q8 �?�(Z�=�kԍ%*�m▸�H
�REq��;2{���6j����?� �`/�s�c�lJīg����ڔ
N��u����k�{�#V���Y�U�����Ⱦ �xc"wKf�b��e:~5~o34�Dev[�Ǭ%E�WPDp���0�/����\���0Z�B��O!�ٰ�}��V���UQN[�؏����_���o��Oυ��5C�va�)M�	���O9�k�DP*���,������#��وS�F{�	5��@�K곥���5/��i�}vi��]t rO��R�WjDi�Z��O�b��-��qd��]�)��M]Z�����M/7	|M9x�fz�fzG�Sٸ�aY*�L�WT�T���x߸���v�>����cڒ5~^[�a0�,l+�����;�Mo���,Q��;�d0�$C��� �RS?
���"�FKd��_x�o��"���Yo:���|��kT��?`�����W'��<���w>��V#�];�����j���d���# L��b/_�#���N]uo�)�� V��Kr;C�������M|yO�_5�Ω6}��ʘ��W[�:́�B: �C9_���ت-l�:��9��v|QC�m`z���5UHk)h�+g��s�o�����&��Z���vd�N&���,c
�ي-�����0�Cr�&[:?�%�� ��5O�4� ���㰚?��V�5���!��>M���U(.;q�N%w��!�I�ox_��H
"�F��H*.�Jkـ%�ø7-�L��W1���MR��8(;l�g����K�5��ua�8��������oǴ��5/��� �=���?hO%\�;3��܆?����M���U/ ��EА fی摽+pT�;i��V�����1�%�r��zF����l���MJU��DG� :�)
)!�Y�y.4;�>ܧ�C��J�b�$�����_���������5�HI��>"��g�Pܜ&����E9^�XFׇ��!��z�u�Ωm�tׄN3!\P�����լ�0A�1�9�޽�_��S�D�@b��Rʟ�;�ǧ��*X#�����]�xT��F%��CVf�N:[)����@7��~��L��ʴ遇�TEp^��Ü��,�a#�׼��Ō��a���C�3�	f�ɶ�B[>c�9�	i��?SBnSfA�>���ٹ��(fF�xe�,�4�{Z�u-"��ӹobS��@|��Q�X�9�Ѵ�v�w��	AG�H�E.�%Z�o׳^A2�,R
�D�-J�t!إa�l��#�Dx9�̬M�6��\�}"���"y���`�$�v����ّ��*�!!Bp������J��t�H�8փU���aCiɹY��v�axO%:���O#򁛔,���sv6��l�6�K�*�n���m�^�l�=~:��`�[��|'^�L��ΐ?)��ML�w@�$��!�D��
D>��X.���46?��	`k�����$k�o���