��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jåا{�\�u�?߷�dn@6�zf��r������;$VF�w��O�a��w����m�f�LG(�f�3�*���w̘�{V�i��5�\�R�׻r��'���4�O��m x뗐�8��=����=4��b�X�d5[Q%[�ç2
Ő`ôa���=���� ����w�Ħʹ�;M���)=EQHٵS�1�R�5�\����'�D�!�9+u*�H�V��i�m���Un �B��W�!#���%��4[����*s+�;���B�OƘ�B�4��/�����kW���);�S�l��sG�C�ے@Ce���<�q�CTW�>I��a�������F�Z �M8�`i�ó�V5B��*��e�G�D8�TE~��iN���ߞBd^7]-�
�C~���@��9ޝ������f�"����R�G���AGN�x�O�4�"�ydIY�NrXS5д���+�(J�/:��~�ֽ��4�$�[�?Pa��"�Rp~�)i���藀w�+AB��wq�2�K�Cn7�$?]����`/��R���D�:&\}�0����f�2�R����z23�����;�������h�yb�yE�/L��%v,���^���p���d�<?��*GYc�[�`�_l�d�oF����N9 �B4?��ߖ;�J��OF�,��nFw�8������|L�UltW����&�2x���.H#]<��!ڰ�
�Z]����0ܵ�z(w�ߑ��r$W����G@]����y�i�E�w���:l[��c9��/����˕p�4rֹ^��x�Z����r�
� �, �/�E�����?�Q,3�C5-���}����_b^�Gm� b
Ve���'وJ��u�&΀9Mb;/��'W���a�-�q?G�^���������fbF�	��!�#�=d�Ok�7���#�;��C�\� T�O*���V7s�%�.�����7Z��@D5��\Aɧ$�I ���~���c��&&�第|u��뜪[��VT0���~��	,:?S�RW�ȹ	�R�4 {���'�b�k(��ƨf`&nX	�1Ғ0�SPb/�������ʶ`:y�?�����"D��d��^�%ʘ�]~o;_Z���4�Rݨ�b D=���1b�n�B	;��t�C�@�"���/�F�/�Φ��|Q{ӽ
+?|,Xg�N^ʹ���Od3c��~fi�IQ�>��T�pM�PQ?���S�q��Y���*Y�_?�Ĩ�Yi�|Ty	��PkK�a���3n�Z{�����{��K{�UJ1���W�΀�T�F���j�{_��y��ʹH�|��ӛ�,:;�\M�JM�u��/s �0�?�f����x4Y������v^s���ݯ}��믯�E���t_?�W�pn�H-8�г!_
\h�7 f�*^C�r�!B���t]3��fQ��� |ѥCRU���G���{5H�	��Y�}���-#��n���8��u�k���G�C��r�{�?����%Z�p�]���s�FVֺ��('�v_����ܗ4���K�'e\Z'=���#0TM8v�$e�ĸ�