��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e����d���f{��@����S��>���4{��ת�AO�Q{���X��F}|6�Nw c1G��_�/�&nʨY��q�D��<)��qj�RB��d,	1�1����t��ީ9K�JX{R-3��6Ⴟ� �~�eäT��B d�y�5Sp���\�����|�z3z��'��lR^����F?\*d��r��7 ��`������o�oZ��<U_��H]"�n)�S��)�Ӏ������Oc���� ��^���K]v�����e��f�!}�7�v��>��kf��*F�3���Ց���f3��Fq[+��$�QCZ/ziB�p�t F�/I�I4��(D�_KV�i7a-�<X� V��G\2���Z��!Ϊ�Gl�)�_�+~i��J?"���g7>����>w�:�x���f�jZ��T�ēcjqU6�l3�t��]�b�A���)�a�Ϫ��>����b���Z��y�et����'^I}����*�/;/�*@m� Eg\ʠ��.c׀7f���)H�̡�m�&Iy�0��H`�� 5�����|�r���:�Ƣ]A��\Y��HG�WV�/P�{�]��죞��ͨe>�.�(���������	d��h�Z��r�ɟ�S�����r?z<���m���%�^��*���h�^���:�̘�[GNpO�!@�K���Ud[�(��QyPz��������F3�`V�2fvc��!�g&+G;��(0m�W����ЖO��sw���+�\���l�����G��{;!���!q�U�K�X�^B:@cݪk`�&l�3�Ь�%�r����';�F� ����C���@�N@�_-,��c溼�G��� ���"����x���s( �h�X��S':��}�dj?^�����"!��7bZVky��K���(���^Ήr-{�k��q?(��ߢ�\�Ι�5)�ж�j�/�����"�q��UD��%=7���JU������E�Qq�Tm���ynǉmk!�҈���1�P?[t1�W����^|#Ђ���N0���`%h���bzp4Ĵfص��$8m�4v��c'o���T�|��g��U�4���$��B�$n�:�k��ܣ|n��A��o{W���ãEDY_�!ӕ�m2���>��_jbe!vb̙��/3$�q�����Zq��1rʖ@Ow�]�f�l������ɱ���:AJ������y_S0��f�q����9����xG��B�H����;�	�)��^C ��!�V�1y85S;�?46�U�Zޤ���]a�!]�����]U�
{���ulG_�d�dJҢ?��H���+w�չ?�|��OD�ςۭ'��HdM�N�JU��$�'pDY=(�m-�p��0�%�"�i������s�sH0���eWG����~�����I����N�ca)̑�l�_�i�1��N#�T(^�S�5��v���M��r��NL����.�ø��\���٤�+��FH/�*�>�H8/�K78�	��EG�-�ZJ4c�� ��TѸ	d+��o�w65D*�KZ��Īc\0;РD���{#�8��"18t�{w�VƀvgC��t|��a�dhR�)��7�ʿ]�Nm#b�����E_�5���.�>#��_?�k��W��c��]*.�L�k��m�T䵖��V���ǉ��c�rQ�1��/붴�e<�Z���6s.Ll�e,Z�ڼ���D��Q�Xl�������)*B������c#y^@G����WX��U�����'Ǉ�2>� b���|�e�W���q_IxbP>�Byn@uG)������Ye�ʹ$x���~>��;��b����
���+�i�'_@j�ȁ��eU6���M�*#Gj���(zr�7��3���zD֦��
��G��/�8�ċա$�����?��m�f���Ы��9Z��l��`�'�̳�'��ݢ���}`gw���Mf���,�kx	����?�dq�A��(BN���ύ���-n����O���L���:�B[g9�YP-��Lp3���S�/��U��w��Z��}v�Ȉ�3RV�,�@oH���ߞY�O�#��uX�b��RA�Uρ�!�.$����;�e@��=�}��︳[�K,�5a\�wş�RI��"Q:���+9���ߗ��;Q�ȴdy�Ӯ��<C��5� u�{:<�]*P^��y�>�� /J���'�5�~JM6�nXW[u�pAև$p���k1p@��z���gy�L�ʷ���}S���
���<%	m���5���ԁ�|�|(�'̣S�g�Jj�P��* y,{O��XڌL���/��:N|��n��m��<�>IMB�ԏ�L���6};:۝�zS	ʾO��Y�uoF�.]`!e���NV�z �u��˻��|z�G"c/�:���+�,�������I����W��H��mF��)G2X�f�ؙ���ͪP~,���v���wzX�\C�2)�����F��8\"���߱��]eFw��
	E���nў�Geh��e��E������!�;�J���l��I)]}�%�q�fƲUx��^���+0*����T�{��K�ert� �4D�56^�W������ �5$vw�C����s���8��(���'�%@���w�W�]�܎V���,^����U�C�:�Piy�mǪ��H�V��pG�X�v�%Uy� ��<k'Z4�f1��34�9���x�dM��r�L�+La���A��_����ę)��`�&�{-��'���N��zrGi~�k����gD s(������M�I��&�%��9����L'cY3)y�^�\�#��FTN��בߣ���x���w`Z=���A����I�dfj�I����B�Q�͌�A�.55�N,:�����W���U�|%'�o�L#-��!�Es̙08޻Ø�����t�D@�5�[o�N�,��"��\��Y�H�4���{�]]V�1��1}���L����n��A�C��9��(9�t�k"�hnC�N�0ۗ+|�G�X�¼��y�ݤVjD����B@v���;A=X��ˀ�@TKK(d�� #�b��>�갥�!4kD$��~���Q�p%��OD���3��A��v@:j��6����ڃx`�p���ֹ3Y�Q�!��'�~�C�-cy/��)�4�:�igy'�Ұ<*�l�T�n��n���D�]¼K8-}��Ee!�؂Ǹ�Ec��BD��_�� {���nx���)<��B�XL^<t?�:(�����Zw�ԑۼ��7���K���P5���|�Ŷ՚?7d��h��ME�S��j-�ЋtTb&'+��w��3���P�o��Q:�۳���WԝL#��37԰�<��S{��žK,�ܖ����e�o��a��E�?�@>^4�i(d��o��^�g��DYO���)gs}�<�s"��s\ګ�+�q��*X�b�:�n���O��%��a�Qh�'� +��������ם�>v�����I�F݋e5*=�wH�6�ҝ8�дN�������;��J�<�b��l�݋�wDu!�Nw�q��iV�z^�|��"�@���	%�:����W�gi�Dވ�Pw��Q(H�� Z�n�w�qi�������H�|e��`D_sÒ�nŮ�S�p6(�mٴ�0?eoGQE[�f����/"���΁������X?J��p[��.)H�X;Q�E�.:@�Q�b�g���7LF��u�Tk㏨���ʾ��,���Vl�xgB1�7�ȿI��P*���ePei���i�IǸ�>[��Ϻi�{�C�E�jo9���nj� �)XL4�Oi1�Ó�����7d�"ʁ��G|m����9	H�\�+��þ�{<jN���N�[�ԎbaEg����p9��Ɲ�\�`��.�+��\$��ō�^,hYo�sc��i��P�/�
���LC1t�9�E3�$ɸ؁>=m��Ŀ��;?� �\���������^���'��( ��ɒ�d:p�d$-P�ٕ��D�6�̪�䡅�n\*)O�&��
vd��1l�LA��8 ���|��cit�a<x0�1�b�(����E��B	{ȸ
����x���I�*���HN��ƛl{�	�@�hb�S��b����!�X�%v���/�f\-�6&�ͪe���R�b"�^%Od���5��wԿa�{���t����{�?+�̅���U�
��	��ݻ_>g�0��7��9��fUv��x]\�O�l���5�u�걾�0J���:���2��c�]�׳9�_f<����A��4,�����.ːu��@��4��Xn�'�IS`%
εb�Q:�?�0tN8�\��6�@�<�cT����N���W/�$Z�Jgl���WZg�Nsՙd�@Bi9��Ŕu�%LX`��x�8�;5J{��bp�ROM���%͝� F���'��BtolX�6��U�CP�H<�T�Af�B	��S>�3�����}�o�f�E�Ш�]`�qF~T��7�
 }��v�$I�ᙚ�>�<�9@�f�4�o/�Xlb'8HI�}�Zw�(���8��'�P �!@ө}=��M��dI�t��F
��(|u�C���O0��ԩ������v=�A ��[��䇪����2VYG�h��ͯy=�Vt�f��<S��:�e����\�?N���B/l�Io�ϟ�,m�l�'��Κ�����F�u�_o֬3뉼�gG��9{aU�r�b���Y����r/�x)A`7Խ��lh`I��\�g�J�9b.Sw�@�����v|z����j0�]-:R���1���]�/55䁦�Ë������!4���ň��EC%�B>���r�����7��6(!�3'��xJ
�W$4Ne�0��Hav�lFL��
R��5�ߘ�5ؘ���>�N�2����lj1!�+�S�Wtq]3O���<��V'�B2�y��`��3=�4޳�-7/%�BvY�>W 	�D�H���ft���M�̄�w��P��tp��~�ۃ({�ѿ3�f��e��H�6]�{W%��v�BĄ�3���H4�n�=���r�J5_Y=*SE�RIM��7����Yc��N���� �bí��P�=�Z{&��S��%iy;�"��Kz4��p���G�X������u��;eiQ�{_.'��2��@˼��?¸��#�[��&+����C�(�يH`9;���?1K��/�vr;ѽ��~��!u43�Qɷ&�L���u�~�`��n�(����[!b�~��W�f華����8N��&�"�Ql� ����w�j����}�����bO�XU��?U����J�3a���hF�����:���Or�w��� ���5�>�zi\O�-��[�{���%�qz���i(��8HLKר��4d�n�jF��f��yF6aM��.�AʟМJ� �L�E4/s\�B��`=i�]�H4���s���)4�}DIQ�3N�`�5����ì��D6+��(R��(�<����v�\�ڬ�W�����*�uJ��a�q��q>U@�/���t������`>1�Oqo�5�߂�ٱQF�=�4��T��ށ�7ޜ�ڽ�.&�M����v`JVitS+�柜.P��Ė�ա�S�C�x�إ?�D��83^t�'/��?)=9KIø��~�rj�7�P=eL؟�Tf�� �8���%��9UHZc��_+��GQ���_v�����d�7Kr5��̓�~T%��5Stȇ�܀����3f�6��ƭ��G}w���Dq�:�7[�n,v�y�ݬ<<��L��_d�R�1e�:��odۯ·?��T���爃tP&#�I�nG����mR���h�fr�hm*[M#�U:"�ˤ�o��Gy�2U��!4��Q����;����9���]��y���k%a�`]�x�ZS˲nɵɆ3�����2[�SEp"3U��$l�%	���gU�ߑ��~H)jJԘ-
� /pW�|�Y"fI3W�y{j> �gr1��St�>~��$vN��p��5�&�J4}w�vF�'�p
J��ʂ�Q��w]X�2�+!з��=���������L+1���Q4�9z�m ��/�����K�J�#�>t��dWY��:YԻti��
���)K��e[P�z�i@��������2|U����(./�m�Յ���8d���e� km|]� �͡�Ŏ"�WUpS�0.��W!����3^e��j��WR���(�x��+<T[{�E��ф��������G�W�����e̩�<Jm�x8��&I����t�>��,A�\w��
�W��c���,�\ӽ$&c�
��T�����]�b.�:!�����"a_�RE~��<���w&ݶ^��5_�G�U�����p��/s��^(-���8pnr�`y*Z�un�1��G`xB�D�?%9�)jo�q�q� y|�>��yw~AP��$�n"a���B�����΢̃`�t��<}G�3����Ìb��4"�ghL�I$|�lH���h�3��b`	���mV����[�4Jv�ą�8҈J�����%�ZK����F �")]�O��Џ�hO Ҏ8h��%�q?�"y�[D)n8rH�ű��*��jb]g��4��V��MQ_*��(;�w���򴳲����>�p��r�.�]s@��gJ�7��D�mI���mX�ߕ�?ba�{u<�M�5U(f�E{��웬� 76�R�7#֕�&�I�N�o����2&����=�@������eKn�U0���j�E�*�$�H�%�=x�=�k��s��Qd_m�eh��FmEڱ���5Ƥ����Y<R^�O1��U^�?#�K`պ�Q2`��o�h����a��|�s��ɓl�D��v*������W�LŽk%y��lZ?��UA���d�*��[:j�U?�Fv�q��K�Q�/_;��EZ���t�>��mmdP���ZR�qK�
����(�!n��~$*�f�A�f�1�%�� �l��$�-�=�q�ieu��T��@�Y��Z�B俷�����`W2�.���:�8GU�dA�!9�� )2�z얚o�%i�������'4M �����Z@0���;�0;g��Y&�xSx�Q"�D�G�G|8Lһ�I�x!����~��Ҫ�}o1*�2�	��D�fH��r`h,��K���[B�����I+��Dۣ:p*��:Ͽc]��*�'"X滩�F<��׎��F-f�99@����/�����>�0�`_/X��M�u��ֻ�.!�@����}�c�,�e�"��-����
�����G�F�z�ۓF�C������}��r)O��R�kj�L�9%����*qwͻ<9��{Tl���	Q�V�H��骚�X�Ou��l$;T1�5	�)D��]Qe�4�����(����CN̮�^��t�[�@��z9�{TZ$V�΁�b��ٽ�؇��[w�لP�8W����G]���m��'����z�fp�h�˅IY}b��0�W7D���TE�)�K����ȍ��F���U�����F����N�dP���<�`4���n\��?^W��ԡ/����۟�2��qY/�^����tZR̿��A�)]��sB�l���L�Z�_� .a���*�,x��Dc~�b7QyH��C����
�����C=����Gl�8�a�7Tل�����K�֗�[�ׯ�f�T��4����7��vqOśf3��D>���M��v	������_5�2|�"6ȐS�.]���������N�9�������ԭ3ݛ'���H0.���u��vfx���܍ce���M/��0,��	%a�\�)O�BBCg+�����,��@�4d�B�uCg��q�m7��hܕT������V�&���E�E�S�L��d���:{;�6^�T�=����"��n�v\r%qz��˱6S��	`���Yw,�Y��й_���8��[��-���Ô}�QIDũ����Y��2��*l�����[��K�Mb����D|D������)Ĕ�0f�A�l�I;��B���Y������r;��8��>ə4v�W�5��>���@�87*E�n�!�	ee���V�V'��K<��UEu��EsY��n5a���Eˉz�jt������3O���y��;�*��t� ��i"�s�qwP��{�Pǋ=��7��Z�d�ZM�qYͫ�y�0
�D�NB��'#f�� �t�	)��<b�d���wMgU�Yv���|��&(���n#4�vlzINV�����!0
��P�q�T���r�E	�qT��Go� ��Ŋ*��NF���k/�<g�]��Ǆ���2��� ��ԵI����Q�Nzx$���D�ee~P��4�Kx�,��NS�N�(�'� ��:?ѻ�ݛc���/���^�C��;����!��Ep3�TVd����Ӌ�J��l�N�m5������js�^�{Hz
�#�����șdU1�Dry��%-��h�����$c7���z����%��6����j�3F��e����H��۶������'��<�%x���{"��.�]�6%Q�S5�3t�e{z����Zqi_�ɇc�^���D���)��ӑH�{y�[�]��7�^�L����o