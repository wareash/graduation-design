��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�uwC�5�b ��ϴ�	+�
Ct� "�J~���z����<
�����'k�z��ߵ,d�.��Z�Ӝ��2�x$ҟdL��h��ʔf��#
����;�;m�ȋ��[F��E� &'{=u�3jg�b�)��LA�u/5{<	����H$�� |=89ٿ��8r�}+�&I���.{�n��k�^����URIF�ڻ<u0w���9��i���fc���>>�*�W�u��AI�&��eASn�ok��>u�ɖ���ϛ��=[3C�ia��KTn�V\~��GU�9Q�)�:ʸW=j[����"��+��CK���G"`��XU����as�U�W��X���)��Ep�.�!���e�p�h4�2���o9����<_�\T�D�J?�Z�8�w�+-t�E�1�Y�b��:����7+�!�Cb⤧�~l�1��7�;�����q��Uk��WgㅜY���|���:1��)P���MN<:x2i�A��C_�m�
�-ʰ��*����Y�T�v�_�ao��wp@�ٛy$l�S�A Y��1��K��x T�2ႃ"%��m�~�f�������nd��iR#���V�~�fP6#��
m���j63R����S�/����e���_��1(�3���R��<	|�� 
F�Ah:L��� q[w��'�{Û�q��R�V��!���D��+3�*���Q�5L�Q�j���sꆳ��_#f}Ej ���,K�:-?	H'�z��/T� �,R�{Q<�??;�M��\�����x���R��p�ys�:C8���%tJ�G!rTϱh�1>wϰR����a�:�n��(T�Á���I�]����jS���'�-��r/_vz���	Ʃ�k˔}9��@6�ES!��(���}�"c���Ѓ��׼ܐ����$i�{ �l�T�����~�<:.�����/V�~�~U!ц�H�G�-��?_�!J>$5��~�?	sɺ��s1\U��2w��yGs�Q`lE��ԡ��G�͋�����I���Wg{�6�����Xj'+a��	�w]��P׭��a��mX{�6�%0�b��Y����U	����i'^�Ōq�V�~Á�W����xӂ�+͠]����,�&|�`��3�6�/�'`jp ��Ŗ�H������p���=eMt}M��&�	���<�&:S��S�:�e��+-��h}@	���u%H��&�q�E�|��"�8�'4�n�/z
�����Aw�i�U,ӡ����/��"L3�Kf��)�%���F�}���>�#�^A�d�a�ā�t�%��%aLƴ���!�	Q�����
V�RC����S;;�#��Oqlx�Yor�M�$���=h2�]7,��|E��',�G�2i5�������ج�	j���]��ϸ��d`E�c�Ѭ��4$�J��l���U���ȧ2�iM�fw�v��������:��/��B�<+�R��Z�3'w�U�R�'c��0��t1�گǀCkϒ�4Q�Y�����c���\�ډ��۪1�@�5[7�碜��RZ7&�����$J�F�66 ޽��O���g�����9AN����l��Ʀ�{]����h�K��b��!l!�(TՅKJ����)�	��q���L��(���xó���L�S7'���p��*p=Ifi~�����4+s4x	q�]�д���}��[T&D��iA��`���!���U,]s�6r��UP�Wg��E�ȱ.\ܢ�����$=�4�PJ�M>s�m���`"䤄����)��s��0�R� UxI=�qsĆ�t��߳u���R�v�dqV�Cr/b�H$�1L��5�W"�XMø���C����x7L���!�m��-�e�9!P-��8^���(M����CL�h�(���=�Z���/��B��S#��&>�%L���������ϡ��̵��DmW����׮�2��>��/M*�S��~�a��g��qR� c8�� �]��Z�>'�~YI���AE��J�lή�KSP�˩YN���o|�Ab�JDp}��C� �G�i�"�B�[�����Ӟ�~����
��8�ig[,�T�i�i���:��aP���@��~Z&tqx��d�d8�	��������`|�i�|&P��0Zz�H���L�x3g����6�D(�F{�@tNY�&JI�_n�ݏz�l.������CLܣ���>Ja��>	;�!������O"2)����agY�$]���4�DM�b�K|BB�b���j��s���+����i5���0 ߃�����A2B��M�=P)�uF������p�r���-�1ql L&&?��iujQ�V.t�@颼�驴Ø (����I]��(�!�5��ak��a哳ƕƫ��k��ĝ׊��Ƭ=<�o��q@�qQ$7��ҧz���gX�eċ�4�(|�Gk�D:��Y����ŘYHs+.���K�$��#��F�����ٵg$Ǐ�?��7����5��ڿ>�Q�s"�c	��6��4��H�q�Sh�[�0p�nE��@S͐�R P���<L���5{��`�}Q���)��r���TK����gŐ鮲���0'�|��[���lK�If��R5,�q$�o�fh�,�²2����8Z����>���e� �4�#k�(�cx�g����W�ג�9OT�PU$ޱ�����/�\ nm��@���,�e�@)����!'�꼲�<轔����,� ��I8��N�h%~�ʹd��(ury�Hz���,r����3���pb' E��0��q.�%k�iUN}��\'�<����M/o}�����Zm��Z�j#I�I`6h�@%6�ٌ��}4s	���� G�7g��A�3��MT6ϰ��l��o�����?�����@�l�Y�X2�����8��^+񑎙u\�Hi#����cx�e$��q�� �!��ݳ���C��&Q��4������@qJ�'�F#>��7i�J�����l�<�^U�S�эR�b��(n�r��cXꣂZƫ�L�7��L� +}2���
N�|�8O�u�����$�M~�o��u��Q��QY �N[�ʺ��Cmء9�=��#g�J�賚���lC㽷�u�"ܢ(�,/�V�p<c���6��		UzGYxX|�ʹE��m{��u�]�Ԝ*�p��>s��(��>;�R
�O���X`���z`j�fD	����L'vb�$�l�'Q#Sб
��!F[�S���aS�TdNf�d(�8���A|�))��16�n;�����{K�%�fλ55,�S�U����Y�I'[M�,qu�ϮP��U�`�"ѯ\���(��<=�Z�����c]7(9���ʅ�L�K	c�|�fx >:2��W'�])nϻ��ƴa�ȥ0J�p=���{9���ZANPL�sA\l�?���`��$I�'����rZ>G��u�U�49�	�?/�O�6��\����؈�Z��*�;#���x1}$��������+�DXڂJ��5�� #�?fUczr���?�i��)�I?Dr'��-�Ƞ�$��ʺ�u�j5Ϝ���Q}��������V(f��ةK}r�S�]{�(�����FH�3wX%]�sS#����f�.�#a|^�ՐmW�T��!���H��í⯪Fk`#�i&Ϡ���у�d��0v_���=#=��#Q��������-0��1�TS˼����wC����kVჄ��=���k�� 
�uM��c�����UkWŎ�U�y�S�}��<�1�|��:聳�ֽ^ُ�+4���%��a�k ^S�?_2�Mh�Y�>�4Եή�VCk��9�N`�E6-��0t��܁Jʫ�>&�;�'�Q>l��L��G�'�{2O�NRz]�[�9�Jӓ�����L��͓��Q�4�qc&T���4�]�9c&m���_酔��.ֵ�t2�d�w�U�E*�Y����:ǣ�?������h�GV4j�dWz�?�PGb7[0�hsc"	��8�N�/���Et� /���䣲�m*h[�]�zBP��.�2�l�.>�e����Y��:�4J�6�M�R��{TF��[�;�d@�2�"�g��{�{��[�����`K3-�K���"�ڧC:�i�7���q�ǳ�"㽞w�V��U������(�D�!��L[���:<#~>�(����㘯D{�=���uZX�g�m�s}�������<}�r�� ]��r�K#��9Uˠ��Y��9��ݸ7ΟbhxU�:ْ��R���P����+�(9g�����┶�;ߗ�í���O���^W�?}�'g����rp�а��.ܞ��!]����:�^���I0#�����8���)���7�d��t� ��$wz�}�Wm��YO���^įӑP5��(|�ْGL�}=2����gkH��o�ѳh]JD�$�����h�K��g`�Li�N�RP�V]��;[�����W�n�L�O:���<��e��8���I�W<�!C��X�G�.B{�3���d���uU��jkg�Z-O�ˁ!�(�/@E�Y�|u��\<���F��NK�~�h,�l����v͔���	��8ݡDҌUir5s$��$�R[G���:���ډ�ʾ�-iL)���&�2t�X)c�ړ��OHg�G&	E�=�leu�M�� ���ѱQq����;n`+�Bʉ���(��/�z������D��.�>Uy�/�,��`nP�e�v�=��K3Z��+�z�Ԇ����-SV�@hf���	0^��_�UGe�*�B�=e�#��Lw�]�����bs\�k>�u�Ϡ�W�=B7�qZO�� �/����(Z�F�MT.�Vc���vIZYpn��i��T�j^�}U��}r9WS��}��̧������r�b�L�-���ү�+x���峓��X�X<(�y���:�[wrV)蜎����M�IG���<�~�|��i���b� �m�C���u^**qD�*50-K�1�PK�yw���4S�vq3����/�}�f�˸DpU3�5����!��5Lw���P���� �}�U�IPd�+S>)¡h�����߾�|��B�wk��-��i�V��G3����%��Cbhr���%�0�rh>W*҈�H~���N������Ϟ�9)�*}]ؓzLkl����m)�'}�3�.6�7����+����{��1���P�Jg��~�f-M�m����1o����y���~d�y��I3p\V�!��H����8Ƥ� ıh�N���$,�ZC��<&-�T������P�a��K��p��,k�TyXEQ,��P�t�Q䁹cJ��D.}ډ�H�,b��������F���cAݡ�(����[p�wk�0h;��s�0��45�_ �b��NhL+���P��-:�B�jE���z�ո!M�C�\Y9 �!����a)I4eD� �kk5=�N�B8�KN��.�q=�\����6b��]�B�"��K�T_Q����{ȥ���<B��8�*��e��O�=��։i"U�u0V��*rJ_�7��ic~�;���.T><�C$�U������_�Z��a8���p����6V�ϡyyN��ډӻ�5;�j�����1l�Sz�f���ɮJ�8���y�}�wZ�b$�P,�ӛjt�e��*oZ���B԰��{k)_R��~	���T��x�-&����ʨ9i/���D>�yr�����nh����N� �@�/��]�ϩs_d����caG��s�bb��RP;�FV%g���I��|��l{�ˋ�K�l����C}_۲8K��s����8i�lA�kW��/*ڋ �rS����	-C"��ӗv�1=�涍��BRٴ���iK�z6�J�Lg����	���tg5��~$�����0q4�bF���"D*�F�I�;����Z���~F��ϛ���C�	��4�����T����#�8���)�Mq�����d[ v��>M����d����r�l��@�2�EB���͜���JDlDhhkBƱb�ܶﴅ�XC�*��\0n)�q70���L��՜Í�.�� (z���^6��\ٍ�vF�2A�����hJ�=˝��xݏ<���PE��"��?����ﮘ�J�Y�A��fl�q
�^y��Ş��?����/�Β�pɿ��$����>Q��\k���7Z5�a�\d�:��?�+�!g�E�!��q�$EjtkL�pRR��
=喃�	������<�R׷Cl�n�����Hh��1t�oxJ��^	�i�oK�����g�.������f�ւt��6�6��I¼̹�e���EuO݈���J��<�7(����~W�\�,�ĳ�/.=�ߌo)��+>��a\vI�Jv�P?t�pn�یf�]��;��]+��g]�$�q�I�KHTZp���,\�"9ka�]�C��Lz�*�b�)�e�>��?�����6��H�N��7�!H��/e�<�k�Q�G�M�_%'���oV1��HT���5��=ƫ;�����&F[�����u���ň2-�߷ᗩ�%A��F.7���iJ�y�KYb��ٓ��l��tR�77�t9�f*�C�}�čT��=�6�a?��^]��c_,H��܋�ER��c}囍�ѭ�/`��'Gq�2P�h=��0R~�J5����j"�U�)XkWӏ�s �4�ŀ�V(���X��%�2��ޟa�����	*ϷM�d�gl��'X�P����>j���[1��W=�65�䜋0F�"��a�S��d=���<�í��#F��/��.Ogd���͔�������!�����9ٕ k���o	#�����_�����ۇ`�X�Wu.k��K6kl4��4Up������kN��?x��)�6�2��A����5WNb�:e�P�\�m�Һ����MQ�:�����1�┱n�x��<�t;k\[N�N��|��Bѐ�b�Uâ�#M���[���ǰ!ڪ��4�����]��S)�@MW�G���P�3.gā��9��Q���S#+��ËC�}��L�(ӛ�	�:,��+�+�-��o�k�l�`b�
��{��2����)�����S��
e�}���.���Ls�P�eA���?<����=��z�Qa7:9�[v31��"Q_(Ji�	���D��Ȩ��B��,�v$|�d�p�ʧ�X�6^�v##�xR�l�J��� V�w�7��ޅ����?��o�g{��Zzj���G#�#���q!�d>�����$��"�ʻ�^��eK/G�av�a�q���;(?�r-0���s��4%��͆F�F�����۞_+���	�W��_NB����%Y�oql'� ���u���ĳA8T�� �$�슽Jo�߫����9nɰ�?QƢ�,Qx8�I�rÙ�,a�T���Ƞ���nt�r�lx_�%��D����lT/r"V���#{P���l^���T�����(=w=T/
�Cl7r&�޿Î@&`@��)�5�@	�G������p��uE��]:����s-���1�������	�{�z-P7�H/9{䃞�gje���,}�2ϤB���н��O�z��d�4���cc"#��,�Y�Ts�f�yN������
����}{{��3�\�4P�\4���B/p�:����u��;�v�+�L�BS��*jH�ny���w�� ��3Z�oK�dX�P~Ɛq��0�h�p`�Z���G5����J,г5S2V��>��ް?U�N��:�>�D
k���K��io1Ͼ�jE��젔�B�
�Q>�?�ڷ�{o�*��w�:#J�����B�r `�)�dK�2O$� ,B(�X�����N�Ll H�u�O^Np�6/Й�Pp�(O��c*�Ǘ��f�)3XpD
e��?��iƗcJ�8$��r(놠)��oX*�]�5�/�5� G��I�E�#y��j7V �F�C2,в�̇X�d��~D�ۈ�c�Q���Uc���{V�v�_���hNuO�C���Q��d�Cah�����ͻ�N����ֺ�6��*��%�s\��WH4ߣq�4�qz�gj&0����+p��=7p����:[�L ��$��5�-��Z�Q�W6���A�m�ĀiY�(��.����� 	��L����x�F����@�?+s;P�3�Ŧ�e��9��Q�S��%�k!&��������)PTܨ�r���i#9ǉ� ��˻X0����C=^d�U�UG�;�mx�B���6$H03_�2�n��}/�cVa-����<�o����7�5�"%7tXX[�5Sң�0B�t���ǒ-�eSկ��;�g�p�}>Q��^�QX�g�>ߏ��<,�\�&x����a|���ख�?�&��"��ko��+Ih&�Z���<�x0��_��J��`#��Dy���k �h@�&��xK�;�$mv��dݶ =Һ4x]�K�����ϩɶ	�����<�h����+�Ԅd��Q��Fx�(������ȕ*��x���#�v���E�,���}�(��3��qR�#�~����fEem�j�G�;r�!�"'�~G�k������W"���n����y�����d�*�����A `ůAE��2���u���#m��5�ܛ�+�Y�3��y���x�-S�!��	��)�"k��8�S�Lm�4����{.�b�1	;��G=eh���z�;�)�9��N��QNG��U�g8F�i^젖��q���������w�e�(��E�s �6��>X��qa��z�.�K�������������K�QL;P�����(ՌQ��3k�{D@_��ݞ����t�P�w������ʭGטU�*P@�!xvZA�Q<��ދ�ۤ�m���+L}Q��$}�������Y��B�D����G�s�AMxY���YSc�M����{��i��ҫ���[�Λ��|���N۷=�k�Ǒ~��")��1�dZ�]�뜁�Z��*�~��:5�1d�m���!��7����@a�W��e�b�5\�"��,��-�d�!J�}o�%�����%�Uû{7f��c�рzqw-�k)'������P:$���{K�{M���X��'�J�4�|�VV�f6�8�+��/��I�#&!W�֝aߏ.%m���=��E1�0��Y��zI,���]��g�P�b�
�O|�TU��y�NQJT1�J���d���R�5i��ʛ8%K�<�U�
Q��X|�f�YT�r�[�?��(Ү����0�9��m���\t<7�jg����l�{r{1��fm"^���L(�K��ch>	�ZH@!�;@̛rؗ��߂2�u�?'YPY�(Q�/Y�c�h"�0%�������Y��[��\}�ķ����#+�7�˭ש<�_T4��V�%K�}�Ɣ����^?-G���|�h�
�P�<��d�/��L"���hRA�p�?�Q2M�f���ܙՑ�y�%��k��&;���o*ݽ��7�0��"�UY�x�\�%	l��ߎ��.g���:��&~ו�Y2����M�?�
�Aj78��P�W3�+�M".���諾�<nf<t�
�Fd��aW��P���~��hxX��	P�ُ�  �����M�=�����]u��A��i�A�����g������|9�fZ [�H�O��;��������r���������Q�͜}���tW4n�j/�B�� �^�#h(���Y{�����7Ci���\1��(T�~"'�}_#t��QT͘�t1��T}��_�u)w�~�����"X��IO�ȤBηy{ڙK"w��^O$�����R��X��o�X��RO,����>s|q�I����e�JK���Q��Y�X�Q��*� j��K`_B�#Z�3��Ӝ�3J�;m����R����gI�����-OoFF+Yһ=�[UP����bq�
Y�_�dS��0h�ߛ�d2��"�]H�-R���D��N��<V�S�'Q���>";=�n d2�I��@n�G��^$A��[d3��#�>���iF�E�gd�z���$D�-�R���R1�mF}�Ao�����m�>�`��f�Ÿ2�Q�c�Iد�GJ��E[�YT�����rd�yWޔ����J��8�}����$X��(�Z�<�g�Q�n�I������� b��6c%Z��1�O�s�Ԓ��[e+B�\��*Ic<�����R�7�<�2�)��Q�m�o�2<$�����Ze!-B~M�@6�OJ�F���I<��bʸ>��w{�Wg��uP�����'hݧK~8�BW���[�܉�tO8���ț��RD]��z��}�~Q4�	vy�90�JwD�'�-:U���E�����$��v�_S߃�L��rC%�a��} �N� �l��ì���J�C��ꚯ��U�:Y�a����>�˹�U(�4��e1J7,ŊX�:{w� 6d��$����_�PԆU[�,�Qq:}wC|�HIZc�}��5/��\�d�v\���A��i2�������>�+�3�2�BͬHk��[�5���s�IU�c`_�لP�Nk��Jy\��H�����K��"eC�F�E9����f��5R���*t�M6ɡ�7�8PYU��v���c��^X�=����ݤ>�/��X�#jQ������9{m�O����&����{Bk�xS��6��Hig.D΂-��|���	/���ӡ:����B��T���J;�թ�KpVd<ڑ���H�a
;!P$S�C�l�6B-�6��{h�ƏL[��5���t �(���0X`v�-�	�s&t�/hƥb�i�N�2�� E���:ɒ�#�Xm���]d�e��%ܴ��2� y��q:��R�w�z����"�}�6P����xl�=Zw#c���`�������".�R�[���5�9P9X��Np��?v@�et�U#�M�4ٸ��R���0�� ����w��D^5��]��1e;|ƃB�?`⿂�A�C�N�!�{�2�ⵞ�c���_A���OK=$�&^�����;��̹��d�[��A��4���C�$�e`�кP�<?��ۍ� -��*g߼�9�#�'�C���W���U�"��E�O
7f��Jm>���6�z#c]�ͻ��)�ń������`1��C��W¯��Ӝj:8+����!���e	*��a����bY�\�am؟�O:^�&��VW�O��>>"(���CE�0�����K�֪�[n[a٦��P���g��Qҥ�V��^_֗."����:d%�������}d����b�!�^;b�U��h��Mg��x��fs��a�	y��wpDZ,v�@i���>��~�V�Pk�=$�sݦ�
G�I�떄�ê��� �w�K�.*Łg�|��7��'Y��3ٖp�_���j��{K
~�n��]�I�F����=p���Z��8���Z�sv1F�̮�5 tDX�ROB�dى�1���.6��^�	%:���o���!bs�M��~/>3�ec�͕+�zcr�zb�V|n���=�%���f{���)%�c��2|]k��x��L��g��O�V�^���������7-:�"���k[՛���,�=py�!A��(1\��,N�W�]�} ���[��p��>,r[k��J��*�Q($�F�>u�MN@��Ia��ě� �<���[�7�M"]����@z���o��(�Del�ԭ@D$s�����`�=�r�hc�Y���R�Ty����lJsӷD�_��O��_Ԙ!H�.L���<v{�,̋�o�+��ʜ������,[R�|Um��װ��߂�EN:z|�(��8%�g ���͉�[2�)�p��$���"�-�d�EOxWj�Y�s��j�!��_�F%B2P���Ϝ~l%��>��rRP�	�(��%.�dd��-�����{�f'W	� 3��Eb̫M���$JqD���^S����FРؼ� k�5uM[�R%���8bt�p���,{j��p@b�E �8[�ʠ�B��
���tN��s�h��,O��d-j��-����RK�$x������Pؕ *�o��)ߊm�A(���^�{$�F��{�m$i�ܰ�vBn�Å�����c�����`����0�T�cu.e��tx����q��ܿpK���hǸ��7��w�` NJ�	ma�&�Z�M�ܛꩻb�m�������v�=a$Jc#m%g��G⑦	����Ė�K��+3��q �0WMȅ!Ы���x���$�w���O~�g��ﴃ d>T2^>7v������OO�Bz�[���qm1������llm�z�P��I}ނ!��'��凍J�cX���,W+g-�8�ֳ�U����k���M@6�#!Ld��� �k���E��E@���Ȍi�{��ea�����^�����:�惝-Ek���c�����mz�^��a�M/\)���\Z&���V^�DI�z��'���͖��w/��t��fV]�묳� 9	���m�3�֖�C�����X<���2t�������%8x�h���W���4�K0���(V���<"�:��0�_A^��G�`���j��<����ln$�7���2�b$�r%U�h}�A/7�j��/�pX��Q���7�����\�,GO��� $�Fw�Gܫ�@ȃ�ۮ��4�2�
���k�	-�%�g7��%�D)�ۦc���¶$r;�J٭��w�(G���'-/y0g峱�e���C�e.x0
����9r��%�joV�Ӕ�#�!3�CG�J����n�
V1�z�$����0�D$S�UK�R���ժY62���j��u���Q�7��o���Ad�������[C	���>�r��0$�7	d��Z1�� s%������1�2��Xz�:�S1N1L_�}�\�{>|�9<ZLU9��#�O�z��lE�����Z������
	�:VCl�����;������k�E��	֍`��8ph�#t;�k���X�?�|����##>A�*���<KR�x���^K����Q��U���o���e�8t��M9l_���f���'/(]��(b
s�曏���C��.��Yn���n���K�>_�|/i;�{­i�\#����I����b[{=K_���Oóh�B_����ᾀ
��v��37H�����!'kK�l͛k��X��UU����i�Q�A��� =M��s����pՙ]�~-7}sDj������O�U��D�K>�:p4R��� �29C�QtG�ӌ%��
Qn��ly�넄^����<=��N��誃�V$�:ע��ޖ+�CM,`��#�k>��X��a6J�ڻa�;�a ��~C���*�S	���ުK�(��hcGY�|�ަXV@(]n�ElyV��E�D�Sۣ�j�\�u��<���ڻ�f�V�,ъ��r�7u���.ᅕl�e	qSb.Mθ그_��2��O��K�(dh�w���X�*�SOɛ�$k6��șNB�?B��2��N��0�.H�s��Q�'�����M����#�]�����>X�EU�V��6CX�+5+E�L@}��9� �O�8����E����zj'1��${#�'>���&�m���(C��^%�Ʀ	��6z�T<�@�$������哶M0qƺ!՚ �uZĘ�+�^��/�މf4|��Ν
C�棂��b��u �E�2�S���c��+,�~r�B��`Xq�}�����I9R����%)� '�\v�Gcf���e�9�?���gp���jWû &��9`�C�u�G;�������|U�gե�G�������%�x2G�����y��X�����˹���;6})�[u��[�Ƨ�JW�Z�ܑΆ����Ew��XU+�DǴ�d�IX�">��:v�����0�o:��OZ���`���;0����49*�~���N01�V�{�W��ҔL,�&����_ݦ�h�T�A�K�0T��i~�AYl�`����E�uS|q��$&9nI+=cs��cD�meEI�����w����%�"5��n⠽�X�q��s�u��eEWzSY��5x�+�i�)��]���=��a:j〞2c�2]?�(����@Ƈ�wRK\\L��KKPm,�$q�/��k�r�N�5"]	&G&�d�>c�����n$��*�y�Z�w�Ej�\n������-��_��S�d��:8��y���ʪ������G@�T&I�\np��60�_,ы��Ձ��1t�t�h�"��{*����������Ѻ
�D��B�)����Q�!��R�2��ގ���V����5��n$!R�쭒����:�4D@�.I�lf�����"��_!"�2�d��Z˞!qvH/\�ִ���5T��?x���xv��n����k~`>�����6�B����I�2��mi��^G>�)D�Q.Bk@�3nS�|����Vl𤒊�g�N��3T�H�ྞ�ܾ�ۀ�Ӣ�U��N���AP�Z�4�r|&�x:�a�U��&X �S��xt�8+�\G���G�j�ɑ�A�[.V��'� V[�`��J�� (���;h���I�b�_�ݫH�M����r@:�؅b�9����Jک\tV�ρA��߆ɼ	��s��zg��^a���ܺ�F��ՠ9��ӍG���M��{��!˨���x�c`lM( �m 8I(�Ͷ�M����;-��XБ�{�磌`XU$���_��6
n�eѳ<})zM[
JK�~�B��I����I�M�.O�4�戓t���(����z3��2��Ӧ-�����M�����ǥ�h3���@�i��"Ua�d���*I�m8�5�x����M����(L�H1;^�s��t�?<���!�v�� �6�y����.���sp��6!YJD`��9鴋M�|!?����E����Fr����2��{G�=��{�G4�B����y���T���u���K�}���ɠ�)lέ�Ά�e������0�������s��G5Mg�,��5�L�x�w��J���X*�ي(G��HxѪ^����ǫמ?��?K�xt���M���]�/C��o�$�8RB�_� ��"�(vDm�`�w�.�A]�0B�뉤��P�Hp� �X|բ7@'q2�c�F���n�ay�e�u7}(���v�f�X ]O�4�Mwڞ�P G���op�m�{$��Ưw��΅�I@��,A~��|���q�BRF���U�x�k�Z��n��j��}F����w�|T��r�%���6m�"�ߤ��R�U�΁��c�'��r+�@j[ݥ_"�&������}@��F0ݴ�WC
�:kg6�U�v�p���b�:2Ȏ���,�L�o��``�N������r}��E�	c�j`��=q� &��>�~�B�>�����ܬ���6[�e��l�[?	�u�:���R8�<FXQ�,�NOg�>�nK�T�'�^�4>�K7WR���
��W��_V����;�`����=�(��Dn
N߼�@S�����q��o���FO�I��mjčG���aЦHQ���ù,ۓ�����A�QU��cI{e��Wnp��Ẃ�k;p��Pk۶�\��O�#T}��JXLl7`�*`΋e�5i;i��֝�{q�f�bJ~��L xJ��	r�U�o(ۆO)�nP��ԡb�j�UK�M�}�1�X��]:���*x.rҎ�I"��#���/��-J�:����0Lz�
�,������\�][}�E��C�����o����j=�G���){��o����_*�t:���s�J��s��m$��Xt,j�ߎ>�Ch��!��FX��¤f�%&@K(��nEӊ����ڃXN�nlv�g�jy��*Y=I��5�k76��Al��r:��jIIh� V�A��xR^@����e�u��8ݿ!��>&��]�z_�2I�b}�z&p�nZҐ���/ �p�ZsM��S���]�v#����؋��Q�Fg�2vƜ	$e<n���G�l2��r�~�u>4�S��.�����=��z>�`y�D��PK���&c��)D�#�M��ݼI&
����E�J��ھ�����ڹ.��D)A��9�Û���d�h�22m�C|s����!Sȳ*�V��F�(ql(W�$��<v����n�حg^N#~C�|_���e��I^��ڬfr7H�X� �}�� ;ɓ!����2`�w6?UC��&�\P�G�U}6X�R�F��4�\����{O� �s��$�6�D8�F/˗~I�Ԭ��"�bT6K#�h  �%�౛�>c�i�v3��*��X%T�Fb���GߦMJ�a�����:�x�N��ӭ�eU�N�P^!y�TV
q��b��f��>Ed8��O�B�d/MvZ1m��A{6� |fk�[Afc���ܚ{B>	R��p��!�I�s��\���&a�w�:,0�c��I��`���!}�Rȭ�ҝ�V�z.��v�,�u<��΋��[�^\�ʶ��ID�+���ɝp
��Z�9��]{u�ܩ�I�K��U���q�ד!��  �^��((cߙF�Cr��zZ6��0F��)sq��~aթl�)��N���"���jT�����P�|�Â<k �e]r�y�����A���y�<m9��&�ҽ�Ћ����&)*Jw�˼c��{C[:L !��ݧ������B��~��$':�v��'���������(}�<=�zg�/qo\-�=C�]��s�&s�z� 
�����\薧4�I�!��B��%W�t�{���Dʹ#�]B���p�%��(��Ti�!�t�yb(�>छ�s���3��^���H���n�E���|q)�u;yq}
��:�����)t� ]�ң� ��<�˿���EL��4�CfM��x�V>����1���ٍi8��gN�]#/�|��*���T|��K�l��]�{o�|\6NL&����<|/�h�H��u���u����2}���Ar>՚�/]�7�Z�~��@^�%o�����ݜQQ���}X��^w̗	�ZB6���b���}:?���k���,���0VT�mā�q�E5�&���P�[	ZG$��s�FΔ��	  0�3z;dH,͌lgi/�d��~�[��~�yk�DŇ���\�V��U�N9�*�;��M��(}a�m��4t0�"���7��2�y��(��[ �7�����u���sjΏ@	qN�1�f!ͽZ�B�݄����vn2�^�l5��i��+&�J]fa��)��G��W�Mh\�)L���UX�&1U�"q��=��N�S:3�����W#�L��|�"q��ś]D�cV9�(j],qb76�?��2�[�(�k�����ys�	&%���T�M��������<����c����z��.)0b�g�N��y��b�T�隞�<�j�W�Y�������bJjI�q��ʑ��Ń���X����
���,�Ld	�w�:;$�K*�ӆ�@O�9zu��K)�B�����[���"��u�wE�{}��a5�j�细�:�3|�xU�a�)�>O����Cݦ�Fi��9E�ތ��Z>��V�ы��r�����Q�y([��,$��6���ذ�\?z����!�ɏ�ޘ���b��1wuǭ�a`����c>�z�����+�a��7p�m`����`:��EO����r8O����z���3�g�W��c@�=N��C»��<?V��H���-�9O-�*���|��r��F5��	_��x���f��$x�}��S<�no"����۠��>�A��������)o�<,�q�K�9(1�msc��c'&e��u�b|]�@�K�i�eku,�x��<�Ӥ��v3��@V��5}f� �TM�\Q�����)dIto�/�V��( t�����ϣ�,X�n�1�e%X���͸����QpY�(�Ձw}ɰ�n�{��&A�G8i�V8+I���ْ��j�(?
S��5{ e��Y�W5�@ОH���Njq5D��7�ݍސ�� ��y1A*l��̫��=�A���E��7�w!�t9�k�Cd`�����x��H�gF�{����u�nm�J���Q���z�c��6AoB��)�E�/�:�\��3M]�7q�8`�_�C��j�ヹ\e�,��!��9�Y*ok+�.�C�c7@���01.�V�=[������DJT�5�����[
�HrZ>��\w[=qF�n~-9�1m�^�F��)Q,%Ʈ�r��YjsR_K�I_�y����=;,��Q��E��-i��X6����N�[�62�V�W��Oi�N#N��,]��.���Rڂ�G�;Ct�9����~�Vz>�����[}x�����5��%%~��4�ϖ��
a�9�&��K�[m٨F�njl�`���V��N��%��D��ݠ�]ME+J����lbA�d� �_8)=�}��dz����5�O=�Q�LId�*�K����L���4A����@A�"I�����j���ƕ�k���5lPQ�ӯ����NoP�����0^�xu�*QX���D�[8�Xp���疈�]fe�v�pcy��n����a�E[�Xb|h,dC����KT���}lu�����ʜ2>��S?ᣈ��1�^��X�(~�bmv�'�``$.�R������ҩs������[�~7��ѧ�Ne��]��>d��䂩�s:�E�8�΁��?6
7��:Ca����Ѱv��bW�˝�ס|���O�����LFK!gb���dE�e�A�8ӊ�s�\A��q� �N�Qp�������g /{�)����]|�¨�[�q��HM7f�<GtѺj��"�E�"��tE_��tL��+�?.(AK�Ɩ�{�ي'3��
5wעE����@��.���&��KWyl��i�f�ɟ��p�4�I/��18cKt&�#ɥ|�t[ ��j�7T ;㯐Y�"8���8.�X��U"��S�ܐ��F� ����I@�}�����{�BlB��<����F*9��̼f<��I^�A��&������p��4'�%�Y�17vʣ��p�ϋ)�߉{*�X�1l���r�*#�A~�Uc͈�+h��h�vW;��������Y[� ��jA���ʪ+�[�q(��NdH����-�b*<�@�0k����PŦ��L�M�CR+���6�Bj!��kB���-g8F�����s��	Ai�%�4+��Y�%�I3^����B�ޭ�I1��z�q(PO^,0)h���\=�xƃ&�DW���)L[��f��Z5������+���̹F�q����L"�0�@�/�PD��1���Q]�`ӷc��g&#KL�4�[0��Y�.�IM5�vkZ�f7��R<Q�%�9}��A��Dy��Ǜ�
�s�wѓhVU���<�8ۇ���-�7P�W��"�4 ���h:��ҟ?��Pa(a��!�p�<��'~z��|�b�&�>�WDL�S���sd�t4�(�������R��V����+�y�\gR�:�8�6�D�!�\��7�Q�(l���h��䋣v���輻®{�hH�D������-����$н��Ro��6S������\B�l_��{�H���Q�W�8�=fl[�LNc5h_F�S �i!��|�$�Ԋ�*W�s������9O?kJ�n���Iq��c	5�����?���kn�R,L��<�n���^��&԰y���(��v����A�.��^���?'��]�r's�b�!49��i��-��/�≻��c_0@|:/Jy]��-���wA�xrȄ���Z%n�� ��+�J�P�Z&������GY����x��6������b~�j1������D�;�P�p"�y��]z!�	��>ٙ�z$w�����j�q��i.'so�1��, �2c��{	��9�*�I�a�;j��A��7u'���70��?F������R��YE&�c���јo��A������m�]�h�e>�.����5䚔���t��*��3���j�fD��WA�d��C'�q�ǗfV��Ch,L��c�j���~N^�tM#/��o��s��Z�KG���!i��jg^pe��8���~�V�|r�߂H9'z���͓9����WmzK[v̎3^�Q����E%��/���P3�^ͬ���8,[�N�@��k>�����&�jKK���-`Am��m-~��J�!�+�Z%������?���8)=�#8�x�1��8d���c�mI�Y��9���Mǧ��'��4� ��FBeV4R����.+ƾ�r��y��v�y]�]bQ��bb��@���ui�*?ޒT'����F0���D_�lޥظ%0�ߢ�<4u�����ԥP�Koؿ����X6�!�P�J����Y���o�v�b�O�	����J(xW�Æu|Ä#A�����[�Wz��m]�9��eCT��|����8DS��E;E��q5�֟�9��2�"$�WQk���8@l�R�͏��&�I�l����þ��-��C�*��@�6�ĳ��Ζd2�r�S�WZ��,��}kN �����\�]%a���ƀb�m�Y8O�� jZ�w(��Ӻ}�M���\��X$�ù�$��J�t�K݂�
SW����ӐbZ�<��q���hW ���̀�]9Y�Ĭ��Fj>��2����!���A�@E9��}۸/L�(v���h�v�޶��U�6�l%vY��U�2+�r�qM��L��xi��a.EM�z�=��@�C���j���[��ҷ@�2h0�@�5_>��j���B�<N8��9>�$-p!�u4�#�_κ�ϸ�K8#�B�8s�!e��U�&Й����u����@�芗�k苈@�f����Y/��T���;.	����Md���QE"oIɤ��>�Y��.����ә�</´�B����q��ȂƋ}fd��Cd��x������-Q�Vx�o��z5M~�����obg�6�/d���<�^��/lu�`�a�<�F��������0=�:�*+��6k������Z@�8zg:T��yX"����2�dM���tج��axPJ�=�[2������*���=�����=*>��
�ɤ��۠v��6�U)���.�Č�R�.�5�_����i�8��H.m"�V�똱�U�cJd���
�4R���W7�4�M˃���(�!�	!&�&k-C'���C�si���E(�O��������S=lh�C	�@�ѝ� 3��J<J�,a��}���,Μ���@���e��crGZ����m��Z�P7.�������B��r���s䠶UQ�ˤ}`�g�����)��y0�\���/~�`���(a��B1%i�M1v3��dm'#��2iFq�����%;���1{чY��mo��X��Q�L*7}]�`͐�ccKg���<�oc{@����#��O��2h4-B�0�;+���2U���TP�r��9%�7Um��in+bY���N�(��93��=��ўBP�4����R�����&n&��x1�W0s��/Mf-�
?����d動���uF�K���x��ӣ��d�!��7��x��	 ��h~vﶹ��v@�`���o��-��@��Ƣ��9p١���i�7�����p$��g��CJE�����L�:_�բ�T���i�ٻ�Kn�p�l� K1���O/OGM���d�o�$�W~Q���Wtٷc�^605�D���
�x EKy����)�e\�+�c;%�(��� ���N�.3;��O�p�_�x:Bv��{��e\!׸uaD;L�ުP������'���&@��`��X��}]��l��}��ep�W��Yң�diJ�x�H�`"�í�D��;Uv>��6���e@�TCl~6 �sG(D�M����d�[��O0����5��>$nlUf^��䀀d����Jg����^�OJ�q�R�!�N��Qes6�Z��|e�E��D��T�y����?}�����Uq�yy�m�4�e���JD2��(������`e�E	�)���V���������nyF�.DmpQg~��L��\��^�*�9}�i5M�AVBnW͠�~�������y�Qmѕ�%���V�����VD?@�Ϛ�K�]�k�۟g|��͐ɤ6m�ڻ'w�n�0�b����O�L��"�2��5yD�첒,��� 1��$���:9{L��=]`!s�?��%�!\��1��@�bJ��d��I��u|�4���z���\E=%[��L��Gʘ!�8,#sX��:/,�b ���֋�'���!dj���e����ȓ�/���8'���a��ʌ������LJo�h����#1�kⴟ��y!_�a18R��?!�� q����K�s������9�/ٮjC�#GK�� �M}��Ql�S��%�'B��~�筰��^{�^�����E���w��$�7}7R��=ø�V�F_+,��h���v(�/�*9���9z�&�]�T�m�9��IU��9YD>)^��X����O&v����w;��/�S˛�>��%���O)�[�F����r{SĔb.��b]=`,M��ѡEB�ԙ?��&�osnzI��rބ�B_GP)�I�#�a�K��,wh�TɈ��:G����O��y��,{��BXl( ��Q���NYrHk�1�&I5ߡ�������4�3�'�L���(A����^N�����X��k�P��5�ZL}��T��x���O�EM7I��R[ ���n��'H��4A��*���̽��q�ZC�����_�T(4�,��<I��=�WM(��V���I��a�=���g�{����|��#���H�B�����Ų'N�RK�? Ѓ�~�u;���B��0c�:�$"c�oGX��vX���&u�g6��0! ���9$���I.l�7��7]	0��-z�04�At��I⏅F٪�dJW���Un��,����qDG�,�Y�&�B^!!��v��d��*(�]�Y�1����z��-��tR����Q~�W��ZgF��S���	O�BV�J�:Yњ}s�s�J1�n2��HC��7
!*
?:}Oꈯ$�C�|�i�F�� \aQv�F���h���1e��p8B�E��J�?(P��"���4A�*��w�J	'����B��YSՒu6h��JYGT�����ƙUz��	?�v8�����oG�\���~X3����<����������m(U���z��;k�S3&fa=L��9k�g4;�i�@/=V(�$�}��KlP��x�Ѽs�A̷'WR�\=��XP�V��Ҏ�Y��
���B[��3��5�H�[ܻ�L���q$j9���0޵�<joO��z~ŧ2�9�_6����jL��	b:t�K����q����k�������3	���<G�x �W	f`̆XD4#�|e��HU���aTÜ���T�R��ЯTr$��'f�TX���3 ��>K��\�f��������\�����Ċ�'�)�$4�ۢ�+ʽ}��Pm��R��n�h��Tŧ��P�O�I���x�����y�q��؉���f�o��Rh��ʋ�1Nx��P�q~3z�ݐ�>� k�Ӫ��D���!?���K�>�!�V�m��/�z��v�7�Q�.L����z�oSz�!'���cul���2oO=�,�t���=�
u�ZX�OT� ��5�ݚi�~�bj��ޗ�Q<���_k�����N�1����X�ݪ��;���� ��JC�������?;�/�Hp7+��x,`o�^�Fv{$������q"���S���>`G�bQ�z�8Qmal��$l��o�ݻ5y)�K�l��ݷ�o��\�gV|�"�P~���_�A�]<��G���Ѥ�����Ű���s�[�<	����ac��)���
~�o5�Dz�C�(W�|��RXݭ&t�9k�nj�ؒ&0�DU��A�s����U^T�Zl����5Rx�9�s�|3*yk����M��@9��TPS�2�@ķ�����_v��m�q�J��x���%c�O�u��tZ�<�b����1C$�A��l��#l?�Ɣ���hA�*i6�oT�}4��:L�]�Ł�p�`ò�2yH��]�.N&�W+I�ֵQkj,1W@4'g�����#gG�2�<��LO�����p�0'>p��1�����`�ý���َ+���\�Ic�U�dP������n �4,���vNq&�Qj���,R�̘y�]�^lS}06=|?K=[�<�rF��J��ǎ��Uw��������b������K��D}Lc���*潜m��Q�Y�}BJ�_O8s�����)ij;fo���\�4�W��..�Y�VI�
\�nk�[����	���N�.��H�#�:���9ܻ�Ղ���6(���c셓�ņ?��4Ψ�9 �m�1�-��b`7bF]-V�cok.����*;y�_'�M�9fSg�M�QO�>u���!�����>0X�ڕ���<�ؼJ��Zf��f���\�떬e0���F����0@�$kyW&��i�4CM����o�W����/��'�A�o�8�Ě�F:.Mu�P���2��Л�f��Ym�1�ǚ+FF�*��'t'�_��6�U��3&oy��>��ѻ���%�Z^_\�����l/�"���mY���*�Q�d��g���P`��[��v����i�ҟ���
v�[�>�1gZ�~ԘM�����	�t <��f� ���ث�h��{��l��&������2�9���9J��lU2�.,��QY\�F9�ᴟ"'t�,,�o�߰�8̸�/R�G� ���!!%�����]� � ���`��Z�g�K}l/%J�N�j��޼TL�MAe9�'p��t2P����Y��(B��k�B�J�mnɴa��1������Btf��v�J���Ri���[�Z��&)���(����G��V�֟��6���18�#q�`&z\f�#j$�&��Sg��k�F���-��祖S|他�.���{�K���GUݤ͋����Z�RA�\�����!,_C�M����c~	Q/����}]�G�P���&��P��!����cB}�P����0���8�$k� �[ޖF�S�gK`Q�1O&��ܒc0:j�w
-$�߁N|��\�g��U�_����%��^3�a^�mPщx�-^:*���fZ6l�p«xLJ���"^��1'�'�+�x��#Ż��Fncޫióжfs�U_�*8}T���׶.i���n�?o��-��3��.�m(6���"::Mˈ����V4n ��s���[%��zCy,�d^M�-��&@�f1�&�D��7P{솆��Hߐ�z3���.�A�k�����*{�fîYD��y���I��u4K�l�T��<���o:v��o��]k�z7��������M�+~s4[M�D� �<|�Ul�*��:�z�/���v���.�Ʊ��ٮT�������v��C��ZP���͇K"�㙑׭P=�~�읜F!�C!��<l��T�EB!�Ɉ�GBc1�-<>��#:�k�Y��.Q%/�XI��_&����|�P�@X��S�����ږ�Y|�{���u"�����[FD�N"D�5�
�<T�:tR�+�I�B�h���a���>So݉�"�8e�����S��uD�v@��;*���Z�I�P�'��R���� ���tkB��v��
k �P�5�}|�*�zF�3�'�fi�K�̕���ݤ�q���P7�~kȰ�����b4�����*���b��@�Wlǜ�	6�`զ9�kޔL���Q%�у\T(�<!�\ԇM#�R?��t�N����>������Gt؜5�6- O�j^�:��V�'3�І��g�HG�����2��T���9����f����]NE7���,�껖�"�v��T�P y�R�E4C0>$�&q� H3�'�e���[�[�)����'�.��\�N!*T�����"�q	���m�L7U����w����l��8���:>����W��f�dNi���`< ����֪ۛ�&n����Z��Bx~0w��Æ�m��J֖�"O�6O���hг��S��X���et�]]�HIa���0j�WwŴm�^G�����^fQ�D`ej�JH$)l��J��p��g�.�6(��j�!ii�9Ó/S�l��1C�;t�ҭ�ISD��y�b�"��>�'%��ݡ��>9�w�ÉU��X#n6���q(���4"�!h^�^��
L���4�k��$-�	��mw���j����*���i�3I3Y���n;{j�*x8U�~&;
�պ�K�IqT����	C�Uh�6��.�n,?�'ݑ3'X����\7,��L�@艎/<`'i�AK�?^��p�
m�1M������ϻ�� ��̊��G�YY^��2�T���[��]&M˥=p��,CN����[=�`C���B�ױ|#���0�h�/���DHW�s*��'{��q�y?6�LZ�����Gu��<��A2J� 6��!��A0W$	2x-���/\+M��.�X�&�=tT�t�w��Ħ�֤�s���<	<�CE�s�Q�ʏ���,{K��$�E�W��W�[�&�2N��}�,w�j�X�7�2�U��`=	�^<l�����'|0��9��4�!ȷ
;�"���VXn�x&9��ס�n����G���xݭ�]�(��F�&���du�?��K˖l�9W���Kԥ��)�s��8-?F
��eL�|��&���#!��O�"�F�T�:����M�ޞ�z�\�])�`9���YO<���������]�'��?�L�:;����.qm���=���i��춰�ʃ�9���9���ە�u�����;��Li	�䖢5�O/���?��|�"KQ�N�d����#����5�
E4&�h����Gg0��6S�����Ȅތ�|]�S�=|'>ӳk��S�.廲��QV3{��ע��ZU#����ey�r��!� !���������,p�Ձ8�L5�[��y��4���[�|�P۔���-�*�#�	�/f��gT>�������^3|�H����P�{��9��/���U(O��m���=ф�.pc�}���r�s/[������ �e}x 25H��Pb�s��b}+�������-2q��q_�|�O/I�a`��ίW�����R�L��Ou� �>%����s�ֈj3���|�^S����mYv���W�z��Ǎ��g�ߊ����l�A�i6� ��O�|��<��I�VA4��'�����:�%A3ҿ�t��OC��%������'���[����P��\~�WV�Ws�MK˙F+�$�ķ���4�a�9���a�לǍ�Ew�ucdwƮ�<���W<��!����U��
d���kVX�g6�J-O���Z��׎j3�<��k��ư�(L¿�3,����B�m�1�@�g�:Ś�����PO5�����*�E5���C�B��4�I�2�WN01g�|1<���tAB�cEq!�Y��&gP�	b��-P"6J�d�rgBb1g\U�^��ܞ�U�\�h�K+UJ��??I;��Ezv��ID1'W�)θ��Mt��=,�yP9��*�,Hn���V\J���p����q�4�M�WY��7����>��ث���[ѳ�I����x_�P��3�(Q簀8��5ɓ�0(��[��g�ʈ�S��e7xe�ݩ��9|�YT���N�E�5��8����B�Hn��{���D��!Q">����.���E/<�B��6��Z��g�����F�{�����UI_�yE�5M�O,����f���D>��b����}+A�L������P�,�MM^�O��|D��\�f�M���@�#�`a�} ��
�q��1���Q]�������J]�Q$���ڝ���8���j��C4UY�	p��<�A���FR�{$>���1�l��eכ��XPRg���6����V�y��[�g+Q�s��k �̦9���
FK��N��d����2t��i[pa�ٶ�	R�%I�1Mʼ���ۺL$���5���7F[S:а+�R��X�|��y���{�7��;���j�̦�>�v^�x$��RMW��F>�3/L�%��e�愚����=L&v�k��9���ƎN4n��/O�Ʉ���zZ�=l��2oI�}0PD����<���W��g+�(w��=���̺�3e�h�ZY_�/i��=����(_*��`*����ꢿ8�+Z!���}0&��C}'X2�kRBQ|�8D��%\W���������x�"�f��a�J+���R�#>r|��˫�.�����z9a�N/	/��y�!���=k� e�o���5��8%u��[N�&	(?r)mH�J��4�%����/>������+ ���s ������&ь'��jn�߻�����$�#�j�iS�v/���!���z��a&���}�������Oz���i�2��(W�DG�� ��ܑ=�A������fR~�n�f�M�<�e�.݌��0�	Hr �������H���2� ;}�	��F�F�ԲU�hĊ�Z�IĽ�����Q׊k��$E/��S�C����>���*���'�,B�HzK�NT���"�83 �PY�Y�
4L�#,�cy/r�rĆ$�z�#v�؋�_���,h�V����9�T�t�qu��թV���Y���G��A�||�R��!2Eg �����I�*+<��X�3��f�&x�jf�wx�@fL��Sm��iTw����z�,|��� m�N��A����aي4F+��6����4�(�m+˴*��9X��l����Gp=�r���^H����\�ѲS���MJuK��? ���VHaEjh\̀u��;�����.Σҽ�S�s�Qz�4�^�C��`�S*��E��g8T�T�:�

fiu�a4�*�����汨�'���u#���φ���:��a@bb�ז�2�]}�Xn�N|\r`xJ�O��I1Z���,�ﶖ����3��pW��2�a��b:��&�ry=٘U��u�O�}�G�4L.$	�o�E��u �M�_
�9����bv���j�Q������Q6�����8{�;7�n��/DP%��@unn*���Ml�<�4�m��zM�L���|�ǲ�����щ���!;HwNt���SbtsH��X�.�?O�I�"�Qx�	��U�"�".�t�+N�T�E~uĮZ���y�A��/���A,�;A�j�)�!w������!�q-�,͸ ��j�������,6/4"3/�1��診�v�GY�W�|�YHA�Uy#����׹,�ex�%.���D=|)��L�ͅ]���I���M�Q̈́��E�2��H��[''���zP.�
�D�d� ^<*��]��'�"���e��9n3�'�hT�%�)���5�P��[���M{���ۙ��❖d�7��/�Ry��1�pa.ט�BG�y��0�#-er��d�4̽�j:]�Z�-��4j �oi
� �����ܑ�`�h��C�د`O)k�H�h��M��AH� �����oB�r���)����&Ɛ-�{�G�s%:�%:z��V_��P ��{[\ڽ4�l�ȇ�]���~c��}�]���q��7aiȐ$����C?��,�7�4ץ;@����&3�4�z+���EE�T�T���[ �v1g@��FI1�A�a9�Z`·�*0�aX��cR�����N��]�	%�?/���47U�|g��{3B��|C�_�}�$8GC�ٯĈ���ej[�C�ݐM���r��l�ź5C�ڀ��o�ƒ�R�r���y ��_D/�ד4|i
gX�DL���l^)Dw�����ٻ�B��������rL�v$�ox�b�޳?�L4$�$���L`��A��#���-}
�{�e����I*"�����^?� ��Axs1O�DA���@a>�_�iM+���)y�t (qLU[�N�Ob�8��tA��6��%��3~X�=}�8��h/���Y��j��v"#x�"���Dg6��mpsg3�ٴ��]N�v]v��b�g��j��Գ�\�XE�$�7��
k�V�1/*z��n���|ߝj����97��L���m����p�j���8�l�v��C�{��[�(�v�Qw�h֗��њUA������bY0GZ��_�2Z$�`m��� ֨=. 0H~2G��Za�]=i6����7�	�=�>��ݬ��앍 5��i�v�>3�C啕]�XQ������TP�^�N;�kwi9�c<�kڈ}o�x�f����ܽG|�ѹ����48蔘�XL@���6�w����Ǭ��l�>{��G� �N�PZ�:�g#����L!�$���ը�Y���&FH��)��.��F�%`0HL�r�r�;u���VD��4��^\@q�v&o��O�/�(�>y5>�,T�LI����|�.�ɡ6�,,a�}��j���C�R�&C�w���k!�jk�'lziDii�x퇡�u�����I���2<����;���t�ƐR�����ڳ��!�{�6_�BNNs+l�m�Wj��P8�;�6�۳>D=���C�(&5� c�Zu+V��H����{��`�1�ύ�_���.O,3�}�쨕�wz:�${,�XEO��z��Y�׳���?6s�=&�6^�_q$��%��?v�EzC�s@屼�=��S��� �h�$ÛnKS��k3�4|ql��μ7������+~h}V��x�s��u����xm�AmDCf԰g�.M�|L99gwX�&�#ɺg|�T�v��Et�L�>^%��ۅKD�'� �TN]pP�'(9Х��c�$}|h����C0�3��g����r�fu{���m8K۱'�o9�#��N(�E( �qUC�2Pv,�ٍ�I6���Q*ܘAu,j����Z��H���x�K>���( S{$�U��6�\�+��9�>׳=�-8g�����'&t2�_��� ������2���^JMy�Hlf�Qӣ���|���ۡ�׫J�b���2h!�2e�mx	����ȫ��$s��RǞ]���{�'!�cs(���
]Z<��V��U�+�|�@���Z��������1uƩ�H�b�q\�*��?�Fī)Ue�\�~L���=���=���7��]9�|�^��t��	��p��׭p��Ե��,9�Hlg.x>(C$>C�W��8(��"�^9Z��%�)���[�ot�I�Dy�,OaR�i��eD�����c��o�j�<�K���oC���:>zl��#V.�R�_�	��_{<����2���w��EO�|x�>ĭ���g7JB��:w��8�6ća�ب.G��_r%�A���pq7��]"Ѩ�^|Ww���-�P��@�He�14���e9<MƸ�J@�q]��V<��w�����a:n��������u`2�'�~H��q�����eT����c>��k�<HE鼓����$���k���M�%f����z�Z�J2���&
6���}d�u�y\���c?����\kt/�@��XRP��-����[�\9D���[��|_M;�a#m�w�Hk�Ip�E��Xe<�;�I�_i��)�Ll)��Έ���]{UzV���`(��#F��.�1�r��{tw��(@�x��d������9�S�O�ۢ��z��$������o����ü晅�����9���g�=�s�?��r�qt��iuJ.�Od9��l�=�.,YqT�O�]�����_!Q�D�|�՟���2=���ֆV���Vb��;z�>K�nSBj��Ƣ+���Ɇ
��@���m-��%�F!��HX^�oG�|V�����u�1xh@�U�ݏ�D��EVb�Ui߼7��v����2,��~~��@��-�EHJ�����I�����߭�(B���x�g^���R�N$(�N�	冸/r�S'N��(X:��>}��N�ZTʵ���7}��|q׻ v*qΛ�[��k�N�I�O1:i��U��T.����i�-E�fБ��h�`_Q. -����t�7:r	��AbX�o?�l(�4{a͐g���搪����qd4D,�]ɧ_�|��?-`-*i�������4�F�,0�]}]���6����v�tK��tQV�;Ɩ�������[<;C�=��~c��{�`���0�r$�~�v�Q��s�|[`�	
�ϡ����nJ�@�<ЎX5�1}�l�B��|3���t'P
�?$U�kl��_b���Lk-���E%��["�dL�<"W�6q���F �a{�YT'M��L���-/�%8�(R�V����׃��Z�g� b#�t�-��:���OAu���8V��P3�U��褋��p��aZ��d^���=b �ĝ�<n0RH�ÿ��0�v�����p\.=�=\�Tb��~�#�� ���n�5ǘ�o�ۜ�=�u���C�3j��F-5�޷��;=*�#�[�":d�{�)����Ŏ�n��˴�D�|��y�zl�U�d�G�!ڗE~��3$OB�������}Bd�S	&�T������"��> i/�@�}Z/�g*�x~v8D�#mgE�4�hG����=�F����0b�.̵0���ǌ�mq���R�V������^A;,�j19�{K����@��Ps�����no��H����W�dd�N�b��Q�Lr����� ��k���<+�8H�Sݰ�G����ccu !!Ȇ�ψ��y���D��1;�=S�Q����G�L�dHcs��U8�;�+N�uM��NB�h�kj���7��%�6v0�e����gp�51�L���b�w;4��$�赬dƦ��+�;V�U˾���!{.�ܹ��������`W��c�lhn��|��R�kl�����j�E!�������VBh�"�������p�9��dw�mJ����F���vM0���֘���GJ�6���j�>L�غ���習�}����2KY�@����s�e��O��FZ�ol��)À;{�+��R�����1����y�`�Z2�:*��ʺ�PB[C][r֫�D��B"��4�İ���x]��x��dD�Q*�*��K��=����1�qG/Er�Z�g)�<�W�����K /+kЪ���l)
��4���)3�_�lm��ٮ:�a��� ,�[K���Py�cx[�B"b���k-��7��^�m.B���6�<��?��LI���n�j�w���W3'��Wl��w�����c*
/��2$��=�z�6�������\;�C��շ�ۘ_&�`Ĝ�0t�{��e�]�����W��)^1:bacN�ZÎ}���#X�ֱpϙ�
j;�a��Ը�u�I-���+a/]�O�V�F��\���_���W`r� ҂�Dӫ%�"����C���;¨AT�s�� u���#"_w�ߑb�N4`���̏)����<@���@�،E%���6�1/d��B�[2��3Y���!d��9,���4�L�9@�u mpK�`��G;����%G���|�L&M*���c�-|����5H?�a��
�C���j���cg/�pա��p!Y�zip �`!U�5���"͟���P #sw�]EM����(��������(p2l����R�ru��9��A����n�BS��C�ίx�kG�Y�,�%+p�+h�qf^�Mĕ��L��K�Uܢ�fMn�
�"Y����z���ܫ������귭�Y�N��ƻa��:�/sz�@��.%����+����AŢv���ne��D�pt~��r�86lw.��m����*�2N�V��A3����C��+��´��ې�}�	 �7���0�j��|���-���'h�z���DG%f�:y�J�G�Sh��j`Cu`��ŗ(�,��DG3\�琶7�Q�-�����L_��My�tC��M6)]�p�u����;�����\�tv�V��O����-�׫f(�зT���}�UT�{|_��o$A�C��a覦��!��K�K�W���D��K����k��5뀃eV�R��9N�k����>$Sa4�I�&�-f[�t\���!�����?�Wgx!�k�d���PGG��͸Yl���G�v&?��B�?~5c]v�~�	�3μ���ܘ=QRx��?�i��,���klJۇ���e'SQ���^���Ȟ��x�[o7���i?�hq�N�0��M�'�?_��Ƚ��s؏�5O�𽛲�Q!\��G��ݡGR���
Z]���=�(6Ċ6���[�"��P���~`7�y���&g�#��,��<��������otL�"4���@FO%F��:K��`�;	����}��*�b��G'D��U,���v���7b��k��AG�b�|#��<���	u��0~��NX
EDou��V�ϑҔL��4<A��@�"c*D8pzu�ax�q=�B�^�+}�^�vd��Np(C]Eʕ��G�
�����[�z�c��G�~E�*żz��y���Y���3���Ӿ 	���R��3"�r��	]�Z]+}:��B�+{��1;ߺ�_Tn�F>^�1;�R�k��:�ؐFrޕ��AS�-.����go4��W��z���w%'D��m}���>���|ӚE�	�v��_A�Q��x�Yh�����j�����?�|^�iF��m2鄿l�����'� ��ms�zK��֩n1m`|�]R�
�v��+¥��#��~I���Rך�!J�Ђ�E$�3\�}���b]�����V�ಅ��ye��[E�6�d�	K�4�Qb'��[���B�ɑzjm���ʑ,%�����jzc$�t�JMus��_(�\D\�|�T_T���\��H�����7dH�+������:yW|jz���SNA$�,�Yb�P�4j�H�̣��- ���������n4�"���L�]��#�h���f���Eћ���[)V�[�}�e���{`P>�H�+��J�5����z��;/���/`������j�G�DՅϠ4~����k����w�1�pe�z�/ -%W�Z ǁ����S��|�	R�D.g���ͤ@7��kH��YF>�Yf�ו��+&�{�Z�8qs���H`�,�=�L�h��.n��O�E�\��%��yߌ%=���L���g�G�k����hd=gi��h果8��\���ج����u}�s�j�Z�eN��k��(n���X��ɢPb�TT�|�xt�3�"������%��,p;���A�������,�e�c^�]e�B��6�����:�;��h�1A3�� ���I�R���	Br��&�}8K�H? {M�`���.jmΰ\S[�X�r�SY�*�4�_'d?�z��D�����������,�_ ܸ0m�'�Nj�_a�M���!����9�;�m�����ή�۹
�z��1��rXH���+j0�����cV���@�H-}��6a:\�k!��^��� ��f�3|�	�kh�d�	�,�mX�ML�h[%�֐0�7OӼ\
�}������2�GhF��^�a�`nÓ ���EW�9>Oi��z��o�(�����:�%o'���	��}��D����5��K�/L�C��Rf�D��J�*l#�#���Q+M�OrI�ﮝL���LD^�)o�l �z����k�d�x�&��vDI�@��'�h��ܿ��M���A�=Ò��DM��+���Jq�.�(u�f��b2]�~�P�q���v����np"���Ԥ�o��h�~S�(�4q0�llW�[���S�v���uD���7�����S�`�iy�yܶ[|8Ύ�ÁW��Vdlq�����\j�l�Y ���B��5i~����7�F�|xqo���fc�}\���aa��QN�����Cؖ,�>��5 �w���(?Q B�����y�^7�מ���Zq�k[���mߩ+$�c�o�]���*�EC+��RM�@nm3�).~���7�������߉�M�!��i��ix�%4�!�W����}��
�7��g5Hկ�×�wH������iu~R���՚ʁ"���5Т0��7�,F�bf�%����M���(��b���ٯ�sL�o<1.%����d-����~����b^��0θKK��bT����KM�������%��f��q�j����k� |:ĠT�#��?�%�A��5:x�Ec�~��l6<]W\�e�~U�7˥~��])��p����T��C��9��O�oEǝ.8]����>3��EF�h����B�� �=�M_�$�����#�#" �ED5��(�d�h��y<�7b�
_F��d���|4�����j&�V��oʽ�(F��Ɵ�6�y�ra�D�Z�[� � 4�q\�r}�Dqk�y�c������f{��U�O��n�l����0_۵���ư���{����.�ƚ��`ɩᙕ������M�jǺo�:�>ۄ4��8�a��p��ś��$�ix���"��S���B�����A���~�81[:	�Z��gtNl'�rNS�E�\��{����*D��Q"�6��BO���sfG��: ��˄o4��r���[A֤�Jyo0�Cm{�ڊ\��M���(�k�):�w뢈��P�Q��<��KF읣L+�8l�[/T����õ|Ȳ-"N��_�,�ǩ�gΕ�w[�V6i���M�&0���9�<2��k�(8&jK� �S�A��2ډ�C���7��g�*�%�єu@�|��ÒF�
�\�	�Ӡf����_ EC���&I��� ��t�e���x�1���m<�^D3�u |Z�\W��pW���͋��.�l��V����6�v������c6+�ǒ�ڿ}�wD����W�N0����d�E�)c+�Yg� ��˚�����%��_�@�^kwof]O��^8oZx���%@E�O�ܰ����|���������°�#r�
���F�E�1|�p�F��qDC���}��N����h�Ԫ�����>�3-�pPR��LN(Ku��՜c\QNG훉��6��6%���Z;�C��R�!^N�D��Y,JWŧY�d��Y��&B�.�4�fS�[�����Ak���#v �}\��u9��(q�#���#')\���Эxi�eچ8:2�2:��C���w��@��,}e�)a��`A�Sؖ⧉ä��ߜ��s5pw���7�Y����3��p_K!�ȼ3��3�_��� ;喧�-%��/������C)�@���k��^�����H-�"�eu-�� ��P�d���[�5�ɹ%G0 �Z�=�Ow�-e����+������5��Z`U�)����6eW(�{�8թ��W�8���MͪcC:=3\^bƸ�8��H�'�w>����[Z2(�q������l�Bfs|@�5C����.9�HUj3w����+9�h9��.�J?�?�K�B�F�Y�iL'"r���Q颂>�і�����'���[����y�X ������2
�������aM�D����vw���4�~��n�t�;b��f�9~�/7��u?�P���w[���zx_.� o�s7���r0�NS��!��s.�!i�(�0�Q��z��f�U�j�y�W�.DZ�����v�}��s)�1K؂\����<�+�/���X�ec������ ��+����RY�V0�n1w����W��u.���,[�3����&ʌz�G"�g�����sz�M)����؛�4Ŕ@�-��6l����_F��I=��U�[5���D����z�@���^	,�U^_wKݬ��g���1��![j�����A˫�^�gϚ48(N�b��FGW�U�
��n��n�ʼrճsc~
�9�7�0���2�"ۄ�\�y���EV��#���˷�;`���l� ;�
O5�gk\��+�
���Aؑ2���)7k��{J��Y�����~؆��h�/�~Z�(7��±w|g����ȁ3 "���i~���/�L��t�Fq��f}��Y�w	~�`�p���W��x�j1l,p':tj�`,]�+8&��/qHxC����.te<�u�A% E?n�(`��P��*�cF�j�����/(�wE�g� ���z:)���l&"9H3iW��,?�lK��qy�#c=���Q�9L�\�}�R2� x��l�,̵ܻ���:��nn?�z���J}�R�/j6�Zfh�/�e���O�]M�!r��9N0�jWaz����M��c������	ޥɢ����-�S�V&�?��H;�_`ɚ�]�j�h��r��<�PN 3�0f�����0�t{�����(M����� ��|���Y�%����r��}�_����M��@��Y�@�����:��>�����%�GS��pF�p{)�lq"[GRc�����