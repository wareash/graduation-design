��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jåا{�\�u�?߷�dn@6�zf��r������;���:B��T)�U'��+��8��lQ���M���8�ߐm�;�Ǎ2�9��d�w�!��]��*�9c����ޚfW��0�H&<K+f`��>�ȄV��N�:v�ߙ��e�H�P*#��[���h^P�ZrS�r���#v�P�!W�"���5;o�%H���ΐ,c_+��4yӹ�s��%��=Ů:�/a�x)����8Ļe�>G2y������2�q��Av�; �ݧ#Sv=�9����[2��[�k �oH�0��D�6<��d�%G��ꕺ5��U�Pm=�1���$e��i��@C��%��t��D�Ҍ�u������n&>U�ӑ�*�D�.��Ͻ�Q�me�\��qT�����m+�Nst@�iu�:�TM=˓��K��{i�����S��G��Dۍk�ЃwRk��yȑ��=�	͐�d?��}t/ΓG�- ?�	�������� ��l��閝O����4�+'���K�k�[�]����lwd���8����k�� ���lψO�����L��T�R��O�r�˞D�o�^�G�zUn�ƴś>
PO�Umܘ*F'&,7�$��=KB�j���5�1W`a�$V:-B�ӂ\�]����@s�"�CV��]��q��+N��J\�W
���j:��c}���	ӵZ�E!#����Fg���vn����X]$�	%۹��I [�[��F1��r��:�	��w�H�"���իdETQ��es�r�����������Pn����%P�o^Px��9E�Nۼ�+g���LX�x�ۯ5�SE6B��ğ���[��k�$�D7�����">�D#���#SD;�8��Q�H3F����E��Zwz֠k �lc�|�ػ�@�jx�M��5;����`~ɐM&+zg�}
�"�	���O�b���$['��@>�O9Ewv$1%�H�D��F�a����܄��sA��JW;[��ۨ=i��9�B����������\3q�+�Y!��-~��e�O"I� ��|/�
e��-en�БQ�7��0r�x-�ǡ������C %�9�Q]x�N��&Fy�J��
��qHxr.P@en�XכzdybC�;M=&�3�"Et��Z�-̘&�JNs���}�#��I�wfy3�MB}����,���j��)�BE��/B(!��pU�m� !����,
EF��z���=�]���
R�!L�Ms�Kf8̭�J/_���]�"��ђ�z=�*�*��w��~���:�3+`jJ.�Tz��C�o��l)Б�gw�)Yd3�z�o�#�L�3���8�"dI��G8�]�|^k.i��3�BQ��t|,�\ۙZ�H�r���Cg�e\�D��@�09`b�w��W� ��nE`�Ub�C�ދ�|kGf�:�q���"z·�Xe U��K�}䫮�Ν\�O��bDC?"����j8۪���Ivo�e�U�g����;��:*&�)��Sd@���"�0�b��w����U�6e#=.�{�L`��������jc [%D�1��U�i�=6�r�Q��?�ˮ�;�t�HrH�`�)r��&�,?�U �u��HaJY���3~�j ����P��	�S�ɼA! ��6��Ȕ��6]k��ې�h�dqS�����dZ�A3���廔�|d|��)�������#I�\&Z�M�<d�K���q�H��n�x���ǣ���/	^��I?��9���,��j<W�� �ly�-�E���2.I&� ��`�ک&�$O�a�z��t��}K^xs�������x�d9��O�ޮl��|N��|u�m/� 3D���2�	�S��{:7���1�ð�,ߦ�/���B��h{����9�BĨ�8�� o�_^�v~�?���g-<H�������޲�e`�lcH/D[��ݱ��u,б�X�WY��^��]�?k�k�|?RJ8��@����,h�41��_F:���}��Vc����L|�G��T�%����᧘�Lp�3a��dU3�F��t�R'�^E��r�l��﫴����� !w�y�2����g���V��!�&eXK�,�]\�������aeҵ�4�j(��	��$�g k�`�T��Y}�����`qoda��:�謐7zfǒ���=��Vi0�|e�������2Yf+*c�� ��ή���<�l�6UOa趐��K+��ɝ��B�g���Vݒ���M�@��~�]�����98}}��������^Ј�������#0��X�b�H�A�#�������w��N,���d�F�P�0D�}B�N,�X}-PKu7�M�V��ҋ�"g�Z$%�59ϳL`��",���d5�Ƌ����-We)�q�����=LEg;9��`��6n`]!��#�"]�䷼�/a��;�"�.3�H�e}{�1��Dl)���xKn�7�U�2������yX�\�X�6��~�=�����k��1��9�ӡ�\�'E?��ƜE{��[��u�oD��Rݠv^��H�xQ������.���-��~���wb^EY4@K'�?��+<֢���@8N�3�k@!*a���#Q�#�5�;<��??� g��#B�k��W�`!�e� 8VD�u�YI�,�-b�%05� �M,���T��W�L߼���4Ao�H	tv3�x��:�Hi	l0O�œ^e�'���'G�Pk����z���bЈ}�������H��?V��82�!ѡIa��#k����~�;�� ����L�`�b�o���C����6�L�!�}G-�	�W촐!�XC/�@Y�j�� �� �J�3�^�����p]}酛�6��qȏ0���3����H3���]$��af'&�`�~�A�K����ݭ>��(2��/��t�A�%c�k0pc> 
x�L��EJ��㣈�K�����SM��O�ܰ� ��D#j�PI�!���' rp��R_�W�S��3���d��qmBfmd)�M,��[��FD�6�К���DH���
��dX'��e'A����h�r?���UXx�*�t�X7��\��ls�����9����"R@�a�%��
C�3�e�����v��ws��ke���g��1Z�u�()jb��!�;C;җ�*��74W���4�d���N�^)�� �����ͥ����W0�Rt燐�
I�]_e��Y^o8�̇�E-��)-f_��&źi�p���Q�R�� ��I��Z#R�>�i�o�^O$(�~�%Υ�sx��P�z� ��l��~���&^p�����0Evvu���������œ�:چ-�Az��Cs�c� 7���5;*S���(Dl���r����7�ŝK=� ���X���Q	��.zs�����SS�͗�����.��[߿Nb)���;��EŐ�t� �.����:&�YK��7f�R���S*_ �vz����-\�&�d{X�O�Z�)2���1��fl�����^{�Q?]����9h�Ƴ&�ϒ��"jnCP�K��9|�w�� �><-S2s����W�S�8��I��&���ǖ��~���֟���ZZ���e��8�o/O����6��6��B�9C�!�N%&29b޽��wO����xG{�]ĘR�5ǁ,��C�g����A4I��(:#{�9�Z:�3	�f��v��:d("ԍ�	�w8 ?g��UBu���UT��c�r�N/+EΛ]"����*D���R@s��9~}�}�?��}�ܕ�Q�t_̻p�~`���؎���ne��&��K�MUe�(�6�j鿚,_��KxK��.G"QB��;j�<�y��T���R�*��M_��6��q�s�ё�AǴ�	�\�<C��T6��p ��7��Q,5C���u#�c����,�[G�+
=�ytZhl��l7ƦL��ɟ�'� 1Gk^[�$u�UG���&����w�.T���8B�0T��=�r�� q<���g�;C��l�.��;%�j
�3!��rU��* �Y�/�r��h`��$ ����ւ���������Q�5 XJ(���jc��=_�ζ���;�j�E4{�016�:zD��BP�%S�m��ߑ�z�\��
�'�;w���)�Y���
��G���^dn(�z��re[�	U���_�Y�:�,��s�x�B�P��0�����ƃ���t6K����wj�9?�/-��e�F����o3	YÇ�l�&��Z�w��Hʹ�)?��CC|���a�À��(�ASc=Py�n�-�e�?����D)�̥]�W1̣��.Q/�XtW����w�:;�ak����Y�T5��2`ۮ��d��D83,h/v�hҋ�C����q^,g����mW�Ue��m�ƫ(P-xU���а���o���6AHNp�<��_CN�.29��4�G;|VM�	x�֌�r�8%��0�	�� ���J<�`���<f�e(8۟�B��2�@�t�6�O�����?{~Y�R;|����)�I�6�RJv��#�㜧��9iMN���B�cme�e����c.�`�pH��cj8KDDk�P,�tF����e��2W Nz!��e	�D��2�m)'�&F/ѵ9�\T9�m��`Q�(Wy_c�i���ҳ)��
�H�Qw��`�*�)�R����@y�Ĵ3�Ƿk\/='��7&�K���|!�@��U�A�햧�[_��ɱB�U��d�}{�pT��;NFt��񋫧'pH������~��k�$�a~x#�
��O�.`.n���K+��k�|�S�IPq�i6%�����H��#��3�G�_��y�7%��D���ŔDx�
H�(Ņ�l�O
=-��t������,���3�x�UZX���3�b�ͺ��\��a�[h�)�*���A���,��|�È�U�wu��x���4���z���uf6HxU
��h��1����t���
{��������!W����H�(Q�z!n<*q�Ϗ��x��%���b���ՐStt��X
�8�i�g�-�StM�M�d#:2l�(�yr�G::A�u+p�ť��K-��<&�櫳�KA$�ftP�o�r9�JAq�C"O"\�#�'��Y�ѕ����B�����f����D����IQ�n�-�B;�D�3V3�K1)h���`+t��]�mI
_�q�D�R^�S�ٌ�;=Yw�~��ٝfe���?��?�Z&IQē@t)�����C;D�_cJ�F)�PK�]�q$Z�;]�k��e#�u�Z /�V�[-Ӽh���"��қ-���Po���C�C.�hň��b]��f}�;��٢��2�m�˃ �K�J�E?�ˋ\/r&�OS̋C8:+�Ÿ�g7�|$�+.`폐������=c6bToJl��6bo���/��I��B�e#ls�!R��I�:�5���(�l�C�ޘA�����4F5����u��?[�>�0�f�
|[����X�)eM�ߦ�'浾'@H�5_Ґ�fx�w4뒸(d�V���Db K�'�����u �&�;�$.�^�v"�I�; 8b��6�<x�
+�l���c��
�,�[p����Y
���)#�;�����{����:����ʻ��xlQQ��U�i�7���D�������7�[=��M
�{Ⱦ^��Xx�a1��`��RZ���V�M cOe�gz���]��f���k���ۋD����\9�񷐬�3��a&䃌�v>}>0`�	�d��mO�V¥�lZ��ax��#�61�L��Ce��7���J=�"@��+q�}�AO����TL·�|�Yg��~�̗���r�첬�!B*����>�s#s���\`L�7�ul�2� ��\	����蔳ɹj9�T,6 ��A�A�����V����������|���kM=;� x/O�
�(�Y��^��� �{�6~"t���\���v���ΫH!�����IJ
��C��������6fp1o,�>�{SP�=!+'g�b�HҶ'/t4�H���u�I[�{�Բ���P�ݭ?�g�39\q��5�vK�Ett_s�tQ��[�Q"����w,���B�b��2�*6\��o�у���/1}w-L�E�sr7\��kF���w� ͔O�H����
H
H����qύh/����71�9K"x�|�/��~�|[��vg	��&�q?z2`��Yt�I�pP@<�g*���C���ɀu�2:S���_X)��`�b/k��n��Q�i��j �Z y�m�Q��T[�YnZ+ GP����A�A�;��G(��{��^����xEt!L�Ϧ��܇TfvR-!�l���s��r��Y ���p�!WF|X�hCL�U8w�U�Ư�s��{x��RKT��\�O�v��g	�:3n\�������?�1��;��J�_!N�̋�'1����&��OG���J\�h�UG�Z;��,{�-0���Ҹ[�F}ε��S4�vXw5YVS��2Z��R��7����`.�-����R�!��D����e�����ug���k�H��#�K�cS�GCa�yָ7�6!���9��i�?p�K4�-��1���Hb1�0Uހ�Ws��f�`h_�m��I�
���� �Zg�N�d��w�3�	w2���hG�/ݤ�*I�H�1�n���|A"��f�V�[��C3#�� �wjș�iָ�]֌R���v"}�Y^��߰xr���2}�t���(�Tw��2^Y�ߎ�_N7mK?���K�-���wQr��%��piF�Jq�62�����/���d�n����ԝ������z���9���|���$M������BYx�����Q0w�&z*DA���+���=JU��j<�
<���T�8̍�o"H�ˁ�'ZY����۳qd]k�]_�2����S��=� �qnl�!W�����.��Dlw�d���3ҡ��J��=���\�Ri8>v��L�w�ۘ�Wbd��b�	C�͏��	���x���*�(�,��o(�����/�Ӂ�}�8У��u�2וR=��Ss��ܤ��E�� �[|���TGo.��:��M(V)�$�+q���J����BJ,�[��uZ`�:�?F��|�>S�9O��d?p�~,���jj>}���+T���4��%�a&i'7�~ә~���br�F�v'�콥F�[��ӵ��=���}\�R�#��`"h"������d��Κ��k{�~a[��.�y���'�zXŎ��O0�B&*������f�@�T�r�;ʻ�n����x=w�a%�eY�N�g�s���P�g��T�GаL7.d/�A��l��� rJ�׬
&tU��Ir�o�֩�-���*D�5�5p��^��0���N�N�[���Lf[�^o������Tzm2E��<���E�<ւ+-��V�(m'������b��%�Z"0��[v�.���>|��"�ݗi��$gP�ff�>�I[k9�&��AYe#�K}'jtq�$S�ً��*�NkG+ �E���1��j�pډb�h�0�x��_S��66�U�	�p�e9�̏�7[wwr�T�讕Ⳑ��7`fG�C�cε���e����p'�A3�9<`�H;|�\��|����	F��t�,�hS��q]�����	[H���z'�+� �@X�����ܲ���7���g�'��i{C�Z�33�`!i׷��h�����(N4�|	5j���g C�{p��5�?z�����aq�
��hMZ��x�l(�uo$�>x������8;���W�d���G�Cr9��$;��Ȕ}��{h|*���8J�jt;B�\zc -���N%Nn�/b�k��y��I����㇭fӁ�f��%�q�lb<��/k�MD�*�Pl]"v)�eq��oa��՚Ĺ ��Mu��$��'1p&��6q5��ML���[5']���H��'����*P��L�c�Ѐ- ]��}ģ�%�8�D��wM������SV��_�m�W�i�f�3�ր�c��\�d�Œ��p_�/)��i̟���Z���R@�QwƣV&��	� ��"�Z}�pjh����7��9��#@(��<Q����'i"v���]R�b����~`���%�
�����q�p񜵅�Q�6�#U�e��R�zjS�)_��K�B�����mC����>q=�v��| �љ���	�A�[��tDb�+bC�
H$J8H�)���f� n��Xڸv�S���
��A���Q�����ma�;H&�Ο��Ew{�^F�N�.�qGHD�õ����7P����a��p#��7h�b/�x�t*� �(U�{�VB�$��p��^3��չg�o۞��6c����	(�-mF�������*�&.�wc��Z �KH�W#�߄*�.�����m�g`L?�Cj6)6���x�4��P���N�|��Y,&�j��>J*����M�S�$ĈB�iR���pd
����N�6pm2)���M�u���@\WI��L�<vW�\���^I�o��摯%՛�g��C���v�7�oɡ��e��h��P�~����o��v���)E~֜����� > y�9l�e?�1��s�uj4��z�G)��} ���B�wA���Ǽ�ל*�}7L_T�d��8�f�,`A�c������� ��43����i�?�ԀƷ�X�=j{9�?�a�	�<_r�WYi9�S�(F�-�5SH�=��Uv�"e�����I�l��1J�uɱ�ܻ�0��\�WʡkGG��Y�E;���#N�K�����C�%p,eea�H��>:�a]�^8"���>M�T5��u��w_>�V��6!Yf�3j�X�� �L�����>���1�؏m���J냂��&�����)�:G�BA&%I��aځ�_��Ǽ��ѝzY@DN-����-��y�ٜTƜ��@d���{ʸ���z�1֏�~�b`*��m	_B?��I�y*M��7�-�lsг�x�!�:=FN���"V�R��_�q��E���!��9]>*�jd4��l�Jg�����Y��I�,,���T����ĩF\(�8\ya�~T~O�N�DU$���,�\Rִ�����)������oY0�K��y%`�=��o�ZIb�� fo5��z�JeQ�z�/ۙ�X�ii��f7A-�ʰ"�W��e*U�7�	���RIT�B��E��Bh�̑�L�`�8dɞ�����$E�O�Ï�ԧgE��_�{/�#Z� �Lk8�K�=��y01��_���
�����K�<V>���t�I��ǉX�v2�Ba��L��i��ɖ��m���SʾْtC��gӅ I#��v�;Jg�����-�t�I}���d�R?�
�C�Xޏ�Y�R�wqL���&�/��{�I���g&�z��h�`���_�xN�ĺ�G��'�f�&����:{�����ږ����2�C����w�ft���x��yi��1�A����h��O��Q�[����H\���%K�G�+�@�‸V���i����13q�5�1n~�����/��A�Y�������j"%��,�ܝqv=h>c�&M��ғ�a�b6��D���5�;7���}�&�D��0����h��c9o��|rA"p ��|��M�O��n��8$��򎰶�f��[#�Q:Q2�­�UI۸�$ߍ�_yBl�֯�}��|e�2�«�PW�8��Gv���-{�mlJk^s,7;!��f�-��!$��5�M��-1��C����iȁ:�hDj2g��3f�!z^>���u�~x(���1�u�\"`������<Pl;�)�6���b�q�d@���-:d^r�xW�5��C\�y��,���C�e3x��bu~b�j�]�|�Cy���|�/W�pg��'�8<�*b�qʜ�+�ƥ�	�J
�����1K� O$�9k�n��2_v/�(�]�hQ�v�.O�rZ"[}-�T�G���!��t'kx�)wQ=�����.�J�7"�<j�J3�.�Aii�a1y�hBqf�qGB������\���O�}���b�����ä;�y�R/Zr&	l�fL�@���^D�u4�	�؋���f�@�Ф�U���D�]{���Q�)3��V{(]He��B���j�Ƨq+�/���9��bFѣ��m+��I���q��=��5�4��x�t�$?�l��(�9��@&���ag�Ե�"���	��w&������3Kg/�,�_�oN/�76��;0[*k�����s�)QL�
�����&%���ւ�O3�KX�7��6I���\[����$���}����~]I�M$��we�"�r���o�ʒP P1YQhx�<��(j��iK��F��ָ���EX?�{g����N�o%���wX]:���&�z��P�] +�7�[V�ZYe]��gk�L&.�W�6�Y�3c(��+8es�Bo�*�=R��p�j��`��+�������:����g�	-���Qҽ$o)������[�/%���=jk7;	/�*�?�;�`�u�(�qndh&�tzP���
S³�mUj�ؐ6�@Z]&ϧA,�<��im������4 ��9%9�S?��m�>zv4q�q(cYÝ��~��Qu���wU���en)U�����Iv������?�q������U�A�L��7Q�a��@�JȒm:r��p��ե���fA���:����V��E�{�Rc�,�ЕN)� Y�������V��G�먹)���3�\�Ҏot�S��A\[�m��A��pW;�T;���%��p=�!�i8��!�L��c�)œ�����`�ϙ��	���5��az�i�����Z^�`��pZ?z@�U���5~�������&���s�%�%r���
?�{^�yMRs���qQ,(	���mS������Cd�%�^�{�_.D����O��BJex�Y��ztF������l%��n�δ ;����*�#/˳s�z���5݇�]��JQ��4����+�?������ڦ�@�Ic[�'UQ5;�1��A+�%���D�p;�L㠉|�g��;<�Rr%h��i0;#��~�Ұ�>�a�|�K2��N�aV��b������";M��!6��vn��"V��K�Zx�QjВ�*���g�a@8^�X@�3w�N\�i��z=���h�7�,:z�8��G��T۠�¶	Q1ʅ"R�,>"��@`�KgC��hJ�{q�.
o�t��(����)���3k�I�����J��锟ÜBbfIx�ٔrN�F�������	pp����uX������G�I�4��'Uy,a��{���U�)�M˩��,W�9�C�\x�y���2��a�-�Z%��?���l�{O	����c�^ND&:�����l������Z5G�-ͩ�FO��Ri#|Y��U�rm��Xje��h"��!z).K�ZM��5��]�`�m�w'��7��޽����.��M�[m����ɒ�{�-��O{";]plB��դ���xaQ���G{���v��΅�.�%�8Fz�8e�I�>%�	ѥO*�y�-r���Gm�̔����Y.�*Am�r���D纪��ѳ® �6��W�>FP��@X�2B�2t���e�1o�y�C���|�����rn�"��~�]�XT�C��[�ZE���!�&T?�kf&5�u�ک+���� Pl����G��K{{C<���Y4u���Wm�RLS8G0A�zJ�u���ůǈT=�7�D����b�r#,Z����m#�*fc<^�t���9���Nsm�x�3��v�^\�t���.��"��a��$�08�oB��2?���Þ����sf-���S�#-�M�&�t�H�%N������<
R>x'��Ӳ)|K�u�%W9Yf�u)&�֘�x��]��r�`g�-�@W��!�:�b��֣{EM[��	4��H��Q�Z�`U����R�zg�Y�6��R�34䐳w���6_��Y�_֚}��[��y���+K�<� ��XxGظ&���!�w�SX�M��kݵ���JA�i�Ql�.����c���I9�ŏswx�M�q�x4?@;e`=�����#l��n���P&�%���pצ,͐0�xĥ�p��#Z��j�#$(AQ�Z� ��U���v �[�U�w�C�&�Yzvl�s��Q$I��7xKY��0�EJW��cqQg�A:VD��&|�9f	�%��/������u=H5�zm?���p����T���n�^�CH�\{nV;-}nn�_M3ĩ��Vrp&k,Ι�J�������-�Y���\ˢ�Z��9SK��e�5�(����ϑ?�|�E�E#��7����}��3 y=GG[#�e�7��X>���G�<.ҩD9���Np��\���N_��X��x8��z�����g�l�D���0M��+�gO�.�~�M}�3�n��2���G��w���� Ö�xp��Ekݠע#s�v���-#B����y�
�,)�f�=o6�y��g�u\�I1�|���ɣw Q��J�fF��� `!��r����{ nT{W�7�wD���� �w�
���i�ū����sU��=��ׯ�����'�-0�i��5t��׎C�%�S�����w��1:"����q�Z�ݼ'-��2mʸ.�Ͷ��T��g�A�
L��q�0<��[��p&��9��#���Ҳ����p���t�iRNeiU^m� ﾃ�O�d=_��|�R0DF�-`+�����+;�U�g��S�e�	zy��A���B��D�L�"R�cbNPV���}���\�E�~�>�VPt�.x��/ʊ�Kc�
�B����T�;����	�oxhU���� �~Ş!��j���W&$biqo'a0���P���;�WZ��#�'��q*{��ܽ >�ױP3��(�Ψϐ�՚�h��꘰-�[ж������K@
d��f��~�L��㍱h5҅
e2B�b<�)���qb
���H�����2�� �>���4p�l|C�b��x��3O\��%1ql���6����~��|�g��ӡsCN*��\;���9�W��+++��(*ht���5�����@�B�	[�V�G�� �p��Ý��g�������	fx����!�<@A^���Z��d[�xm��J���m,�mF���T�(�X����Y���=hUa�+��Z)M� �:
(a��}�.E_�Т�ŧ^�_�ک�x������GL4�#�]�mU���oB0/�X�?f!���>}@����2�b+�{���k(�:n�&��+r4�����	�M�\�(���e�ή��Nb1s�	 ����+^Z�}/��@���o�ކ�mu ��~�s@�b d��cRf�!<����P,�F'.��jD�|{���z��$F9;`��{�mLTTCY�MNGQINsڅDi	���V9���L,�M����8�øI�a]�<�L���ۢQ�,9�G;�� ml(�4o��6��;�2 ���I��HU;���YpM��V�1e��d�� ܅b�PvB����3E���ۯ,ʡAN�Y�h"�!�^�%�2nU�T6�qS�h�9ɮ\���H�(���	�F�+��[~SӢr���StǙ$29�O��G�# ���ާ�23��rSL�qv��F�}8�����m8o+�T�*6D�u������D{/�P�$w6]A6���z$&���HifTHY�Mh�(�w=���VN�⛂Oi�E���[�B�ч��-�m��Q�gi����/sd��E@�� ���/>)�f%��m槲#(ۊ|��H���ض����o��^�DdC��qK�\�	�f}$b� el�/Т!��	�O����"����H!�,��qRk���vgP�$ڜ��w�kla�IB�y����Mߨc�3��Cj��̸ͥ�R�ñ'%{����	u��v8�H �����,�{9X���S���E$�D욀�`�@5�����^؈��X&�
�/fO�|��ے��N�O��/kC�Y-�np�Ԁ�i&�x��D�̓ M�2.�W�K�2EI��`�s�}��8s.�1�����-�įXf67.��I�7˚1�
'���Z��u�kN����xԘ���a�Ż�ǧ���g=���Ϙ��JLn��*��UܧQ�<?��ٺ��cc���f���>��/>&��U� ���h��;Nڗ��``À��7eѦ��qZE}�c��<�������B�z���J /��&���M��wm]m�M(�i�OM�ꌞB=21�`��3�Q� #?*{��-�љ��t���TT����{�Th
�� 1�W���M�����\����r��/$z)LB���L�aŭ��5�=n�̫İ��,S=���{ɣ��|�G絎��z�k2VA�x\D-gNm!ճG����Cp k�?uB�D��_�\\[�ᚆ
ʁ�ӏթ^xo+��L#����s2�w��9�;��R�(��w�ǂ
'ߦ�T�G��_�J$���{+x�c��JW�WBӳ� T��&so2y<9�=�	��B�94/�2M%�����8���A/��A��8,�v7=��)�~btNs�1h�&�0�ܴE:���`8�5s �b2��[g��j�-[�R'A�e�2��(±/��.���j״.ᶰ͉ Ǝ��䇼�K��s�a$�0WDC��[>%�p� ���)8�?'o���X�|�W;�ٕ��h�n�*b'�ƒ��CG@�8���fI'���
��Ы��F�l1p5�p�l���j���ϲ���[U�St~���XC)�u�n�T��3�|�^ޡ�9�|�YF�q	���K���l���*��)jΎ�L9z�cH�n��J�|F/�D���'��ڎ��O��s���)� �:"K���)�k�ou��)}qg�1@LSz��}���:!�O�*� ���)@�%��P�+
�uٴ�z���{;�I��olW�]�f�ᓏ9�-�������\��P6���+�zM���{�	ؓo����۞m\1EŢG���#t�*�CM�c�*�|@��O�R��7ӕ���U�.j��XH��&�M:Ds([���X��;S3��%O��%�y�!g�`ba��1������!!J�)9%T昄>�W���T/>�R%Ȱ���L«�O.<��M$�B��#��V7ӈA$����K4�,�b�:�5�s%�g����bˍ�;�\���}IV�Ey>d�2�x,������E�1m#RYp�2��U �gr��O�����m��pT�V6q�����426#�Nt���ٺ���&���r�o�l��S�OO���r����P�70vF�&��K�Ą��( ][(\|���3M�m}�Ѭ�u�bL��/�b̬�EN�c0:���MFt9�Mer�	9����4Ȇ@e�^���B���'}�����gX��w����)�"C�4*�.�|�K�f֔+k��<����LX�$*���n���<qgTӤ ��O�.A���B-����:cj.��)��:��/�[�{v�71���hA�8��B��r-��Z<]��Rl��T��+8�T�'Mf*-�;ť��ښ�X�S��ЯӐ$��F%���%���8)QǦ��X��]Rj�����M6��;��/��}�gBxd��i��Q�d��u�]8��3Z�ۚk������� ԰v Ϝ�ڽmv����伽=��9�������k�S>'�+�M
�9��w:�����3��_KI�x��s��	y�!=���j�a���#rɓt�R�J�f�87Cd�%�2��� �@߄�.=�9����耦��%<���|������8P7���P�)���'�6s�O��0)e��-׺��^�P)��������Lշ+����ñ�*�(`��H���kO��G*B-\6�3S3�.�l�5l*��+�E�V!����Y\b���b�p��^Q,��z�gg����樜�yCh�Wp���ч���Rze��S5\8�9��x��{[�w�2�e��D�9�ن�I�ŵ}\�H���WC'^�o��Ou �Y�Ǯ�OW�{R��$0�f9��17�o��"�}��c��\��$��]$��TŹ�/cJI�ى0�U�Kl����e�u�wH�X:R��֯a�9Ax���NJ�GӉOm�q�3Wl�����O��:u~gGx�h�H���٣�{5������i���i,�P��àG�lb��������(t��N��d�=���53�Ȝ���a�-��T�]�O
 �bX(��zo�
��#שN4�37�c�����mG��b��\͡Q�1X�pJPmЭ��;4�L������p?B�C�T�Xӝf�_�[��XW(j���!����p՛��䍟V7��?��ӷ	�#����t�Z���Y��:dW����r*�u�eH+��ǣ�1"�9��S���ɒtK̀�m� ���@L�So0/��@���RS�\]���`�8�Z\��z�ȣ����@�2��%�?��rZ������)�~S����5�c�m;R����:KW�5\ҿ�mfz�݂�3�,t�^�X����p�xvRQ�r�J��p����3��)�X��t��I�1d/�I�i�/f�.�o$�O��#�ԅ�������("��e���P�r�tn..�'��cO� �W?���H�>�cC����jS�q������`��0&w�5[�D���g2^!���p���N<�2%j�����-�=���r�`u�������3�3a��p���|O�7�0(Myk�0�J=
�:|���J���1@�	V��H�[<���Ic�$T9F��Ì��B�������oJ�%%����f�l���=f3)1+�ҍ���k�D�HI�o�3�[�ͨgZw��*@�V{\A.�0%��c���$�/�!qCG������&Q�94.Q�����U�;U%�-�j�5�F������.�+ws�ʻ%�5�������6G���Т{_%�\�#9s�нE�m�a�5ӏo:8���Z�?b�}N�ϒ�0��:_��H!;��Ews�������=F�l�8M�����$X4ԥKz��t_�&��`kpg��E�!Ν��>�#C�Sf�NN��E�H���D��'`ɚ!5��'��)�2�VX����Sf�,xҺ]o�[�ޒ�0��j�Bz�e�:@������.֢�G6���Z�cTߺ\p;��U�,�/�̜�)M#Bc�(Xe�}l��oug�9��r�*2��M��ߝ��6�RF���hT������Ϳ��(����E�����S�
?u3�)Bٓ˷Q�;�)B���>�r�VO���jW�����	�U�_֜×���JW�WG�&��q|�yna2��t��o�����z���X����[Y�S���X��:�o��
=�Fot�S�� �1~��Ĳ?1�XL��"G�}�VYlIH���c�������[OW(�l�CrE(4{�Hnu�c�e������v����h��"��_���p�=�"��4<����U/���Ԍ8I:%g��oY�3�};yLzp��� _L�9Q�*��j��e�g�*~��������dvգ�~p��D����E?��5�q����D��k�kD�{CB�I�ҩ�ҡ1�Kպ�~�*{�f�,��J��
v��B�N��"&����Ra�_���ܛ��sx�1|�dM8���a��`��5�d��I�dnߝ��6����	t�r�!���.���JO9�!����M���28P�����T�c��N���?]����KH��������`}��@��sk�#g������5)�T-�l6N��<� I�����jz�xD�өQ�|��i�%�cCkg���aj��)���ި%����Tڗ��0��/K���~��i��EK��r}���Z�KݎY���Zu,�'Q�(6Y
��a�U;��z���rǏJ��=�W(4�#!q��#1�y�Qud&үUuv����EI�[jZ�s�l�z����w	:��w.�]��L�}�|�+���b�ժZ3���SX8�%Dς/(08��al�FFLb�zf�֌4\A�;0�g��3��8�|�xZ%j
���W��=�����A������J=����!e�D�g��V���Pd�*&8�yV@xF.d@�4�2��(4���� ��N��4�\g�0��ɜN3�����X��6��a��U�H増�����k��7���.��x��L���H�l�rz�o����K�n�F�&;F�,�c����Ǧ����t��u5>���X3�^h�׬:��#�ϓ�	���E��e��,�eA�D�iJ{��y��Zlv�������K�a_
qa5:���]7ٺE��]%��z�>S�jXߖz�8�')�h�	�zn��Sy
���@������\�=U�y�!Ə�8�_�3��A�0`f�'Nej,S��&�u����4�f?���9~�ce(7���j	��`��4��+w{{O�s=
�s-D�*����#P�k{���~�#�6L�����c� ȭ?��fS�<��Qj&��jO�H��F�J��a�#���j�j�*@�#��)�p���j�T[�>Q"w����1�v4�Y����ݭڨ̰�ɚ=����c\�j9�ly3B��f�� o$��5XN/z]�K�ԟ��-�>yuuH��E�p���[s ���i���.�Х�,:r�"����!�TH1	�˦�PI����M�V �s�m�R�z$#����hJM!�Ձ\5j��l�j�6܋�f�l֯���i�Xܮ,�1���o����g���C�K��O'����t1��L��|�����o�q�Mx��/m�]�� ?q�g6]�0�(����o4���d/EQ{Z�����i��ڴN5Y��r�q͡R�֝�0=����.���΁��F�8s?��L����\A�Lu�ǐ��<����Uy�_�����7á���.��d�)F�i�J����d�z}�4��j���H�T���j4�a"9+��#�f⊈���bt�h-lZ�Y�����ٰ����v#v&ax�jK�z��os��p�S�U���nM�n�������<�O�=6$��Q?YZ���90<�qb���ty�%in�$�}��9%Q
�Q6�wQa�䜆�WK��pR�E��K�w�ԓ-پ#{u^�K�EP�&�#�6�yW2���D�l�G�� ׅ�N��`R��{f��C�4�;��8QU�Y(�3q��p;�Y�u��w=)�8E��r�!;�f��+ P��'/��h�)��[���	1������i�M��{	.�Ĳ`�4�b*�NO�.�%٦W�A$�E9�E*��U* P�i=���A�%x��VM��Dy`簮�
sϠ�E���ډ����*��y��ߪFg7�<�L�����ТUXհ��O)�[��`�+xH���PK�x͞�e46�n|Ͷ^<�h��}�]�ѝ��WA|�����0��Ǽ�j���e��|��/���@{)o����ƂS���C�`��UF�}�͵�4}��U#�ȟ���ਇ$V��Br�`�89��5aĤ�!�^Yw�I���~W��5�>�����낔�H���Y ��	��8dQ ����v��d$L�e��!�.,��S��L=G�j���ꎝGy����	�XMD�0�~��6`/ѭYS.�cF��_��Q�nPŷXpGh��k�!�p/���3���2�����!�R)�HY��j���ZHk�,\� �}Ih$��@�_%�R������^���c&Z���n���"�x^�	�%�k�o�����Er�C̀�y�?��ܞR���Uϳп?���1@ZIJش�9�9M-���l?���]sU���y
�����m2��f��qS��a��_�����a[�aG4����o�:��ޜv�*����$�$�R�{7L	Q9��;�(��� �	����/�J�l�)��˄$7U�mӀ�K�@&�{'r��p��j�Nm��<�Bȗ�0B�;�h�-A�.7�I�W��$�[��_�G�����?��j�?T�b��,nj�X�:����`�����P��[�������%�6�ҭ-L8���36.��b�Wޱ����B���ʾ��2�$_Y����;�j��L����1Y� 0�b��b+�%G[�b6�� n��L�cfZ*P�JJɣPp�mb���Ԩ�fȇ�c:������b��6����	t�B�
/���� Y��_������i��S�D{�t��;���l�2en�AxF%t��v�W"$F+�?��B����8ֵΕ��"�lv�1Va2Q�Q�C��ߠ8�̌���:�$t �RW��Rf�1�;$<V�8?$>�J�T�� ��8}@<^��tH7�n��֨�؏DH�>딜��P/�(�{��KC��d����q�;ĺ@rj8^2���&�q$L��(Bd���o�i��~t!~�>�:��P2~�qU���A+6x���gE��6�mp���~�#�[���z�8PhC��3�xZ$�j�#���*]4ҵ��H1\D�������I��#EU.�GV)�́��YZ|Ͱ.0���������-g	�,��g
�ȫ.������XTv�/H�����j�\pY�����Bl2�p�Re!<�Q<�P`u)|�������H�����2�i/D��G�_���$�_�Gν,�����>	i��9yE��ݦq`�߆���L��	%e�Cgz�����t�;ľ`���pd+d��=e�b"����%�E�+V�zW�8k�'
^s'o��:�%'YDO�(V��RX�ȳ�"җ��b(�~!���p�(��ß6ed|t����B v�*��I��hb�o&��PȮ]�qT���O3?e�!�J��σ����CK&{q���Ӝ�B��i���#�1� �#���t����W,f�fLwjK	��t�kڎ�2�Cص��>A|Tj*��1�R��t4cl��e�p��=�כO�7֯��D�X�'�Uݢ��-L�L��x? fG��Rq��%�甍����يm����χ���,s�d�g=:�O�"�R�qc#a��ȵ.s��dI����	�Ob�g]찓��غ�ɟ�*n�:�Q��FH��*���k�5�cA�j����ᰔr�9�x�
��xiZ��8���tu���%�iS��;ÎD�-�P�dk�m&n�By��'k�o.o�v��	G����'6p�}vS3^��ҍ�x�;$�v������,�#�j�Qx<,��qX�atV�[�K*��W0+���U����n�����
�SZ`L�D򥈩�I�9Q�_ʬVVX`4����(l!?���N�`jn��c�Wo��h� �6�sǤ�A�&M;離�Q�E�W���nU[���,e�u���.#���<lc�D5	�-�G��� �^ڤe.�HNƛo�jsڹ�阹%�HJN ��E�leցkK ��{�wa����#;�m>F�������.��h0�>�l���Q������f�Ի%�9�AѶl�b�y��tɂZ������yE)>ē�_Q�����ʧFPq��4�΂�nX���r��.iVea��N'�O��>-]�6�u��N�pP��a��x�|Bgxx+^aS?�6��ݥ��Z���,��q}#�9�e�-�@Uk�[�� Dq6���0�6��B$�Y����Y)��X���c%�L��8���5)�O�����I��Y��b�!DǇM��3V��5����Չ
�Tw�N�ʇEr�y�@-����n8��á�~R����|0o�
h��H�UD�
l!6��b4�ʒx�Ս$��k�-�W��y�S@F�Erɜ0WW\��/�G���f�3T��7&��ah����8���f�(�.��i(tI/��5X�֫:�{��U��D�6%| *���=x썉&�ϲą��C����N5y��&�7ے���<���q�_X��f��L���h��c(��[���%A�Ҍ��:��E!�?�tT>
Y���W����_�����b����2<0U~�iй>f�~C�W�ދ�>�@������P=m_���I�>�^������(9pT2��3�����AC���w<�s���LV6Ĕ6�mb��k�����	 ��#;���>Sv�G�=iI�J�#;�6��zgZ?�����B��;W/�'a���T��֩�k �����?�5#�U��zfV�7w��i * [
��Ӹ���{����(ҩ D�
�I.H���d��H�L8�~14�,}{2��c*[��a����J��	UZ���Xbd�wd8�8�5�3��ֽ)���i�j�LT��I}6ɋg�BaEy�������z2�M��
� �4$T.D_^;�;G>�͚�)�#l�o�.b�n {R���X�S�!瘞���uMF#n��^�C�o�2��yY�;���ͣ�*�u�ǭ�,��o���Km,���G��#b}���|$��*H�4�UR.��=�rR�~��;�J�%�.u8����<x�~�8Uh�1�i�j��k`5ٌ��#]��&DK�K��pR{�{��(�sm;��>�m7<X��D�O�) <����4���K�3Q�wY�z��ҠɂX��EŬɆ9`�?�	1ЎZ�4���/�U~��:��5�N�C�ˮ�Lh.ό��	qw�bJmm_�3���8j�u G�:+��l0��N��~��򍟉ԋ������*�L��U�<t�l,�c�.��<�L�d++�!��O%�	���d�8���>��Q�C7e�$�H���.i�=^.yR��7�އ���x�2Rfc�G���$G(�\�c@8�����:Ҷ����O��o�t��5G��yb(r~a�^���p)cեo^ۀF���N<N/ �f��#��G'[@�������CW���m�W��5�7��/*���!�� ��|g.����Qo)��.��יJ�?��	�䲤�w]oK2u��Q c/���5���.0D/���rk��53�����BPwl��ȃ�0���BȉF�B2@b��0�i��>��@�) ѕ�ɭ�p��D��g_��u���}}<=������a�n� ���WO�x�>>�:t�q���9�}8+kYۗa0�i��\%~��@��k]V�{���J��\�F%V�S��5=�&���x+��_�����;O��R"�}W�xK�ܞ�W�ُ������I>��Ѳ~Zq��S�zA�����W	�2d^k>��,p��E(SeHo9�-�7�R���Z�ay�'%���0��B�o�xu��M�#���Yq؇j�"'�s��+$%�SW�ޖ��Zo�,��]�t�)h<@��� s�ڷ�͞�|
f�V'*"��le�h�Đ�/�Xh���
Z����ŋ�{��{� ^�f,I�+D����-}�� �2���J	�P>���k;�B4�l�����dR�������ߛ�iSH�xǬ����
=T�YY�\0��L��aiԁxjb!�N=9r��Ca
^
�;�S���ɀ	|�a����M�V�)�31Mѯk.��"���:~Hٱ�2T��rIOlk��L��򜉬�C_���ߤTH��6�տ����)�ۿ
#�� ̩�N���m��W�^QK��p�!��	Yi��(�Ssa����Xw�"�5a�fJb�c�h}ƹ#���|qO�IEP�قHD7]�\i�Z��_����z��Q�:-o_d�k�{SZ����B���e_�a}�;|mX�Y�mn>�0��|s���;��7��c���P���42�� /�vr����Ԝ�M2td�*��A��`��ww�#d����c�ji��"X���DP��RxD���%0���'��~��pl�>�,2�Z}~?�/z͈�"�U��oR�t�\�K_�K8a*��`�ı�O�>	vU�$ܲ���BV�x�#�;�$#�o������a)<q<��߽.p������2j�tH{R�Y��Ph�B��,[,�����n�)�aD����w�L���9=l��g�#� 99{cF]Y�nX��=ӌ_���x0�ZQ}e� j�u�|1K�*��ISPw�M�ytcOZ�5v��]�RG�*����8'���������!���+�J7���KW�����牜���;��m��p����;t`�$At|�aU/W��C$�� ��+��-gJ���E)���d��x�bLyt�p�D��ܲR�S�HN�!#!��Ρ�ɁxP齊� �S��TZ�O~"��u�D}I�'�^��"�h�^��G8DA���F�&��5o�����y���nGQC%t��\������^��bE�Z$5o�Ѥ'�^�#ܣ���z�Q~ )�mΊ	�%�Fry�T��2��O�z��M#pH{Ԇ���p�\���P9�O�\�_< 1"��{���E����?a;ՉR���oQ@��Ԗ9�R�K��x�l<�n�a�E�v6t�Vo:@�?f������|�㥀��H8�m���Ĩݎ���.g�~��ՒJNg���p�>�bKu�Fe�-,9�8��Y����9�v��X5z� H�ѩ�v�M\�3��N�u�}�jl�,��5�vJ4�,2�/�ϖ���x?��#2�"�1u��U6 Ɍ��8�徭��M
�� D=d�3��R?��/�$K��@��T�g�JY��g�=��Wd����;�?f�I�X�%��l`��[��9���c_ml���w��A�P�44�V��R�ۄՑ̊)aY�u˜.�N���������2��O9-s-���G�z!;��x���,��o�	�{ܪ�R�S�ۂ<X��x�G��R�˙���P�m�я�,�b����u��%��M��J!�����)�;���xm�"N�1S�,�b�
8'w�	%ŏ{�f�]�����%�(��D�m�����)u�@v��Ps�~J�����I��7�{�f/xL~L�����@��+��w;Y�Ӫj������m�=gj,�!��n�(X��&l�fa��~�Y	nH��Y���)�i��/;g�˵*�%Òq��شQ�0u����H��cC#x�!#����7�"�"�8���{茔^x�*�����_���I���o�9��0eI�o��3���Jй��{)[5f���?�6���=NKQ��*����׊oR����W�v.~Ɠ��\ ���p��g,;Ed��
���փ�T�����B������,�s��;m>�b��mn~d�Ox�w(�A��L1��p�;joɰg�v�#��zkR�ۚ��j������]�d�a�>��)��ޙ|�[8�)*���p�.�����4!�'l�^z'��Fc{h���%��n����G�����#���iZǁ�H'��?$�hrX�\�:�)�R�:�6h�$�t;�_Z�(����M{:����
�Q�B�O]���㓈�i��A�phK�T.IRe#q�uV����É�߱3�.=�A�U����}��+�����枓ϛ����l�f+�0� 쁶P��1x�k� '�&{q��я�����U9�$��\Ӽ���f ;�3J��!Ӡk���F�S��%�,��6Ñ�z�Fn�*�J�'p�4-�H��ZT�:����v�������V�O��$3	;�g]>4$�r�*�R�]�Rbf�o-�^�Dl	w��'T	Q�Ҡ�G;_����H<�����?@�/�r��֐�!�6<��9���s��2,�́��W���S
*�?�1,h�a�̹�t�'�>1?��6��u_}UF����N���LL�����0���z��:5��(�i>���������=�׾s嶍yd��"�ꝚAg�-~6Z	ع�'O��"%#X��]�P���.
DU �l!+�p���L\�C�O&X=��S��R▬���WT�K�N��l����1l��-c����&�m�׺<���5�)(�����ou�}/S/�KN��t��y�n$3�Uޠ�эŉ!�c�"��f*B3N���E�#�����q��f,z��"O��a�0�Ͻ��P��V�(��E�S6�]�����f��(	���ȱ��堈R�/O|=VR�02���P���G��/��̋=�x�,l���e��T���eW�
�l�z\�?����<�3c�}Ӷ�a$�<s)�yb��k��t�[ܛ_0�e���Լ�)?�I�B��j�͟���"���L㞒��Е�-O�4��m1��w�0�^�́X���Ϝ�pq\�'JOq�s�|*�q;c�S�{��投�჉$2�.:�IZ���"
���(Z[I
s+ΔV*����p�c9�Pt����[tE������v�(�`'��_�cg��Fj�<�U����0��&��C4i�ZqK�O�`����Մ��v���v����(_�5N��I)2\��jC������z��s�W���M �-��q���<k��hGԌm�b=��(�L�!��0n����擯<v�9���_���r�|7�D�ٟ++!馩�� ���n]���]���Ė�(}A���L$�V���c׉X�MNd�6��{��K�nTO��$�R{�X	#MĜ�f|�ghA��^���)7����0a���.����V�H�C20��h>�k�`�+��
1�2�:{��t)�P%z4:� 
G*; �_#�P��㻴��e�Z�4�F�S�ΰ�~�5G�?��e�|�|��h	^Dq�s�*=O�P����T#���|�fdՠ�s`ӂ
(
��-��5�(�萸�"���W�ձ�;r�~��T�R��l���{s_\��| }0:aWz�u��	�=Z6ܟ�7eop:릏����uD�C,�7��A��U)D{�}�7�j��aK6<p�+����(܏�~7 Q[�>�j��b��z-�G�r8��(W�n��vILo���x����Si��XUɏOD[����	��6��L��r,do�4=�y(����g�x%��[墲d5�o&�	���9K3	,��v�J^��/�]�̇�9��(2�t4-��� �`��0fa�4?�.�\u�q����H,-�[7�R5(��hRh%� ;;A�t"
-�S��$���p%)�� ����d���	���q�q�c��>�K�ҥ"�m�@if�ى��ғ�ʮ��$�_׎����M�zj�W�/x��^���%�������т�fvv�r���Ѽ�<��|.���Ꚕ=w�a�ӪM�HZ��V}B�����U���Ƌ�o	/YZ��Aüa-c��萭Y-y�&L��Ц��T�͎�Z���.ɚ�q������6G��za͗�%�\�s�TL�.��cck�F��i��S�G�hf�{�1�Cx�N\8O��F�̗,�RWu8<�۞�9�Cŕ�'T�A_�����8����z��~���F�6��w�t�G��6���4o�[������gh��O^��G�ת��
������vM�U�@��a�N��&����L��̚�.3�����/��I�<\�l�M�%�Dn1��<!.�����K�Y6^t�xV�E��8eķ���p� Q
�&���a.�o�Q��0�$����XD��SSP��L�Qa���"��[͆ݔY���+���(~���bP�x-�>�>�=ܳ��֛����B%O�K�y��_����V
k7�i8��Q6������c�
�k�2%,���5Р64��J���f{Џ ��y+����u�e*w��\W��M��!�Y?��(�Vq?��d�N�x-��� u*"K�km��G-,1�h����)��7l�G�t�fP��X؂���.2�ssf  �육`;��e �ŎJg#~��B#���/��ǰR�oua.i�d2&���cB�$����Q��Z�x������-���O��yGh� LSW����>�x�:x���(_�c��w�rsͲb�2�m�L�V�˿:�s<���4�2�?ßv;������3�s7����9��ͬݶ\�B�1�,�E�5%�������n�=4V� �Pf��O.�~Pp��r"��u�$����v]_���+OJ����1	�6�	Y�m�j]��kXm��tf��ͦ�C� {�$�v��&�99ld��`�[A*�����l`\��$%
���Y�Κ���H�I6�F�|:���Ǔ�z�V�6	o+)M�R������3�Lhs����5i��X�����j
F9��THd��ې�������0��+�j]�%��y:z�f![�C��&a��?�����ݫ�lQ�B~	�s�ڳ2$��N���]�+�nUU-��'J84J�%��u�s�Cc�q��W��v���\lv��eOT����!�~�ea󿨼�y��Q�I�[�nW3��)br��Pt�v8���v$9U�����=�`��ߵ.�r�7�C�OG��%'P���c�n,��f�9��%�Z�����F�e��]�oO�P�*w*T͢ 9����u[�Il�>�Ʀ��"Wp�I�~Yy��!*En� ��t/(uK��~�����aS��Z-������%$�X�ݖ`\i�������?��bWv�W�rdm�f�u����/Y�?�k�> ��I]R�$�]��G�t�H����B���8\^�0k��ت� ����yI�wvƳm���8{���oYp>������=����-����"��'�;��T��h�<��.Q�i�N�l���x���-z�5�V�[p7���d�,�/�/�ni��(dڍⓦ�H�H��*K�S�~��U�޽D��ǂ��U�r�q�������V,��%}����������EV���B���'#B��	�L��W^�EF7��m���3#�"��	N�0B~Q�^
���k	+ �8(R�'�øu��>����g�Wg3>� �O�4���e}s4�-�"�P�[�����{�$;� K��ƕM�c��a#m�I&��g{�<�2��O�/�t&79���8�
<3�i�7k�ַ�l_��G�$~��+;�v��T65)�%du<��D�OW�����^I���1sԳ�.\Q���W�W��S�u"�{�_��-Q(pD�$s^�^���Ͻ� '��Ϟb9q3���*3��`��u��O>�T=���2\��W�Ws�+q���^{��p�z(T�*��ⵂ��NΞ�ť���"e;��XJ��8����RL(�;�m����9��	����Z��./?�8����g�7��"�xOmT����?����@|V��X{.��Fy����-okG�8��מ�m󇣻��$��
���4N5oiR��9T�e~��������c_[a[E��2�%�Ӱ�Kag�z�U ��0}?� 3iJDf�iad���h�������v��"��Y�g���4,���>K(�g8A$�Z����p�m�CX�֥PRS�e���m�e�t|'{`�TW����n���x�0�;���rc �؋/�H�0�{a��S�Ʒw>!f�w��Db����Ÿl����%~��W���y	�����"�,B�t����sIҰ?�=ـ6߻i�}�<�1�;������5��1!��Q���A���2�����MӐ�� �=v��r�������;�S��<%�>�h�{�0>�+�,�h3�MI g�fe�N"�"���KK����oPcG���Nvɮ??�3�e2�b�o6�w`YW������;�6�{?N��&8�
������W�	�f�B��j8�K�F��H��(v�T�-@���{��Xx[�)S<&RK����؛堑�����k���W�XX�H�(�l27�*HB�6�=K<�P��^Iy�t�*��u���:���h�S]jR��a����%S�YmO�і���r�/��݈���Q�� ��VY��C�B��Q\��p�pT��eG�ٽ�����1�u�r����3��R�0B���#��#�g��),p�Vne[iL5�-) �&/��0g �y���I�&Pk9�'��7_�n�MU��=-'s�o��m�^�E�+=�^eݙqW��W�,�:C�����_*�i���2�-�۬�E䩣^=��sw�Hs ��¤����d�%�4`��P���7[����n�*}.,��V4�pB��o�)�%�����6@�gÕ�$�P�bfhq�ImT�rڈ1�/�n�ӌ�b=k6����;x0����vY�"�"�u]��`�+G1%�:Z3h����e�35s-.�РO�� �M�@K�mX4�o��h9��A䝦�\W�* � ._���~���k�d���`�֤�{l�6����n*2\S;�I�=�e�p���u��~�����^^!�e�d���S+���#��[@����V�o����++W��:�5��hshsq�d�PhpkC����n��d�zl�7��cw~Ǌ���'5��g�2�*��iB���/�fHBl ̤NmGĔ�����vS�M�ڇ��i(�\��JӀ}4z��+���M����	Or#Ѐ�Ңdu��N�����X)�%�����'����r�[�@\�nH9ѻ���#��_��x9��Y6
a�/j{��?����h\c��ꪅ�
M����b ��A)I��뒔G۶����h�g�sW�����`�=�N��K�$vvl��<�qؓ�O<��y�d���tc�EC)�p�p��I��v�=G�+��K�i�.��T>(U�>����T8��Q�D�N�C��:L3h���Ή+�+{ ��.Nn�$4�T�G�,yOV{��� �Sw��6�^���k�GF���HKVN"�֐@oϫ��G�Q�#b���o�rL�CZ���xF�qY�ۀ�Gz�5WFZ��� ���V�1���3�'V�v��`u���Sc��>�߻�%x��;��պJkLq��N)�����W�EC��c<��\���+�y�@gp��*l��Dّ��1���3FBo԰Tf҃�'�ih�����amYS���g��k
S	m�:���xI8
��.�'
�ۜ�)��u�P!�~*��z��v��͝���K
Zr|��M҄s� ǭr��!�:M=�"Pϒm�Y�NVx��wb�\"{���G���T�Ǯ�w��������0ȡ�nh�iRV��i6����Q�c��T�E"�?��}�ޥ}J�n���q���e�0�����9|D�?z��#�%>�;��òF惉��q9�����.��w��Q�&>�b�C�	�B77�����ob#���do�x�"��L�\.X��344'�� �و�h�ǐt�;�.�S�?H�.>dGl$�`f�#�g��e��!�M��&�F�T�B{�N���:1Q=�Ύ;jAA;�"��"��!�\�!%��D_=��Uҧ�c�o�j���qg}��""���;�,�#ةC��/�W���j��;��)�S�Q���Y�r�xo��atr����iy�~�:�ţĝ��$<��|�ڻ,�5]�����9��݌y�ӎ
�w�R�.&�9�%�(�0@�<!�#ކ�'��P�z���� �y!z��|�n��m�y�9�:g̟��"�ݜ��$t�ͬ�J��5]!��sާ>L���b���Ԧ��������m����mREb��Oe�VX��x��NB�U1����v����n�#�v��S�z˦��)�	���k���4�v�w����L5�.8��zQ��T�~e��S��'Ne��H�h�tI4�|�Ʒ�iߝQ�yI9Uj����Ah�Բ,`�V�*1K��c�����e�y�#C�>�F�o�б���AyB�C�*�f�ȼu}�M�~����W�����a����L�[�:�C��W|��V��Ԥ3q�pĶ&�Lr�|��L�\\��!��D��.�xL��?u��������i9�>���	���$1!��w2���C.�|V�J��p]
��ܤ�3�g�=�J�BMI:����k˸?�A��u��$[�E=���*:�0�
D��yZV���]�Уn^�'RXTY��^u_d��"*���W�Z��34L���(���t�\��5�0���T���Z�J󶻏�����[����-�����}0��m�����I�V��Pt������������<7�g1D\p���;]�od��b�χ*p�2k��Z����ƀ���̆>��.���0^��c�T��BD"`>�h.��yӕk�`�M�r�:O}#AwT�W��^y0��Y	�?!-��M��h���T�)_t�`�v�2��T��>.��GD�r`l!�Oۃ��s�L�ϵVw�'��Ƥku[��w�4��ʞ�Gƚ�L�$|Y��0��O�	5'���H��Iߛ�O���n9�g���s4���T��Kbf!�)����]o+��6�Ab:·�۫�{��3EC$�F�Sė���+��T,�8.��gI)��=����53?�G����� ֭�7k
�q�����.:�̮���\1^�an�$jf�`�?m��[���Q!]-`rʤ 3o��rФI��*{F!tr;>��P��Ս1��|�l��k��p�����d���	T�����R��0'��.#~&����Cue���+}��� 	>������c��)͙�0�j6'�X���4S�Ÿ�yS��W{�R���:��74ߴ`�v��Xf}�7�%�2ߗ�	��y[����O�J9"�󼛮{�6Q[�Ӝ
{Z�Y��k���a`l{j���j����@���BF���{թ��K��1'�����I�e���o˽��j1u��RW�Hz��S&��s{�3���iUG+�6|�R���Yj#Z���^���x�ǝ�$�A�y5h�i!ҹz�ʘ6�&�W��ڬ>�yC�A$���+eh�=�b�����-�V����f�
�=����� ��)m�<��f��?
�Zc��ͬ���L��a�EW��W�w�E�*�<:�n�TJs�zHYk$!~Re�$���(vj%��h��.�D!(�̜�ퟴ�9tLE�P�8P�Gm�g�J|k�y�_��2G���I^��c�@����Z!,G�ܨY 8x��˒�0D�Ut��S'�A��ptu�F�J�>��z֌E�y����y?�Z�j;�u@�*yĸ�����6r����*����vb�<���X.Z��r=%פi�iYo�)�=L�ٝ~�M�Pb��F�k�H����u#� Zz���Ѭ��\��;e��/��-��V��\��'��q=�+�7#�����c|�����#��bd�Ժ����&M���/U��ٖ�3��I�7�],�����ʌ,7������~�Ё�Q�@W�=�A&�����Q@d�Ò��4���#�١ob�e{t@>Y��8�:�c܏$�S��)w����o,j��F��_<�H"W��oT������a��I�
���m�k�ig_��U"�q��-��LqV�)V\���p�s��?p�7�{���0����s�g<�~{����b�M=�Z��8��	��+��/N��!�ESXΰ�3���N�Y�Lu�/r�J���p~����I�V~t.��W�!���F�6�<����\��`X�����(��8ҿ�B�ƣ�������".;�~�D3����7ݿP�
�&l����|���>�M3=��p�}����ͤ(Xm]B~r昷���z�@ȁb<9��"a�d2�*%!9Vx��_1�D#�3�2�u��yR�EK�ey�o���ɽ����6�0�=��	�"��q�E��L�p�m�y� X��O�y2Q�����2����&m�1-E2Ɛт����q�%�@�y���5e*�4n�K�}Q��@�����[j����\'g��"��0��ҍq�;��*QS�W����:�q�88�ȳ�
�\�x�BA�{'!=]m6�v:!"Pmk�'��(�C�?�P¹/އ����[7�� �W)��;�Mf^%����+f�<-8�7������z���@- �C8Eĸ�m���@�xA�����me��K��%'�����i�ԥ_t~@8�^ܐ�3V��]% E�0{$hK�^��{$T&m�R8��Kc����.�&�P-X��ռDL\�����a��./z��|F��G�_3��ǜ@7X�^�C	��#����5���m��i�a4x���&"{x�Mbf|[;Z��J�׌��g]���/-oh�ՀM�U��β>�&.օ�*�&h����A}=�Л��	`��B{i^R'�;��s�Ju�y��;�(KHN�t�i��;�m�	8��cD�輀V�bc��)�O�q��6�Dc�<�8G��F��<�a��ׯj�O�N��Uyv;�&��7���S�*�������	����C���s+E���(>p�>
�0Sj`Q��|�{�i `ӣ��h��
8�kqv��6�A���K�AQ=��<M!�,\��C� s��=G�%,?6B��)����L�?�J�ny57\rHE�8F�m�!ˍ2XVԷS�vI�{Px���+�`;�Vܵ��2f3_q�
�����C�����N'����nS$�>I��!=L�Z�}=��K����bW�~-l��,s����x^�0��a�������A��~��Z���ђۛ�k��P6�b�`����@��U6��U��ug(�i�U���#b�`+%K;X�y��6_����nś7)��T�,�JP����Z�x��=f�ȁ�VL���.��}񕜝�Ev�$g���UYu;S|p~X��� R^ִ��;\�xYB<��2n���*��8�����g�� �.����Y���8ƛ(]Zd�w�)pr5?YӢ���m��e%��0���W��ކ7�20]iT*�A=�f���U�³�T�kM�0�,�oG�_"���b��~*��kϋ�_4f�م&תo!/�ײ@�$�H�\�m�.AZ�e���<����`u�|���7����S�q�o���W�J^��o/��B�v��N=Q�D��x��:\����REb�錁�%K-�����`�*����H�#��	�j����UaF]�8��1�)��f6�|��^�/�tsrw5:��_�ۄ��_-F��r��Ʋ�Q_nV{?SX��z��Lk	�y����7E��<(��E!����C*Z� �:[Z�H��6DuP޲^!d���$�]twm�S��H�)������dc�DPd���3�3;�+S8W�����E�G�eM�z��˻���^XI񕌖m��� /�S��_x�;�s	��M���-+Ǿu��EU��m�d�j��ڽib�ϧ�������ok�����q�6o
~�I&���%�0VM����U��5�8����|&�?�μ��E�[���H͎�F�ti���P�6�NN(���jQ�6��?yC2�ԣzp��]�	�޶Y�MQ:�$��cH��@���Y��O�+k���d��><0����5i�K� =QE�sE&\��9p�!��Oy崗b �>���F����(��Q&V��{�~�
n�`ء^��~1fD�$PRvw��%y�<�"z���<���~�x�jL�#<U���. �Q��n��D�a1Zec��ƆА�� �����#�z���Z5�`ԉ��xf��4��RP��Ap	�ݠ�`�>��Eg��m��B�| �5�3�p7 l�7�1���)��z1���u"b`�3���?�?n�5��R+:�j�{����ء�'���I/)�\��{fŠq�ݓ��%:���+˪2��w��P�O�H�'݇U�z�ׇ'r�e�ra��m+	�̲	�-�j��ѐ���J�	���0x�d����;C�D,��+���8`���襧Q8�$�)q�G 1�"�=14���a��rh>��f olOk�g�J�l>����$��`�J?���{��f*^ȹ��-�%_S+�|:+c�P+^F̭��D���q
��ʥ�B~`�M�8Z^���춉�����/�:�H�,����{]��,�H�_�`hj|�u�%��G��HDswN�8B��Ә1��D���&c�<�⍲�t��ir�}N�4�	R�b��>&�q[�/�l���lÐ��[�j(�W4��PU�?�`F�_
J���D9pL� ��ju��T���x��Y��G��!AS�)��4��>B�8<e�jhn�_�r�4���S8C� @>_c���?�;/���i�JU��cb�	ꓐG3H����~�KG�p�/�]��l�0�T�j��c9�u�8zsg�:����{n=���d],>�9ί�(�+	���h�Ncp#}I��UV�y#V)�>�0
�t�ӈ�_��F^O;���X�6[6.��U�Ơ���"y#G"*�ĕ0�Dٗs�bc������B63�Ÿ+����Q&�����zcP���dF��E���/���E>  �1c���n	���A/9��d��l��{G^�c�]��.p7Yv8M��r9J=������5/<���Q�b-�M�e�+�XZ��F�:Я�k�G(q�K��0-��F�+�)��s�̤%�3��1�=���ʔ5�@x���ru����C(X ʲ\y��[e�=#`�
��sL�PqWN��˅`|�M0�W�k�ltZ���xMI<i�<i���OB���q�ő�PG��d�u�B篶���+�,�M<�-�w\�"!ZHq7K��=��*e ���!�L�/�l��@a��R�x�hrAt�?�6�T���*������t�:�T�(�
�׫�Dk��9�f�X�s�.%{Ư{�n1��M�4�t� O�*�Q#5u�/�b�����&=N�XL:5j$(.?�>c��A���8�&)�͒|dm��3 a�Sm���{�I-F����<��;�BY�nL�����\ba`~�����U���UX��)��t��@��Q:�����E�a�G�����}���LJX�6����F�����r��B���v��[��z��}�m��/�oQ�|%�}�"���6�N�_h�s�C�'��|�CI��������x����0���u�g� �Z�k|��f��;)=9#��m��h=ZXPx�>�D��.�I�9շU�J;��T.5
ߠ7ϵL���$�u�6���v�zR5c��!���%�Z�T�QaU§��ꢄ̫��9&�2ɔ*<CK��xl�N�QCrU9Da7?lhi}����dhQ,�r�y����4��,,OfT���_5t�f��5; ���4U���`�|u<�<���9�l�{�0;�/�x�S��a]g�H&ǀ�zGP����!�b����,w��1( ��C�BЊ�@@�i��l[\5����]�ꤶ�T�bbK D�'��V,7� f�p^�@"ܖk��8��=�R�7�<C��ς��N�?Dm��ǥUF�
�`�1t��L�f�o�p�:��������L6��{	Ú$9����(�����1Ý�;^F�G���&��{2��%�5�8��q�j���R�O�V�cXA�
��=QgrΌQ��"^���s���)2t��5�|
F�hJi��S��f��"2 c<y[l����-�p�W��b��h��iWdgBUA����RQһ�vo���*�\,`��UM���O����������1(ɆDRO*ꍃ����_���C#RT��q�K�t*�=np�?Fw�3�ш�����������^��B�셃����o��J�0�crC���?�w�['�<���*�k��	u�~�s�7ޣ�)e �Gc�D >Ww�����Z�W���Y�ظ��t�+��-n���Z���x������@?����T.�"��4kl
��9G|�JB`�|
��Z�O�8��w{��\�g�k��"��N�#�{G�����?ˊʶ�\�~Jad���r�Sxn_�jY���b7���k�ւ�XWf8?j�f��Hs�ǫe2���K�9����{��{����Hɯt4F�����&���0����ȅ���`���x��vͨ�h�cDco
#Ni`ob��:�1�7�.,#���8B����=U�=��A���"����Q��-�&�}]e�T�n��>��|��)��˛�(�iy��p�Ϝ�˩=l��Cc����܈%u$>a.�yV	�=�\=[")<��p}+x�C�9��I�b؄������3�ik��f}�œ�K���^Ec����" �[CD��N���И�b	����l��Y��Ƣ)ˌ<�6���;���7H=����p�Q\�:���-H�j����h�$e���=���,�]?����bj�▢�q@�.��$���fy��AŲ��r���n��A����S�'	�n��k�����xz|28k� �x�4m��D-~�I/�*K��\nζ�7��[�rr����b&篊�|gY���@i�m$%+;E�Y�Ĳ/ծ�P���mg��<�e�^�_$sA����C��f��,��L��w�����T̤+q$�a���\�f#4�s��<8��tG\���+��E�Jq~���-a��ո��rFj��n(�����k��J0�ћ:<��Ӵc@�4ҺK�WN�_1\����Cg�u���C!dYP���p$��8su}��X�ެG~G������^���f��&�ɰ
e�*E��Rg�<�!���VJ�˴x�02�0@]�l{h���E{���S�;Cy�O�J�� �staz����yZ��O9G0��>)g�N2@�$B�J�{
���,Yo�'V��x� �j��A��Z��ɤ>�,��v�O�����\Ju�һ��H4A��8/MwX�=�
���Z�1�9/��Z`m�����mْ��daV�����qaR�xnIڇ�hg]v+�W([�2qئ�mK�P������N��l�\�Y=��J)^�q�Cf>~��q���0�g>����+��-56�u���Fll��o�@�WQY(�Ƭ��x�3V�0:0���zB�^���7�U�)mh� ����ZY
����`�t�Fe�I�3���BSI�:AY?��NE<)�N'<Q�['.�A[�����Q!��V.l��L����Tљϒ��Ò��x�����h�DX5@A]֠h����䐼2���7�ϑiᩒ@����!ϲ����˚��T�8Z�@I��mٟ��`n�Q���P�b6��e�X�Ѝ�RB�d��`�s�J!� ��"�۲��Qu-��S���P ���o���d~���Ƌ��Ş�7݈y鰗x2���|�d��~���L{u�FD��1NM$��2�`">���\n5Q �T�ƁGhR���Gz�6~'6:�6�EL��hl#׸4͖��h@��͘��F�J�v�Ao�i���o�9��Cd��2E8�7�طi���	�)N~Y�LZ�U�R�(*HR�Q-�M/�@�a6[�X�(P.�6��߄a��#	|7�Gf�������pF̮��2�H�Z0#����a�tM!W'�iz���/�����e����k��L~h�&�����y`�U�σ���d�y���P2|X�Ul��S_�˩��{���1�r�ԁhl���xTDA�����5��G
X�Y`3$� j�9���!�Ci�e�ھ�?pŔy:7W��=(r�jm��ڬv��/�/��FϏ)e����2�_NnK��X�����݋yR�r�0�v�S;�Ҿ���rd�N�[��T��,hnh�-�$͇����`��&{��,�"EuNj�c]�Nި�@R�AT�B�_X0W�Xf�L�;�8����-�B��X}W�j��[ N�ΩPc'�O(��z�ޮ<dn�@�ێ��"W�_���O��?o�J�1��JB,ZD�5���i�������^�IP("�1r��&�3+��n�.��x}�f���q����Fh���v%��FF��eR=�1{��K�/+��gQ#��w�K���f�+���	�2}J5�"G����3�Or�f��w�
�Xo����k<А� ��AP�m�z�@����P�+Ӽ�01@'���b]�؄T�Y�칀$��N��,:T��5h�C=g�&���ƺx�ӖQ��߱wRcW�����N���@��)YEC�u��"�c@�u����!�n6*=u�x�#�YbU����s�˗z]hg7�;�%1y4S���0mj���+���2i?Ŕ&)/b�0�%_A��)C�i��;��b4l	TCw��ys,��IB�*�Ф�d�R���Kq�Ze-�:쾊��|Iqg}�)����4Q�y,�8�;t��SҨ���%O���υ��m]#�|����6�	N7�ϣH�ն�,#a����6n\�\�$�h���Z�KKN���b�NT򓹨D��a$�{���V$��솸��5�/�6$0��X{�.�
�f���_������Bh1q�&�Oޢ�|�g�m�~�%�x��o�d��'(B���3�$����F���Z�Fdꊋ��v�+���{*����?<r���=^F�T�ie'���p�*@eê�w�.o�x����գS|��0b?�2��{pJz�ց�����aH�*^�2R�佴�A]�����7IJ%j��7��d����عZ��
�]��+	��κLc�m_u�"���M1g�	�>Q���Y��ݙc�s=�7So��z����q^撧�X�E��,x6�y)�׋�=V|��Gb��O��Pg�v�M���yeZ��7�ܺ'��<��\35�CD��[�ckfr����%�-�ɏ<k�>𕄄Vw]M���f�=x�l�Հ�	��J8����l�D�ߚ�^����M ݎ��@�be��1�zh��I����"%OjGd�]Rӄ(6g���i��L�O�淲o��S�0I��¸������0H=iLmeF�m�1T���t���'U�#�E9�P�ϱ�����Ad�F�O�.�*�8{��`q��W-:�lH�ō
������tMF��/��|�քk��n�b�l�C2�- �^
4�����QCކ�cw����g��탫�v=�f�����CZ6\��0<
���M��W��.�-{*��d�v��u��;\�o��*r*ʌ��a��?o��ޠE �
b�G�C�S~P�CI`�/��$:� F.�.[�W2Nu��2���΄	�����`�+�L��`_D!�CA�)�4��"�����T{wS��98q�.aJl0�6�hί=G��T�Q�xst���őH�Z+ã�F)���5y��e)�z�+��^�A3��q�!K��d(�R������.�K<u^�[�Wn�p���W&���i�ܮQ� ��Z5�vN�)���U������n��s�'×�묲x@m�L閰�C���E��d�5y�O�۩Q\}z�]i�m�1$��2����^��,�'������'��f'�H���jx���[���J�\�հh	-���k���q �ly��dP�ܠ������osZ8�"�E*|~�7Y���x�n|+���ݦ�kx��V�V9���v�u�|���-�\��	ٷ]������q���	_a�!MAm�v.:��yM%�m�t����g A��{�sg��C���<eT�� AD�|�	��z�:1u������9-
��.K��UFc�J��y��r�(^�/�cs��1?&�����O?��Q�]�(�h��Jr���O����-63k~�ܔz��P�7�ciTnB�o$�6`A�U���� ߯l�!͇;a��M��iUm��&+ԧl� ��׺�&�?s��<­��:�v9���j��[5�	���7�[:C�_���2���lܟ�I����<:�+?f�5e�?�'}�<��PV�3��M��xM'�D^��c�W��� ��է	?�Zٽ�MU	���PH�4duVLq�kc�;��y�c���˚��1��\���9�����lo��V״�h,)����X?ǹf_3�!�ם��<���	en.��(
F���� �|0�����5bZ�V�Qi@�~!
����I�A�J��ٲ���KA�H��V�##<!�@��ŕ:��狉VRQ8�>t�+齳�@<~�E �%C[�\3,MB��'2_�xbRL.�$X���#^#D�*���r��I��2�/}���JF �/�4�'�`$��q��u�!AL�VH�X��a���1��	@����Q�-��%��Ĥ�!{�3'�7?��kDH1T,S�<����jqL��뤪	W��]�m	��*0{��	�����VA�9#R0�t@
���v��mQ�2�4�o6���K����k����Ø[3g?3ƅ'�֡eVg8��C���SQ�G����� T�V�h�)>5��6����a���{RdU1B�Σ��~s�n{ȱ�1��J��^�;Mh3{,Ωj�;�;�֑'�K"��J����ZP���%���cX������<F�L�9A4-ǡ���X��ԃ���C�!#�H���d�u�!�<�`��O���ǋ�}��Ž�����]�c�$�DgN�N�x���xN�&�$3.n���������Kd�����^
|�Ah����L��Q�o�w�ho|��xsǚ%ү�{�O���9s.�Ġ�1A@t������
��4�=�	Z���,}{�Q��_��Z�dO�:�@�c�qKK̴j�R/�b��$;Ji�ڞ&������~�ƄH�䫛�����u�Xy�%DL��
�_����2R�$��݄o�M��-if�z��s�4���|�rK��k
�a���^l?�.�8!�X�S��:����k�L�;Υ�T����͓k���v��F��I�n��0��m���տ'��[f;���vT�MT�����!(7�<oB[>�����&V��cA&�ؖ�{���v�c*���k���r�{@�'^]Kk�`xǕeV�w���UN\��z���.�j�'�wO+t�����z�^k\�F��|�\��/�|�5C�j�q��/���s�S6!`�{�s	�o�ZV��86-3xߑ�u���(�~"�7_hѕ��K?n��]�1!��6G��TI2?! ��~ �cD����Xus
����StX<�?��4s�@S?:H0ZE�4'�\.�ǜ��� ~�E5���2'%g�8gG�����6.UU�wxLx��ф.��Ypg�0���۠�BJ4�\�&�3�m�ls� ��0�,��7��I�u��H�C�zO"�w�#�f�dh�خ\&���m�j�H��V�*� &����7��Ї/�e+')�e���񥵶T�OX���<�������t�b"8�o�k����,c��.�
=�YM��'y����%f�?R�������\�@q����UP�Y�e���b��rB�hИ^\�bE8�g�*h��ȜX�0�LI�i�\�TC��6(E�]Iz����M�k|��|�{>�㵳�ڋ�zb*UHg_E�A���1���vA����2��{n4���8S�'�����u�큾�1��,�̜̓o��b�����J�jR�\��B������M��5���Tc�Z]�^�[yLp�!��Ր�8!}/��y�Y��D�7
b��m��Ra5���8X�r@�S2��zRj�)����(�h��$1�FF(k>��s�u����^��geڛ�+���� SM$������b������$t$����B!��lU������gGL腶��/R��#���es-�}E�W	��)��ѓ�ܤ�l�#������c� >d�R�����������H����%�	�'�[\�XK;:08�@��th�O�{SY�z�}avV�N��*{=w��g'a<�:(&�e�K����H�]��x�E^��I
�Z��<��?��X+p,?�>�P�*@�`��r�;|`�G�!?`۵T�M��B��6��Sh�?׶�Z	f���K9�9��O�0ö�����_��Y~��@Ѷ�����O���m/���odm]?0iL��_1J���$�<B���	R{y{F3�w2�Fu^����:@�j/Z�T�(S��#������~{�超ׂ�Mra�ļt�5���lg���8��"@�2�gF~���L���4/�Y�8U��~�v%]�k� �k�7��>�8e���=��Г�mm'���v%�����bq��{�R�%v��y!�� �cA�����A&�����X��$	���7{�
n"߻���7(aU׾��jU��'�R��u4�C[��\B��r�g\������KMn
�Q��P�����Z��l�>ڪ�߮޿� f��,1�P�<�}U�p	��HC~St���ک��a�q�2!`��+A���@1�jn��u]|d��w�U��w�K�>�1�7`��	�U@����I�T%t������\1 d���<l��H�PbŇ+�
�%Q�d'$4`� 0�r��������a�R`�i�weop�cqjo���Z�f�JP�ל����'�f�m#������w���PYi��g̾>`&�[���m��(��p�FUw�^��v�s
d�����qU�U e�����&�~��t�2QY��jIa�x�\P�C�PS�a7�R��5u_�8�ܯ��A�e��CR�-�(=��@մ�J%�j|��kՃ�ѕ�'��4E�hS���SQ�V"�g�y�����Y9z��*u�\��O�E30"E����oD?����l�o\�Ů,4�_�ӱJ��bb35�żP����'P<��]�CsH*�R'N��ON�{w��4x|L+8���,f��Y�z2p��sNQͪ���[b�
�^��6fV9;�����x�Q�ď ����}��'刧��̌R�&����ޥ95Nf�ї\�p�9�@\uR�Z��]���ܽ$��Z�!���ҏ'I�����)/�ah�r���Z]�[I`���-J��XN������S ;�(��O�+�mI(�on0e�l�F[�+Z��;B��Vf �����~N��ж��Z�#����>#�L _�����k!vӜ1G�ZӚ�������T���6Z�4���jQϻ�y= ��E2rp/�fj��l���{���F��u2O:��f�R�c5�~i6$��l�`���.��t����(����� 5V��S4\ƅ}G�"�7ku���-]�V���qq)>9���F��䆣M�����NTɗ�s`�ûV�[�Qi�8��%��3�×�Z���5�/I��Yc��� �g
k�X�S�u��Pjo�P�����f�TfL�<{��a����M
�b�������'�`H�8R{�t?�ܶ0zYaQ�ф]�j+{���~ܚ�&��{;�P:�+�	�,���/JJ�A��Z �9��&h�z���Tv�K=��ҙ�`}V�0	���	HP���iͩc����i�F�����:JJf�#"�9�VQ
�U<�2&�}���-�*k0-G'�X�
b��oZ��l�땻�$�8ȵ`���'�a�*,8�f� �g�e�f~�ː熖��̜������{HwO�(�����γÆ�v��t�����y��7�J�b!��1N�P��c��}���R�7����@�d�P�;��{�,�w`d���b���$M�!�F���25���Iv�]ɹ��,*4��s��IG`��ջI�N��K��WHֺ݅�	�V
���R,n�3^�<��mX���$Ak�NH�{ )��,��ȤȒ E��id�,����X�ڞ���jI��o�å�ͭi��zt��m������͹=v��D�֫0������7�G��,(��`"���L�2�L��Y:�RG'�<���NPmInܬ��]j��@0i�eA�\�������o��ٙ)VnX[�a�������B]<-��m.Ǽ�~���槁�+������������t��ϛ4��':S xK��US�1�d|7���|:�,W�_�3����@�o�-���꒩@����a���[a�{.c����'�V, wHa���\��M�F%�>�j>�L�~�4���@����t<2��jz(�ߌn���j�'��3�3�?�����D�������cM��H����f�œɳA5s(��a�͓Ii%�l�f[n)=��f?�H%��R�aK������{�����[�T�=,0�kJ��<V�Yj��#�|����H�` ��l������磘���n`&����RK���J}?�h�"��Q�"ka���1y��Z0�nӜ@;l%�^�F��Q�CΗ�_y�3M�k)�
�>B.i!t�,��a-Ɣ��v��ŏ��2�g�"�d���q�['�H����a�j(�t�N5��#��_��N(=w����(��̀3mw~ �ʾ��@� %�378HJ�D���Z��wW�3bT=�R>�s�%�o,�V7��f'3OG�V��F�@ŕ.������������P0h/wd��P{搊7�Vg��f�c/Cg�C��1>��+*�"��q�K>�dH`��/��8����Z)�""�f'�#i ��EXiv��y^}����]�"�Լ2������ �aR��[��`L�j���(�����m�#a�7�,K$&�f�w���T;NhOEG�(sTV�X� oʒ�[2�����<�E_A+�Z3���Y)��/�M��8c<�w� nmPX�I��c�I�hz^�@�� �n|)���Z�7:�SPd\JKv:��bH�u>C���?%A*)2�y��������K����&"��Q�9)����[qG��.���\e��9�HB T��Q�O&Q8h�(x3�Y#��_Y�FM2X2���e��@�S�Ҿ9 {pi��9��g��. Ok7�Z���m���W��Ŝ�i�x� ��j�$��j0���#���?�.�2*{T���O�<��y� �tR���!}�!9�(�>�����#o7�-�Lҭ�~��B1#��v�<x����*T@�����n�ղQ��Z����o9��Q/ x@\��R�=����2���ޣt��ߌ�`�AFퟪ5�����S�n��%�nh$�76�{�vf���k��7��{�GMmP��b��w�q�,U��WKdZ�z�e~Oˬ��^1V��S4�d�-.��ۘ�U��Do���k>oXޖh�Cf��t�z�j9,7��(s?Kj�l�Zڴ6u�O%�JP�Dɟ�ng�(�S�O50��Gi@xc�>�|T)��߰48��V�+�	F�x��N�bxd�Z��.\#!`Ѻql�ۭ��v�<�~P��wa��Y�A�E�v��2B0�[w�|[l6�֡�z�]}�rf�˭?�B���T�ZJVP�Qf�f�Q�q�fM0�:å��m��(,�XZA@�o{v
f�<�B�|����Y�0p�ԫ���`�P+�p�D��aܘ����+�7�~l*���q!MV�A�fB�t����+!��f�����nf2����պ����k�C�5�J���p6c����;b�����U	[$���y�	���N�EO88���Br�ڵ	�C@iԵg���b��G*�a����|����5�+�+lC��bO�E� [W���eL���8��4�ܘ�b\���5�����1�,�I�s]���+�m��5/":��Ћ ��X_��R�>=S��'�IiɔZ��Wr-�.���W���iZG�'֓�nr�o ��ʲ|��A$bqb-�q>�s�V8����P��I�=wQ�e�*C��PY�>E��F�5�\~�Z��idŚ���2{L����c`\D����&������L�^����� 9�x���{�S��#�ꃸɃa�Hw|�DE�s����枑P� B���A���G���`�g���s�]��4��n�������J����e#��E5�~T��Ď[6�Z%Yk\^4��{�,N��ȭ��Z��NV�[hU6�-[���r�h�r�Z|\��#��&\�q��=;rn`�W������%�zx��~@�,����[����xg@9z��	�M���@�>6�b�:0��S`T�x�����{��$������E�7�I���3şcb�� ��7t�61^3K��]iC�.�ɜT��R�ĀZ������(h=K���{1���Y�qT�Y�	m��Sp�9ݻ�?�O�q;"ޝ�"1�ƫҭg����3}k���u&��p����UFP���ֱ�7���P�h�T[�t��w�X�!Đ�֎z�#�r|-��)Es4���?�uJ�6��6 �.ɱ�A�v�U�i�[��xm�m"?s��/��ʿ}�>��*�
�'����x��\`�Wg�6�9iQ����u��g|��<����	����i�,���5!�I�(#�%&9M��|EЃ`i���+X�o�D��Z+*ۻ�{�[R7f	���P-�}-�S2���@�d�#.(�(3>l+�h� {�m��a��"'(�o�㲨���~UP���!�3�9DoP��+������ؒ�u+�o�(t`�\�������cC֊:u�Ԗ��v�(K��rZ�y��#���Y���M=M5���i\��� '����x/��5�	�� �n�%b�x��h�
�r��a��T�w��[��k���.p�b��gD	�a��"5�?SZ�ԙN�2o�p)B뒟�8��H��y�m�]B�͊T狄���qDΚ��⊈��ƪ�veF�e��8Z'O�x��2QUX �˳Ӗ���<q=0�<�B��&��!9���*գ7��%?�lG0��X�܂u���m+/����ﲻ��F��!�k��8aO��{�8���zX�s�F@�dv�4Ɉ���Q\�6�x|Jn�L\O�V�t��q'��<�\�g��M���s8���k+��cs�+�[�Xd�������z��c���YK��	Z�Z�2��z]�Ӡ��_c���O�,(G�?�Ab�__�<U���7��r���-��X�
�e�Å��:�~`����,����h6����^y��SIW:$ybqG�o�?jb8;8�omE>�R�h
H����{�Zl�����Ox��N{b3�-�{�s^�>q����߮�௓rP�y%��oCս�R.�FP����_k0�ǎ�J,;�{��y\Q�������kLȏ�ý{���D	u�ZY���TXn��%E� �:�������@s�@�h��g��*}ٍ]��e+�����r$�{�0���O>�)�_z �h�-��ȯ�치������9E�����v.bO�],N�ȁ����0=�g��O��B��#- p,ۇX�o��&��������`�
���A��*�+}�SA\5�����]����":�0��m+8Q�֧"�3nN�Z	b*1XCR����sG+ajˀ���vt���+ֽq2��ݳ6?�a.�B�\@R�u���@&U���2$MT4c?�2�8e���k��y��DKzpt���g��'=�C�+`15�� f��`%���co*j
*P]GP�}��m���wrբ��ӵ�����f����"��E��]�>ű�ɩB���A fv�c4r���@Ei7��~OK!W'.j5�!�r.����rҊ����*��#�(q`�D�f��@vO� ~>|-�Ӕ㻽T:�g����R2�?.�H���)�,s/�t�\,�۞�z��x]?n#��� w~��i��x�#3#�в2P��Zy�QxJ�QJ ��3���t��h��S�v��y�7X>w�5�i�pB�S�_v�rVg�L�صH6���3����;E:�� �1��s��rŒe��_@W$H�B,j���6�=��[���)�Ѭ��(1�l�W�	�Z����_'9�*�gy	@�W����mi���G�	_�����%K�U_���J}��Z��K��Fh.�_��I�"3y�i�d��2O 7�h�2�>�p�8�%Րm�u�$�>=��G�	ΤDҀD��$�R�����^���t����M~h�eŸ�������ɘ�$��{@�Ν���>�0aXXĉ�0/�,�� =nO1�9����2Y�aqp;��[4M�?���ZC	�do4�I6d�	�I�P�&��.9���Jr�Lr6��>���hj���Rq�q�ύi$h�i�����f�t[0��~�H�Xd�ڠ�(�h����^����N����,:��ByK�Hzٍ)��м�������4�������w��sj ��!�̋@y�$��wL��$vE͋�7�7�sg(�Kh3��@�I�c���P_�~�o�o��E)Qd쟕�)��oI��G�\�ы��J[3<�]�|{�W��i	U�H~i�1)�č�5\(�+�8ڵ*En=re���G�~���h��]'M����:a�J+vv�G;�������P�ղʊ�|&��*�9�/p~	�c�j��,����A��	&u-�����������
���ȇ�q�H��v$ZB�Zy�_U��|��	$K9*!�����m�U�x��Q����M1�ȁ���tY/r
팒s�{������Cu�h�sa���� a�ܜ�>��YR�l�άXh���5ѩ���O&��Ƅw�(ݻ�u\��'�����!D���������$���?�1�QT!B}�c�IPu&�E'Y���[�sk�W<�����/��qCqg�^�F���N9�&�׮$�Wx���Q*M����B
��X/�{�&�]*_���8V	��T<�t6�Ɣf�x��p��<�#ՄU9-�E"��^�6QLH'���2�1{��c���nC���Hn�dI����Dx6(��3��q_����c��J舸�, {T�ٍ���|�$�*U�����x�Bd?D�gރ���ZƗ_����s7S�d|Ť}
�o��W	YT?㇅5O�Li����[ \Z<o���sz�,���RUsҙ�tRoU�􈩰��ݧ�	'�.!��Y�w>4�QӍP96`������>�+Ќ�i�M�6ķs����2�bA����0�Ц{�ò�W��A�+H��!��P>x�u����.��wЈP���aivV�5��C;ŋ��׫�~|�}�A*-�;
'�A���C	�J��Wt6�e@ݢܖ7��Z�ΙNG�Ũv�-�q8�����6e�5{��ђ:i�݃8<^���`�h��-��St����V���ʋyo�b��_�����~�jҍס�UM
U�V�'�E$àk���\������-�VfkP��y�x��Q�2���r����Q�J�Q	�|ئ���rv��j�������Q���j���|��x{a�����]��	�.u�s��<O�sr{�eE��+$r�Tw��~3���k�
�~�"�"��A�ﱠ���K�yYͅZ�6�{d>H�Xڞ�������P�{c=�,e����9?x�q$�M
$O�B�bf�I9�=�����]�=��(ǻ���ͅ�'9����Vz[���G�o`�-�v���H���+���^Ox���-O��B2�c�B8	��k��;&X�l�|�
���q���F�? (>J���?a�B.���뼫��4���)�����:׾ϡ3�MPLVG���o�q���0җ�tq�4FN��^�Ɩv�������%�n��� ��=��?~xBT���s��9 �l�upSBԘR"��SB.~�5	�$��pC���3�̛����.�Iz��gĊ���i�Rbca��Y�F���>ߞ�FA�����> ���E�m�T7����-���`6!jِ��7�4���<^ڥ#� ��r�{^�m";3�E�sfX��V>������%�8i�������<�p�(�0�z'����di8��m"���#HP�b�_�aI��a3Ψ�t2;�җ��<��E�81uu�������G�@��d<w���}�͚������S>xO�=��;�I�7�>l��Pp���Sb���ڈ m�.I������H�E���Q���sv��YA_ ����T�S[�gؼ����~s=�V���K�[��'�s�WزW�n;��=�|��zz�r�K��C��s,8E�@��5��W���	.i�Q������W�8�<�fj��=��AqI9���i�C�nR3�jc�eX�0K	\­�m�JxHPW�]��B�$�Rq�ߝ��[�L�zBM�����,��>��L�I4������ʰ��T�$���K��RU�<E=�������.O�K���C�|�`�i'+�q���?$���-�R�>�ǶH�&�M�6���<4�lZ5ޠ�%�����H���6� .���Rv�Ka���a�Y�����\���%ubX�AE�k��k흓ۮL�S-��f��yf0�bb}K����6��#i��b�~����T���EUɋ�x<j�/VC�Z�+�Iz/�8Ƭ��m��N��`$�����|$J���푰q��
�Ѳ�S�*�ͶY�a�.�Qz���P"˅����E����1��j9l�%��U����p���G_���1h����:�_��&�H���N���`�
��KP�?�l���!+���M ;��W�d�o5�������qo��$7�n~o�������"�ܟJ�*��K��Gi�׈�j�xcJݏM!8����ы���4����U�d��=�J�Zݟ�_��ų�?�I/)��=��z�<)#bBE��q|4��C�e�X%���!J�`�y_�̶�~�)�)�5{�B�~ט�Q6�f���X|{�����1k����.����x@�@n���ͱ�3����	Hr?�ϺLZ_�l:C�J�i��j��	�@{b���f� �њ�߾��:tc��w�=Y��1�&.�o����P�&��[�(�����翐��(�:�4BP�@|%��*��x��U���ZԊ�E��pgK��B�0��0WI��vX�y�򋓐l����*t�JN)X�]tbk
hwO�IT������{�ŜNn����Ni�h	�/�J�j �A�wlߐe3TWx� %�T����_B�O���Mއ�U�w�Xٝo�W���d�Q�,���A��d{�=c�G��2��Q<�G��������P�|�P��ˆ�ד4�BR�a�ߞ�˸�cC�{yҠ�_0Y9L�MChF!��%� ]4�i� >n�rꤢ+ĸ�Q?uҽ^_[F`.A;|<\���b(� T�	����v`D&�PL�>G��sT�̠+"����x�� �<h80����7`ʙlh��F7*��)�\p�M@?W���=�@4j�\�D�z"[�iKC|T�=�Γ_8��;��^0ރ;�_3v��k�{J.�o� �h"�� >�S5�Fb!A��$c��o��<���;����g�����K��0�hD�j ��T��*��~I^�e%��1��@, �s��Fӥ��}��eA^#=}`-� �!j���\�S�5j���?��g5k%��#q�pVU���?7V��|�KȟO��9oM�Q�i��	��J�l����uR��^N]��0��N�V?"���)��MΌ×!_r�	�I���u���5���u>O�R��(v6���[@bW܊�f�Pkp�*ɩKτ{ɩ����X+�@U��w���w9�5��A�mH���&Lq>��*Qo�`P��r���ψF�V��;q_��_԰p�������=�����f 51& �n�Y�Cңm菁���D�t��M*����.Ɉ,�T��.aSϦ��1�B%o����:�N��e}�G��Q㞊���qtIB�pgIK�
�}�ȢC����'z�;�SzheX9?��+�@R��:��ev՟c�g&�Ky��s9ډ2�¥*=['��M��O�#K���I&w��V�9m�y
����*r����Z!����Й(�T�α���Ϗ7�3g��D>|�x1*B�?{6M[ ����l��3]5E�~];�zN_�Tύ}�_^?pA^�8���w��L ;h���C�v�⚥{@
�rX4�0�J��M��V��kc��"p-�L�v���r���2^��w���朡�E��Fn���xL�U(�"�H�|e��57tQ�B7��[ՁJPLԄ�ٰM'� ����0��-K�,R^��Y��ݡ�z�/�(��'�N�+����ĵ���L)'�$�\��
s�2;�L:M<�pra��%������X�kg�}B����o )�M�yg6nOA�G�#����{fnIs�i�8�l��`8t�Zn�3�瑝Tcv#�|���;�p���{�� %qy����@6{�9��ڰ��4p��R��O�a�6m�L�)\8����rr�"!Ʃ:&�9��`<�|X�긳�uz�c\Rle��xd��<ѿ~�+�7;��q5��e���VN�=��u�!�A���"aR��/��Tlߙ�d� $�`�]�cW�6l�� ���6A�A*�:�U|��x�Y��=4�Z�z��3���L{���������'Vg��b�0PH�@0�[��v}��ݽh�Jb�V�-�Ң�I%�?N��ċ�����wtaSvw�M��Lfo�F�!Ga$��u��u��(l�5���f1�.(ba��7�������;L��&��z��Y�n��Ѹb.-��:+�*�\�C��t��Y�8_�h�dd??B�f��a�a�뿽A�]X�-��T"0~��o�Mvg*��v
Ƃ�f<���Ҙ���rYߪ.�Z��}�yy�I�~J��Us{Z�!	����aQtǷ_18�����8����QkRߜoX��Vy����O}#���)��$<��A���.�.�Kw@��:�hw������;�s�;  �zG�v�@^���_��Cmm�M��,�C�̲8�8m�EI�}����j����a��ύ��0��X�M�R,���O 0�E�x�b�&VjG���u"��"�n�N�+32-�o��s[3b�h;-S3N��0�L��ݙt��p����hT�3J���R����v�&��I�c��Pb�WbV�C����ۊE�J=����6�@��&A{%���E�����ek���D����N��x�Of�y[i�ܪC
�����gڗ0�rv�d�������/&���.�%C��m�=�E����c��aאо)(��f�;�u=Z~��{	KfH���i��G�Ƨ]/�䯺���w�����|?�0�p��0sU{'�8�+g�8��*a'� ���	��O�Ɍ�;.�:��h���.�q�c�9�?���F��d=Z���\�߄���(�u8�PTqf��Ӱ(� DF�tz ����*cU����i�c���{� �*�*��. ����uӾ��\1}�|��d�3�^Ԍ&���Ř聆I{j�������E�L-#����7�u4+¯�^�Y�0�]5������R�s�U9�z�?Ԡ#}��ͣ�2+ḍ|�sa2��;�%
|����l���¸כ����;g8�xnA#�דd���KV%������ڷs5
\j�s��^񄻴�>�Uߧ�s�����o����4J�B

G�
�z�R�r����r<V���"[{�������M������z���6;5�%5 � �rҒm�ߟ>�W���{,e�qAmR�衊b���������@�m��Ԛ���d�}�Z��6�����:����2k.h�;����t�W5+�ĭ3?�SrǱ�?��rN�0IV0��q��kPx���{4��YZ ��LN�hS�h�yw��6H���*��I���2K\����Zz^���|����}RDƃE^tVO wx��~&�Yƞ{d�x'K��_�<���MB���}F~g���rN�V8�qj�^�&8K�pxH���#��rG�[lq�_��J>��p pe�ˌy�b&�)� ��G;CJ_�H��_�U���%�>'�Y�ԛ�A��Ɣ�qG���aní%-N�m�5�OJg�i��
�z��U�S��e��I�?f)n9@���#o�ǒ�9t�5�q[�[��=h{ۯ���9d���"��܄d\&]J�̭�o���e��Z�Ad�.vB𻒐آsj��ԍl�LY~���pn�E��D�YA<�؏�jPl�zq�0���8x�������HgQj�NM�DQ>fP��'R�>/%l��hF��
��)(��h�ON�w�۠����Zj����sI΍(�_�<ɗ�э\pE�|�Z�����Eh:��،�у:�n��=p[��Ϡݩ�4��oY��b��ļ�qK�І�w�2��$�+�)"����L�܊�M��.w�Q�Mhk��Fm�>��+� ���$����R�B}�>�:=�I7�8�d}h��|�m�ƀE\p��Pfb�ͥ�1$O=�yKqs4:��	�}^.�G��E���(�7�.�p�Vz�|���Y�Ŧ�@�;�����<�k$���ס�\���m�ʡ|��:�G	��p:|��~�q��n�V�N�;�V�Z��:?�&�SJ�*�cR~M����8��"�J�*��)�Z2�ZZ�<�|�s�Sn.\�N��-
��z��s�
:��N(�̝lFu�0���x�%�B��|�`>q��Ooǋ�p��+Ģ.�[X;����_�T"�2�Vd{¥<���2!�y�]�Yd��_U�~v{��J��*�|�*�r�O��� �GޱYPy�#��D���Ό�_񽯢��c~^8���g��	��x�<�94>�FAi=J�`�u�8�s/�⛠ US�>��|�qV�Л�0��~y3��B$4#iK�HNX�E�&%!n�c��̀��剳;�Қ�z��г��g&���"�j��3H!ާ<���a,��v�4�_�c� ~i<�*~��$��v�Y\�}��s�H:m�]�M;b��N��X}�7���T��O��1F���A z�3Y��px؞��mf��G��
�S�p�#�ܧ(��u^��ЀqAw���2+�x�*մjMC�ꕊj��O�)��Ȝ!0����xcK�=��z2�:��P�<�����?�K)60c�o��Om��&7�C�BO�e�F�W���BA���ܔ��(�'�6P����Oڣy���G��"9p�h�}�^�IUc�w�xJXl��ENz�����qC8"ǎ�"�2���5}��R(�+�v���@�g��\����3{�E������#;M����s0cp�
z8��K�\�f�����P� ����W�\׏`�q�W��w<��L�B�*�j��2�֠���ĭ9f1%�)��D�dzͰ݇ڼ�kV	�+$1��4��l�К��y������i)�Z�ʔ�J�+�OS��x3Ã�B8��:�Zw���
�(�#4��E�Ǐ	�V�F��������#箯sWk�������к�+�O�-�������O��wu�N$W�E/")]hpSIΏܽ���)\�4���At�y��Z��b�~h3�������jt�MȰ��p'��e<��nQ?��x.ϔz��E���=e�
�0��t���#+N\�*�߻�H�`l4�V,z`��q��ݥ�E.��w��Q����o禝;�#���\��.���v��,�.��c�p��h��~,&���_��E�^A߉�m��N6ؤ�7�S+�p�)cƭd����%+L��^�d�I�L?�W�z���Yw�9Z|��X�� ;W:�X��<�٦Pha���X)>�5Z���)�+�h�؝�.	5�YRᎋ.��"%8l_�����{���f=��z��f���Ju���Z�l��+ve GL{������x<�Wo��[��_�=�L�i���rQ�J����And8{��;b����+k�7�m�C�R�*]�������̫EiR��=���u�ʇ�꺙۪&%����X���W��)����<�2�7)�����x��U���o
8�&F�����{�P:���-i_�k��~��lK�j�Q;4�����i��פ��������gr��[�E�W��Χ�<x�-S�
7�noRJ����`�voVZ�'�S�T'���p}����Vo�qʗ����lG�?CDYR�Q�&b���|I6�x�h�Q�#�K0I*���-~��D���0��1hTp	Z�맯)TG�"��b�G��%��1J/M�k�3}�^�f�=�>�ѭY�!P��|�$؆��e~�;���V�O��dR��R��GW߇:J�w?u�����#`*��ӕ�����=�)Xׁ�_5��Wb:�
eb�D�8{Btʼ䟦1(y<J]�W�H"sW�~��Z�=�����`by�?f��$tӿ �"�@bt��]-��|s�2$�sdnb�Rfh��f�:�{��3uJI� 7q[3�{�dQy�Y!HJ �}��,�n3��nQ!r�_��S�C���
 U��W��*k���/��(Ԣ�ku�8��G��fx����3)yGl��H��݋*Eqi ��wQˎY����榽�h�t������l/�XU��@
+���7�=e��?Z/c끲�<�*��:ڏk�������om3�C�H�Ӎ#��Ϟ0�U:�a6���Ϯ�¦�@a���m��Nԓ֧�s/҆���=�[ۼz�we�J$�҄�C�u��l�0��]W�9�ˌG-�����>J�@�G�+
�/��eF�%���>3���i7Z��g��⡓��O�IE�1h����]���f���Մ0�+&� �9��"7��_z]-�x�.�	i|�6���ӷ���
t5+�Q�B�H�%���{~�&�nK�����Q��r��b�ɿ'� *D����NA��ĳ4��yl��<��:4���Np��f5�	X���	��8��r���w�Q�K���Q�BAz(�,�3P�.�0����$�W(oC8E��{X�<A��.�ڵ��v׬rR;S����/&8'˭~��|G����h{�Ff�I�k��7r�i���ĒEA�2���2�W�eN~�S3���M4���,Љ����Wj��b"�-��k�*��F>�{�g�~�1l�D���aŰ�*H��g
��ݍB|X�C�U���-��q(Ai�I�f��LR�������]����>D��x~<�HBrR�'�Xi2Sx��7S��KW��l�P�/C��v�8+�5�X-uڲm�UUNE}{�ö���5u�ՠ	�����NW+�9^A�YQ? 5�W�i�E�+����pd�<@-[�^ٍ\ц07� �4����{qP� s�S��$ߦ�;���1:I��9n1�u�1	÷���K�L���$���#���*�*���l�u(�	�в=�Ou`�I��#��eW̀,��uJ
�� ��[����m�1(0v��~|�|�Tp88^p��բ�
��f̃t�,#_A�k���H��ǲf'}Gj��V�.����׶Z鸌�p�[�7~VU����ړx����h�n4kY�������<lM��0g.�E�E��Cc��ɬ̾.oa��Y �Mta�N���_ry�]]�2^�a�_��^��9�ɻ�)��@>1�Vb^?�r�6�>}��æ���-��dxxh�A~VM�X�����*��(3��T�)g��4����x��i	�}�b��5�g��ƣ�EJ�|b@���1�ǒ�,�M-���N��9�ƫ�d������(u6l�K�ӆR7��MjƷ���
�	ͳ�\��w.Ƙ�45�N���Z�����2	EiE��q*��PC���C3:@�Z��a�[�ׂ����Y�LVf������%nZFХ���
&'B���Ƿ�q��l-+�qШ�>�Ɋ0��������G�ؖs�w���/$7s�	�im0a�w��[��������GEc�a�'~�쥡yTZHIoǽ�2�q���	i!���j�1R����P����=����@�訙ŝ����I�.I�݌z%�\={��'JJ�.���6�x��y0��W̛�j	�H.v܊W�Y���-���O�/�8{�r*,�����e�u�ZEK��ֱ�A�I�VN��#��Fi�Ʈ[�������٫�z�u�����΅�yϰ�3L���n�Q-ѹ��0�d���j�$�D�wD�ˬ�7O0Z��
�+�z#fh����ha����+������ӕ�gﾧN�9kn�����y�m^UIp��s�2C<*c��A'd�S�"aB��S��j�ٕ2<Gb��N��k�x��'2������*�vdS�Ь��#6̯��\��)�6$�N���%�j�CDq�m2�[j�����i�0��Nb4eY<��S#��G-i1�r�?��[�w?�9J�fLi����|���3�&��x`M�-�����)�
[}o��j�]]�����q4�=/�^n�_���_��%.WqYn�,o����%n� �7x��8�l���#�嶅-l�v���K��(4������8ڦL{�A��z]�5���<InC����7���]��`�"��"�Gf|$���wmt�ԓ��5��E��P���!�b��U���~.�[j0���^#G�冸�W��[{�+�d83lG1�̟��o�kQpG�Þ[�n�{L���^[-��G>�
B�����̚<�{�L����8I�����!g��d�ˮv�e�wA��/R����/J�d/>iC�T���t�
i�ʦDˌ`�
�<��%�Ddk0B3�`�}�y���B{����~es��5�5/TpC�rt�F�ӽ���U��J D��-|�"�wV7,�
k���D��Z�ˁߢ��z.z��gR�w#}�G�������"tw��s���{����F�u�y�������:�ZRQ�l$�V���@I�K&�Q�|�b��nh���I����6�
��[�ڦ��ٳ�"W��:B���F�䳁 �IY�(�|��?�$�d/��WE�	�
��Li;��i���� �W������� C���^�3uP���<�e�O.:��������z��V�Jգ�-"'�܉F���M\�x��l�E���Hr�F|{�8���,�Aw��ԟg��\>�R
��$�-
�\� '�g��s&@=!��V�
��Ż3F��-�~U�ڎ���Ggۍ��Er"��$�o"?m����ܸarڎ�H,Iѳ�GU����ޙ��=�֝�i�1Ҡ�-���hK��n���k��w����K|��m�i�W退5�,p�����i��&�U�k^q�Ý���Ǿ�!R���CŢ������a�R�������R��_G�e�Ƅ� ��.�3E�1~$l�U��Њ�jp�5�,�	a!�x/�F��&��*E��p�$�&m��(�������>���8OV���8������7M�*��4�r���2�B�G���Li��#��1��Bg��A'�d�U6���`��@�d
&k�zz����$#5=t�sz�!D�RR���9��H��.�9���ۺcD��>��^����RI	"�M�-�����"�����R]��Ex�&(|�e�"?����W��x.��K�ܐg���ޞ2XӽOG��� #/h���-!,�`�xK�D�>p�*�fGE���IL�uD�9 �3��.�~i�\(���\��ͪ#1���iA�e� �=Ռ���˄���a���� k�˵�^^$��Tk�s������.�>-�$9�'��q�kq��S��%r�t��	w��l�e��J���޺�yeR>S_O��uu�ў���v�.�n���*KD�$,��0��=Yb"�
�������-���3}E[|�h:��pHӒ{��La�� !R�$�JIR�d�>���BS��l�M� @��qYՎ����_x�}���Y�����Ų�_6���`�A��+������˛>��4�TA�*h��v�Z>5�6(_�[[�+���.B7�\ډ�,��Q��s�P�F�=U���[[}�S�2��,���E�{������m 0)�"�@I�hh=�r���s�00� Zo�3����ɼ;L�	�p�u��ˉ��rm:�"ޛ�d�:ެ�� p[0H��cͰ54�R���j:��܃��9�=�D	�jK�7T���F0{�z��ᯱƇu;�h�9o��=/5����@ݭD�4#�]���wM�_�b�P~�}���}���n:�c`Kj��������z�b�&�_Ӄ�a��f�G|^1���е#���j0Ԇ԰\4'q���f&��`un|������뱉l�xQL�K��C\�6X����X�������2Î.����.h6��2���>�ro����j�S������W���U�D�
	�3�
7���ˍw*�*ړ۞5F��i\lX¶�s+}�[É�Z:�z��:_��%���ɏ"BpZ$�SF�4�ZZ�L�r������_ *dOjM�Y-_Қ����Q��L�ȑ�=&�!���l)���q�S�G�u;���JOti�)z��)ZX�5�۸��|e&!�Li�q���3~�+�s���1�G�~��~7C!�?�u��*J�����;9e��":'v��B`c���������]��"|���=��Z�h���q_����z2ǩ5���["|,��3�$��-��ޖ*������ $]��x��ܪ�b�A۫�y�3ہ;F�n{�1:h�~�'� r�`��ݍ��h$��ϔ�'��Ҕl)�L����༩���>?U�)g^�dҘ�bٽfS�����&Y�6h:J;R;��V���̐�.�k􏋝Z;�V��A0�D0�c��z{������aYI*���L�Z�q�	������b�qd~� ����V�VA��c�>��ݹ��7���É��j'�e�/%���� ��w�<��{�UIq�`r�ΐ����	%�W�)�㩃):O�FP�諸��&s�oCe���b����fe��Q5�>�����V6�:.�~���,�A7
�IY����f��㗵 �)Io�?�/��OƢ> 4fgW_����ZW
I�4��D�@�5pKmfL�� s�<l��DBl?�0W�5�L�:��:�)0�w��R��JDwTI��.�C\�%E�z��B"��E&�b<3�N�CF�K��;!v��V��%�ng��d /�ӎ^�}ì'��y������m�Q�Ig�x��*{?[��&V���ɚ��h���	
�vq7����]�N�y1� A'��?�$T�P�w--a��˽����7��U֝�b�E)q��k��q7r�pZu������� �|�Y�7T]?^�,�H�4iK�WŲ!��qPh�.=�ڌ)l@n�/՘�o mQҖ�rw-����\;!��Wg#�(�\SwY�7˙$�� �{�{��S5Q�}���~a$k��E1����X��)���ិɟu�L���+0/x��^ͽ�e��2��q"���nV{nzv� 2�e�����AM�����ZN�B�.�u�q����m�cqaس5�0��&��/���y|ŜI���K��x�q�u��V����� �)� ���ґ�?��������/���N�|�!��$
djJ��p�/H�!.��/0C�j��2ڳ�xn���d;�H�K�5���JU�v�꘯~{��ɬt"k�$��掟�&�0��O��Rz�d��ճ;7l��_�� �$^��6�uZ��|��Jl/��$��5LLd ��$^�`��OY+Eu:E�!a�Q���" (���
����-N��p
3�� ���?ӛ�=o��8b|Ӓ���! /X���y�RG]����N������5w�4��Ye�u9�X�"�;u#��Lo������ˢ���T�\*����8��^?Y_��U��s2��#���@Ԧ��^�!F�&�S	@)O! .͎[,�
�����H<q7P�{��~����΋�a���'��K�#��_�U�^�x�6�K룞`�Iǐd$a�b��_�9^3� <3b�>n��Y55��xT�@���tGj'�k�2���@Z��S�g�S7���&>�a� *6����b3�r.��ZE#y:_��-�䇻�� �!v�q���r���Awv**���Y(�Ph���`�9>n�� �B���H�HWC��] p�a�Ww�(��e�J#?�����VU)��c��h�P�O-�[g���i�	Wh�M@߄.`¸WN�2uyk������gO�f�,~��/��RCKz?
��"O�c3�9��H�yȧS2��7��B�m��}��Ȃ�j�\�l�wf[��\�I�ڪ	{�k�nY�����ҨY���Jʌu��)AG�_75�|̬��=����z��b�4��y��zV�=11=P�z<8��ST�����hV]_,\�Þ0����U���E,G��Y	��'y
�诙ڲ�Dq$��yt�$�M��!�[��4fc����Y����^<&;����g�>�Bү�0^��5���-�m���d�-*|��d�=Jt�'�ʥ��iY���t����+�W�Ugp�pʀ���̚��1��Ò1o̝Iv��g����P4J��2}8�i�SR��!'t*��0��&ۿߏic���xh�A���́3���P]���m�d�M͎Y+�m�Cb �+8*|��_���y��}��2;�\�sU�Rz��v���h����� ��P'j�*zd�)%kVH�o�W;�,/�v�u�1lȲ*L���걾O`�������89U}���c@�S(��~������S�'yN�v�xڙF���(#Ǹ�	�����1�[ 2s,���}������c�gA	�*��A�+Y�?۴0�vP������� l�@�X%&��������>��&��K���W��حG(Y���xRLj���=��gֹ9'��� R��%�V<�32�����	��Di��N7w;�����ՂPL����V��c�,v���U^YVh@�$<����Y}7�OF.�o0��sΓf��%)sU�
ބ��WY\�{��:w�!�*�0������@�t^��ˢ��T��*�	��Ay����f{ſPƭ�H�H�dfx����`���[�nԕ1m���󕱩(����{�Q��oň�8���5l���[��5��+k�
ܲ��dca�S{�P
npk߰Qɓ�1�<����ؤ�KDj02��]��7����?�B%	Q�-�����ɖ��r�<_ n��ʾ�� �_|����Px^Jۗ�0��.C���3�T�7�������h���l���Ȏ��!��(�SF����q!0� @�H[��Y�U����Fe(V��'=�+�#g��D��x���h��s���bVϔ�{0D�ۅ��h}�M��ɂ��?�{�*�yh���<(>&�����Wx��[�a�[}�_��jFCGm���7q|gk{I�@=}ޣ-P#����(�����<k���;XYMC�H&rlC�u��DNE�?��=Іa���@O�}��(��J�\�-'���
�V#s'��T������ze:��S����U�,����K��{��"ay����B���%$���ܮH���[�X���:x{v\�-V��r�� ��+�D���Վ8��k�T/t"J���.�fy��]q��ě�� F�1��^o)I̠�U�t��e�7O*��W���]����W{{������-qWZP�8� 0�& T<Mח(Y��Ϩ��rTa�d�è�l�\�5Q>���@f�lR���wqG����805]@R���_�hë���!$� ��Yq��M&�]'B4��e�}6���޹J�z�n��e��κQ�\t�������J�>FN�U���I)4�,�J�b��r����R�=�a%��^uN$��@�ZG��� �lc�f��S�%Y����N�2`���߭��l����-���˳]�қ��-�����g�������}�V"޿��sR�g08@v����>i�M�����p��ԩ�ܡP�ߎZkl���A@�ք�����B�M��;#?�!.�r��zGW�Fe]�f[ǯ�dQ��-���v�u��+�R�Q�5�����M��ĥ�-���C�x����F>��/=%�b�QK~W*�ê�i��H$�g!�^�����Lh�6	`>�"���Q����(�X��7i���%�u�$�&��"f�`�ۣW��G�I����2�h�5>��E����Ht(�jՖ����@�~N-�ۇ��P�_*����Y�LF��"�z�5�pQ��i����s#+q����r�+�fAG��:�ۘ����S1b�~g]��h0���Y�S����2�3m�V�ą�=�{3��Ȩ��FܰtL�,$q��l��4$�Q�wwr4��8���G�,�� ��k��d�Ui�o���16�M�n�X�	��zT���#=�Hi�[����`�~&�Fvgx��
��*�����ʣہ��	)G�ݍK�.�H�P=u��=/6w	���QrǪ����)�	HQ�)"��o�
Y�/��m�Q���C�#��g�g������k� ���+�r�}��S�Sе�����>'n
3���3}ΐ�8a�o��I{&�(vn��I*\��v�M�h����Z�ל�Һ�ы�j���tS"��qH9��ۭMN��;�,�K��Ť�����P�H,8e��q����AFpՂ3��Rc�?)������A��Dm7��J�ts+5�5ޠ�cK��'E�%|W�V=���w ��OP���r�a�kHc�4��q��<!�O�����0G��]nN�N��:2H�dÔ���d���'!??Q�{���%:i�D"���4��p���N��>Pٮ��6h̞,+�L�2j��!��-��;o���"�?DI����T���;Y��F����3,��-�D�Y��p���&>^��:vA��c��#w�~���a�����m���a��Z!���b��Vǫ��iK��P��B�6կ�ݍ~���7LPCҚ#���1�'P��~�<KLUN!=oq���"�d9��(�&^@Gn�� �s�}��I��0"�	T�U:�Z�K��t{r�/��蕀�d,�f���C#�����3B���Z(>�����J0|��v��MG�г�m9F�5�a? >���g*s�ɃMD���z1��q^�ɵv;`t�G4�*�K-7���β]�;���Q�9���a�	�V�s �K "�[�:����N�J��UN��-z<t�}<w��=��T�DJI�~I�l����۪3�F
�_������?�^s�f�X�2���RG2��Փ;���L��ZL�h�WC����N l�����ST�,��X��]��+ǖ+O�o�?��X8�7�'Z �M��/�h��¸�>����׃S�|'�@�&[��HR�p�d��q0A]J�o�Gw��+q�O;Ou��T�O�a�8���)W���we}/�-{��٤˖d@dGDÒ�}�܃*Wl���/B��Sl:���+������� �w@��Y�Z�v0�,���hG��%!wL9����Ր�JK3βu��89��``��SJ�m6|�m�l����a�$�l�Ҕ��U�r��)9d.uF`0�N�]��k��0�w4�J-x�����V<Ξ�w�h������^jX��I���ʋx�?)���m9����<�v����F
�%�^�?u07� ?o��|T��13�J���M����Ҩ]���h��� �X�^��;��Y�1"I?d[�t��W�2��sq�[n�đB�E�S��?DB��0��ϒ�������o.��U]Q&�H�1���s �X�i�#�:���;�[$������Y,�0�݁�U��杏/#ͦ&�NU꥞FU]�N�C%ӄ��7�|,���Y�x&���4g�d��5%"�����N)���1Hl�ƒ���e�s�|D�#H�&�5K�Z�M��*�?[U��k�µK�΄����?LqVe���~ww�����2�
�2�F&�l�ɧ?��'y���_��:dH;5��e�7��A�.I���FHÔ���J��1�L��C�G˞/J*�֢^�Ȩ�_������H�d�d�2��:���l�H�w���4m�K��\�uA��Wx����K�T��������5���U�6�_r#{�Y��pǦÐ�A��Z6�R�mg�o�.M���Ζ�Bqz�6���$�హ_`�Ҟ�8����*�8<��a`ݬ��ŕ
QLՔ<��'n4�O�c�`Xk�;1﨓�И̒�����Q��sK]��b8��D���zϗ߾�1�'��a��8`��E-k �8��#[�j�_!ǰj_�Q,V�ʦ�6��P:y�d���k==8�|ٯBuG��r+xUe���P�s��N���Ec!�"�l���{8�u���}�ck���(�:f|���)5BK��{��&-u����'�C�W��M�4~��t2�������ma�(=U��"�>£A�L3����g�w�lZ$\�J��TXzb�c��I�x���EVH�b�����+m����[?���
(U�e˟�Ұ^���hj�M����4�����$AK`K`g�8�7?o����V�!`�Tr[H���G�:����+YH�|e_�:�Q��]g�z�p�� ��s.����[��ì���=��r��7°\?Vx��S;��Z��5@���g��K�}?�+`#B��A��N�~-p<Y�3@u]=���n��pu�bK?<����u6��,*����1���/��N�k��u�@�o
#WD-��K��Fxh��A�����:,���IMYU��v���Ԛ��R�"z�:p1|w��v
�K�-�Oro�/��f��𥜨�E��r�B�Z�^������U�4p�H����=L��Q&�^�2ǣݬ��Hlr+5�e��ħ{%������Հ����.�I��\�hOй)@k��y�8���1�4����@�̗?}� u�7�W618w� ̗U�e���vL�s�u�g� �]�a���Ľ*o F(	�jN�ǎ�R5��=��i�	L.�9�B�um!V*Op��|�>�%�Y�BG �:��#*�5u��H�_Q˨5}�^�1�՛�d�����7�Sm��L�/�AD��K'����kx�$4�{�H� O�(��>:�-�crf	�� ���QfZ8:��
�z��hk2L>�c�Q��`p��~Ү�� �nb�:+��x:.x*Q�&S>(Z�IC#���	*��.�c�F�l:�^7@bm)͈�"����%��*AE9�� Db	!�f%�]҇�*k}���x1s:fN5�Y��g�Z�1^	ϩ[(���q*`
�݂����P&�Hj��:U�j�˵6�����FtEB����q���U!�?#q0:��F�D�B�jxOű�_@Ϲ6N�;/����"���Yk��N�&C�<à�{ŝ(���)@�=����n������>5V�`�|j7/�o}�d�s��?[���95R���QyF�.�S� n.�N���%pJ����kԡ����5�dٜh	���D������䣌M����'/a�xNM�+�5���v���r�$���4���7a����x�xx�'�t��bA��c�Ij��{�\�&�|bL�Ҟ9x��w�%w|w|�4�7�pN���,<��s�l}HY��7�6I��RN!��*Q!�F�"�j��e�qUŁ���y[�@��3�����L��e�]$<*~V����vW$�A>=��Խ��&��hI$���������~��e��Aqx*$����vj�`c�'�-В~��FL�@�Q��Ԡ�+ƃT�9��g���]�gFeCX�J��TE`^��6K*�>���N�-N*����G���/�B2���+�j���/D�7�S��1mu����ȶKkp�������OpN�>���j�j�P�8��ˌ6�&���P�i������-�����$���jg�Bwnb�HY]?��ot���o��
'$
\����rx�ZX������Oà�nSH����P�Cu:����OzL;l~oBb��=�?t?\�*���$ayj�W�C|ד���c˘I8Cpx�è�+c͵��-Oc�<ʘ�Ն��G�|�w9ى%ȟ=|��W{d�!�� �E��ʶS�M����{L���sÕ��ߋʯ;S8M���VL��>�ֻ]����ͩC
Æ�T�"���g��%�`l7zd�(i������#O�/���y��w\�S�|�uM��$����`�e��	�G�h��>-�c�����F�0	�'U>����\��5WB�����!&a��u �6�`�48'�bA�I�G��'>DX5h��x��Ѧ�(�&&L�ƺ�)��^����`rw�����9Ojk���2R{��l�6����@2��72��nN%Pؼv��0�+cN�N0Ҽ�	�i4� ��𲍳S�Rx|��_�t�'�b=�������	�|�E
�P�E5���i:�>���-�@�V7�M��ɟߎ{�9�HƷo_��P �}F �ٯ/���\*�q�7����|ow!�*�}H�?;�F����z`��:��?�����.e3�,Y���d3^��&�U6�!\.���{'L83+g:-�2�b�i,�f�8(<�X9*���r���=kN�L�<�����=UZI�%��-X��b
��E�:�7ch�1Ԗ
pQ���ˆ���=;;g�:y�\��93�����<9=��t̽�er�+����S*~F�<�u�9Ki��,G������
!�:�O�L��ʛ�����ҵ\���m�O%����i�x��S���p��9(}8�;Gv��;kYI��<�E_�i�6�.:r���Ԁ^b�&�j��Ѻ$kN;��:����)W]--�91w�cGT��ѬMX?�Y�l3�f��D?곩߷�v<
	��ߓ��w�,qC�z���f��1W��w3�Q�dǲ[-qW�c1�Ԗ�M�nq\���NY�_�l\z��G��0����'�a���Wx.>����u@��,;d����vO�W��?nd �� Wg1s�Y�%H�-�_�픗�֢��K����Ѿ�����h�6wpa0MCf�4& �h��f�ȩ�1�|�scH���m�\Wg������_��ʩ%% ���f��I�jd/����O�Q������P����d��0Nm�o��i(N5h&�K%�w6x]H*��MG�_��	��d7����\�yÕ���2O�;$��\��v��j}U!8?��>��e�!��G������⊹����n��n��]ʷ�O�z���RV5�b��-�GIXw�.O,�cJ\���33���K� ��e6`���G%�x͢D"��{�P(���c0�M��f��"VY	x������yf��[��w�^ �6�d������0�X��0�[�aq��R1O?:��Q&�U�ՍRE0���敲��3C��lP�̴��+�����k<մ��5��������-���޶R��f5q�9z�i�6
�/��$�i���SZB�N0#���G�/���<}��(����Ҷ<U?�z��Ϛ�꾴�?�k-�۬��6�&9le�'�J�x:)��o�N�� �@}�����޿�R3R.L��/e"8�#����N�S���hVt:x�N.^#�������E��Pd��{���	,WH	d�$�&R6�	�g*9�b*ʳ{Cm�}��W��G!D�� lRE��'X��	
g^��G�w�w�l�t���<-d3���dS9[��l���D$�OI�@:�PW��\��1c���;���EN�0��U�`�Z��I[�0�M�RA�Ag��t��1���B솭&�f ���d�����{�k�T]��n(_��96?"�4[X%�m�)�Z�"���G�9��I^�jg�F����C�`u�kn��� Nw��,��5�,>������$����1D~)���@�n��7����>әnɃ�z��Nݝ����>���i�Q?��������đ�f��>D�:/������Q%݁�F�' �/��	p-�D�-�RL���:qvK�b*�:)�em�����U���'�u�Q ���l�5©a��8"W}��.�zSKK�$`G�4�iK5*��[O>�
�A��s$�=���I�9�I[.M�����8!��,��6I���!��&��N貕z�v�����O���(ӵ�$�����ؠ�2�h����X]��Vã��i�N	'����R�]/��p��4�V��i!���R�9��51SAE4c$���q��d�\�zAn2�	_�����w����G����.�j$��_�|�J�N�zi��喷�ޥ�j����>ՠϟf�d<�0b���v�=1����8��7��-��>��'[Xz"�\| Mc�r��� ��-�E)�=?�_�i;츖Hպ�0�u|��O�UV|������W9��!!ܡGm�̣k����]��[2P����1˃[�%�́<@��X>�}�b*��w�]�,[N?��g)"���NO��fB�Qw�Bp�X֦'X��\�e�o,8��ʡ}�!��3�J�2���<0�|O9 =к�wK��0&�:P�S3<�O�Z�4��_(�c�/��h��I]z3;�s��v���M��'"w�
��{�$M�l;�ߒ2�@�֓�q2Nt�C���3��>q�V���,�v�]�M�*��a�-L�W�T�Cjil�a[��k\�=��Ĝ�Q��Wٺ
� uI� eczDx�Z*<qV�(h8Ve����w�8 �e�`/~Gyb���^�Џ����f/����!1j?�����hTy�@u���Z͠%��qa��n#F��Y��#u���'�N���N�hXwB��b�g���8p�˒�3�2��WK�qN�c�<Y�P��m����sU�����@H(��σ�~�9.Uo��K7�n�.;S N�����T�>��i��l����{����z�X[�S��W1Ԟ��	-�7Mf�
@��JK�%��Wo�/d��h�^z�2�U��41w-M\��ǐN�,0�{M�//�L�u�_%L?E2�H�3�G�I{z�U�WP��d�Bw�����7�&e���Gc��(�}�SY@����X����9t=�_�Qy��s��_�z��e.)˅P�f���^�Ȗ	�eOm�"Ni�� <���`7�{�Sy8+�����Xl����E�*yC���Z�y	�D���!l�ʭs��f�/��$iG�P�{��2�b9��&Q���������7��	�-��}��ꝶ���O6��G������>���HR!��^ͩ<����z�Y�*@�""���;�N�N������#OO��w0lJZ �e� 4���o�XY�!8�+�c&62dH�`2�ؼ��� ~��ՁZ����6�J��� �K v��;ؕ��eK'�C��?J����]6/C��޲�H�ʻ���Ա����낙��ӯ'�SE\L��4���W�bx'FDO�'�s�>F���9��n�8����I�&�<��\��sj���5x�{l�K�σ��m��P�Ȑ̡|_~d\�(�E,gy��'8�M�Ԭ�a���n~g;���v�[�N�WSӷ���,�?�c�'�d"�{C��1ڗ��2��N���� �H14�_ڪ�شe	���t��H����c�eJH+�����E��|�GC�&R9Lf�����ͽ_�"#( �������&�=�N@�E4�d�j��b<��P��v�#�/Š�
RPç�$�b@�dQ�j��~3_ƶ!��k���f��/^������L�*�~������@����(��UX�����ʹ��,��ΐ���>�3@��B|&��V�~����Z��X�h?��ܚn ���7[Ē�{||�.��7���,禝�&O�@��&щ %�o|ԧ�F ��Lz��I)*[?T�M�(\�WXY���j�R�^������R��R���v�Zk��&�'�^��i��*�N�X)���ც�����\;�'��2{�Ob-$u�2l�c/V�B�Xj��&� -:-��01NS�XdjHL�����3��#jN(�t-7��^V�T�5����*�_���B��`l/jE��b�)�9v��n;�aڈ-��ه�!�$Z�Ja^~`O�G���;�������l�O�"1�O���� �~��	$m��El�.�Vr��Ig��d���P�Vw��JIɑ�4e˯��o"��7EG2�A��e0�uS��g_%���HEX�01��c����1s��h��҃��iUU�U��*|���;S'�/6��V�{~��.�����X�̎��ƌ���A6���!�^}�^�d��f({�,�� ¸�^]��S@!��.W{l��oEa@���@�ӧM���hNu1!u���$��@�Z��^;�ơ�
� 1�N�+��͞��u�` q��U�ό�Gۡ��$`N��D���}}��GL=tjfu�qL��F�՝�8[���3eE7Q�$�50;��_[���z���F��[mQȚ��`�@�!����$/w��F�h����%u�_��+gK�I8C�B�x���R�k�lYoa�e[N�K��Br_� y���#����8�W��/}�j�şO�lr0�Az��@�kp
�C;�~������	x0��@����!�;�H��Iq{)C�1NY���%�Pɭ�L`au�P��Ղ�I�\m$;X����dQ4�^�t�����\�A���M:~�W
��`7E�s٘��|Y�Ų���r���R�ʞ<��44�V�gɤp��:�o�D`�SY)�;��G�G3d�9�x�ǔ �e�Y�D?y�Ob`�كRn�Af�P�o9z�;���E�h��
�g2sr�8�?7�8��T_���W��g+ҕ&	�A���m�����|,:s��2���$�L�Y%S/��]���}�e|��@����1�e!;�u4#׉S��1�!B܏\p#*�S�B
�0�;�����y׍x��w'�C
=��N.�(��|���+8��]�0At"���͍��ؑ�=�h����ƨzb���ϫ┳������kҕ�CO�3/�Դڐ�xV���ʃC!�
?x�/���&j�*ƋLh`��H�����ګ����N\�_u�i�Ə�t ����I��)�~����f�l�Ïۈ?�#�^_�� ��W=�dαZ#�(|�?��س#��Ne���UŤ!1#�t�:�����HՆ�r�������ߞ���|�B>-H��.�i��0�O�x�b���m��5�$�D`Xm��j1^�ɋY֖Dl�z�o�t�A�����qZ+�V!��%|?��+���]����g̊��W�l���t�Z��:�G#ﳅPA0��Ȩ%�)5�df���h�Իr6Z�D��#{���Z#����]YHl��KLC�x*y���ֿ&:����˧ް%�<p(H��`E��N��qͮ.�ͪj
�]ߤ��G�ו| ����T�	�ӊu�q[�"l&�0xb����";TVϬ�a�s���.�*ѡ�Q�C�:�S&ق����u��G�槶���
���k7t�
r�Y�'7ӂA�������^�qEt�L���c\�!�E��I��D}\�*yĪr&!O�CP�-��j��=���r[#�3��|�g��&�j+VB�P�J�R�ڑ��M��⃲֪R���"=U�c@�%Z����6v�u�OK��}��P�j��<���ʼ�P��ڦ�RM6���ٗnq���Vg�;������lŢ���θ��������x�썟��h-�?��O�?0$�T8�Z�&�
)�64��	�������J/��*6��ة�v�nfǹ�ӒyF��;���n6Q|����!��c�Q~����{� ^4X����v�W�9�O���r��&���5*��^ؠ���e��,�Ō�c^#y�x(��w�~6g<-ac2�=���~�����sO�N�l=��ik`�N*I��s"���|M�-�B�P����m2�bhQ�T
�~҂��h�!���ʝ'�)�����?��BI����̴F��i����hZo��1̗��e�?^��k_m�Aa̪��>:Y@��(e~y�1t3�+eڬ�J��\
�h��]˙SE�i%�9�8_� ��Y��#Ţ!��/���@��|h�0��6Y����Z��;�����P��acWwTEĦֽ02�s��a��l&�+�"�_��W>X�:��ϒ�!�Id�2\��eS��;�qO�6y��m�Ͻ֩}]:u��E8Ǔ��1���"/����{w��]8�m$ص|w���jVݢ� ����퓡� |j
J, �:��q~ �r�����훻��p�v:ϧ���h\ ��J�k���Y�V&�ݍm������5�1,O�V£��u�y^�#�h�~��Vn���
o���KM�z�a�R��A���O�(����� sx�$0#� �GZc51�x1�9�0�j���M�����%�-�d���ˁ}�޸�r�/��E�RƷ%��Pڠ r۾�ܧ�!�!�R!��tZ�1�E��{�|-D����G�nɡ�5ѧ!g�^F	�z��Y�Ki�붗`0#f+J��(��W�A�uR"Vi���b�����u
&��<x���U����D��m��
|$m�f�6�Ʋ�-U�#�/����ɬ0���n�D��*�Ռ��,�0B���E�������wxNb���J*S�g �f��|�®�*�̈3�s����n�xRƈr7��xE8J����)��!G�;��C)�bC�q�'��
���-7'��ǫ6o�@�"���Xߜ���h:���C�׋�����xC����	c��?f�����q��A�xF���w���Zh�,m�ب�BRS�X# ��

#�~)t�i,�^�zD����-�%$}��=quaOxک�Ix^��:0Q��`m%�ն�('`]9�	H��ؖ��,M�Y�gp�y�G�t���$�����wV���:3�i?��ٌ���Ny��Z_�|�#p�xb0�ٖ���<ȇW��: ��2X<�	Pr�7�"K�l�[9;�]�a/"I6�?��.�qu�̎N8>:w8}�(�-㺘
��ȵtrD?�wj
�D��ߠ��e<����X��sb7Lu��Q �c���?N����1�DEC�� s�	�?��O7��"g��gNN�F���A�Lź��\���8W��q���wge �a1�$t�*�(t�M첛C��).v4��1>�-5.V'*�����[e�A�!&����s,�*�TN|g}?����Cz�����Kr��hbWD�h�Qz8!���1��gP��G�=�����C>�	ZH����R��'����Ҏ��1e�mް�m�~y�kd������v�l+�Dq߳1��慫�;d�J�#���)�����M͆�6��1��gK�_U����mD̔�	��e}�q��hxVa5TF	��D�fu�m(�^�5	ߙD>E�@ota�}^JU^���}����
k�Ҏ���!*�;����W�N������Vo�rNĬy�<������03!@��}6s�8^4 g��{�
Z��Q���I���	:�`��,)�����4�E�G${�yPq���ls�;��#��/R�
]�����=ݠ������ʁt������&<o�*�;���!�4e��0Zߍe��3�ɐ�B��/��h��^\�v!�޼����5g�Y+t9��0�p �0t���S,?S19�5�'��E��#����[�@G�<������0�ˎV2O�x���g�>U���ۥ�ڥ�F4�y=J�l��P������`٫���/d�a��r,�c�KD�O uG���/�Is.��(f�H�ڷ6 q[m?6W�(��4�����y��(x�����kVB�)]��m�%ܪ�X{&�U�Q����l?�&+G�ٮ��{�f�s7~o.�����G=O=ڂ!�V#4)�8D]c�U��}.+�7{����JZ�y�o`a/;3eBM�O�a��N���A?���}�Eq����C��C��=��5�AU���P��u�~{ngR���wY�;�@y��,hB �D<Y�\dLl�E;�2O���)�҃�n! {�uG�"ϋ^��~���	�5�"D �O�5Y��|^�P$G�vRZ�?}	�l$��54N�o�I�=�W*P=�����9q(��kw�\i=~l�S��9��&|08�!�_�S�������ةY���i����#���]%�И�4x� rN�����#]��pY(� �=_�[ۡ�W,ܿ/�ϡ
����� �@?BQ�f�^�ȟ�O��|/S��K�x�W�+%8��@/K4"��ջ*(#ߕVʷ�{o�V�!�I��<�L��aY!�&���΍/Ģ|h�B�KH��u.TXd�ҏ��0��������0��fI֎� ���Σ����rr5�K}= � �dFG���hw�+�\����JA2���;O�}=�]W�SNx��KЅ���xKcZ�vy���P����rOu�y���q��Mf�� �o��pY�Q��M��V��g���?�0��U�q=J9`�M�����Q�Ԃ4t�6Հ8�������3g��]���Ox$9s��W;i`���)fZS�Fd}��oɆ���7Z��P{���8G�g���x�1Y=;�����ab�$�~�9}�S��tح��F��61w�~z,���0殰�GS�4q��>d$�#�H'$��<�5��X� ���oAW�s��RL��W�3D����g�����O��?mi�*�p�,�E�؀ͤ�쾦=_+m��7���u�kE+�tM�x͵�N)�H4�Ҥ5%�L�0I�A���	
��Bܧ�����ɕ�D�,4�	@�xS��P������`56ŕ[]�|���@՛�yW�;��UԲ&�f�8F!�|�b�-I�>[?����ٚ.5��W;V��|�c�"/�-b�M�Nۥosb�f	���t��`�C8�O�B�G���ڹ�gI�׻\�(ct,"�$�ڥ/]A�yιN���X�R��X�U��{t"���Z7��ϡ^�� ������1��~�CI��H�s.pL�T���{e�Xv��8�YG����6��ڧspTT\K���Pv�,Kwݬ�q6+h��l���u�fO�3K�����>���� I��
퍋_U�+�yb����"���BSs`2 ��(J�T��M���!�88,�<�n釃��X���B;�^��Z�� uy-�p����`���%�2��)�<����SԱ��$F|�(r���l-*o4h&����t���A:��%
_ubP0u�LZ:?/7]�$�#:�.	����#;Q�P����L�j��٧��Z^�b�h'����	�9��)�'r>&�- �e��m�����9�u�=����<���������{.0��/QD{d��]<�)�+�b�L�3.���7��M�b��)� il�(�іĠ$Y>�rr$Xb��C��B�\"u����<W$�Pͮ�_���-�e,}��������Iz�x���U�<�����V��=�j1��u8�9��Z���%�,�y�v-X�)|����$O7�fRer��^���k(�Ƌ�b�G��S(����AAO��Zh�j� �p���Jur�W'��dq��&\	��$�(Q��-�>���V�W�A�J�""��9+i
'XM�:4u�R�k�OV��L_)P�aO���X��x���Q��J���o���I�0,`����2b��#�-�����te�#��hw����	�,T�*.�~_�\z ��2�̡���Q��?����%���="���J���L����"�!���������t�$�*cq���x �S.��4�s �I4ʹ����f��ɉ����[gRo`�y:��r��#E(?+.
~٫����~Y��D��n�h��Oː�:�EKX�g_�tZ�����fׅ����j7��AZc�A�������{I��7gY��ȯ���F�Sa�&��d�tk���7r��$K������7�Y�I/�q{]�x"��QY�CD� uE�9>G?v��Ix�:���r�7��/�\f�|j*<5W}5�,�x�[��B�D�|���W��"�q���l+C+|��g& ��3s.Y�z�C��Jѓ�z�,g!�X�<DD��	?�]���ԧ"+&��O{I��\��?�ľC�2���a����;��_J�a�x 	�!F�!(q�`%�Q�������{1(�1��j�X�J�R<pԣA�P4C�8q�3=+�K�p]k�zr2��~8����g.-��'	��B��i�Sտ0�5'.�Զ\��Gk�
FΠފ��߯�\j�-Rh�K�)�ka�)�\ �K�}h:P�v莰N��;��&##mo&�*G2�OT6��T�&v�cE%��'��Q�!��ed�1;+q�؇��S��/K�HI	fv�o׷ɑL����^�i��K����㾝̼���D��:'g��:mM6�+���G+HP׸&w&�5��u`ES�+����}�n�bx*ђ'5~�&#Z��`��ZT(D[3��`����e���8��#����~�����ʳ�<���PptE�rD/���R��4� �>�ٖ�VMUx�r����\�s�t�l3�<Om�S�x�tKR��目Ml3M��I�_�9p�LR�;���83K��H̄�@�B5t�Lc�0�]�	�ꇫ�l�"h��7�)\~�$����ZoJ,bC*Z�YGnaX\t�g�J%��~܈�v�|������I�v�Ԧ��~���v�c@i����>�$��v���nT#���Bɒ�Pjf�ce���T8�4s���Z��F��f��s��7��������r�7�p3m��	�����}��X���6��#�"�g3Tlɛ��՛IG�P���~��=��Fs���e�B$�y�3G^c��#b�ӦH��+M�v	��5/�'i��s΃�EiH��˩�+���?��`�J��-&t�*��3W�$��T��Q$+Q����R����
�u�N�q�V[U�/w������������@�s���w���[(�zqݭ*~�
��s��hu�R��9����q�!�ro9hLz��)
3����M��ڣKO�Ǣ���Sz������m�f@�轼��݅%ns~�ɗ�JަwOtI�e���v�����)���]�u&�Ia#'�W��4�UA�������F���N ��t)�h��w�p����>d��꟪���r�?����-��1v_��!�S����IjT���]��sy��JJK�����7?5c�/k�T����(`��I����!�����:�����?ut,Q�0���������ע��:�/�ъ0
_X�uy��V��+;.��9?^P��0���8���A^�� )���M��&&/�ǫk���:0˻rl�XR�n�1���	�:���p��Jȡ�GQP�� �%@]�U�*x�zN��yQ�f�I&J�M
��<C�7��K���Ek��x�^��V�yW3�����}?
��F�o�,����H�w��S�� 7��E�%� .�=�85pz�nǠw�)cB0�K�*�Iq���TZťU�-�����mA��9�*Vbi�39"E7Nt{�T,�aC�Q5X�� '��2��yNR�&�О������]��k�-+Ӵ3�}	�5}=
�{h@�F�;���I}a8֓n�<t��[�G�g�~�h�GHC�����oS���Ѥ�`%qU�U�D7��<0q���^:M*�_sY�R)�	#~��<C��NV��:�G�4H�1KPT��b��@M*|A`�a�B(Y��`=����z�7z7IU`��O ���R�(�î�p��gY���8�h��#�� P�_G�DZ8�vG���]&��D* o�]A5�[�v�J�8�_��$U#Y�W���N����ڰ����>y�=�F!e����Kj��Ь*OC���U�FXff��R��]��,�2P	79I �k%9s�"��pEk:Ԁ_�f������� QQ�*	Kfz�A鑣��F�!k���z�Ҍ���H�2 *�yvj�=���?��*yt���P��e�_��/�.\ d�ڹ��"���� �]	7
yj���,��G2R�s�O%��޵\�������;�-��R ��"u{�)8j�mG����${wKx�]�I�5��qO�d���|{�e���s� �c�b �3	�_o-�.�� ��Y�w����|9��4�Ad[�x\GQ��,ߕ���M�ˌ�0s�Q¾�\	Ps�/dn��,��G���������d�dj!Ob�����Pѧp�cm���3�g��LpTW���g^�U�vErF`7��W��9�b��u���\�?�r!b��$p@bt<FZK��o��w	�eh�qt��g�D1X�u�V\j�����H��.M(��ͅ�擦D���>��&Y	��s{�a�����j����{��/K�L0��D1W#N�b�aX�?���"T��hrcQ�e�ZJ�fӊ���(_mϐ6�
v	���w\�K#h��}=@�HO���uڨ�G�	�g��JLqJ�������-QS�Uο �����>���.!Ƚ�����������Pn�wp���k����I��c!9�U�6�'C����4����RX�9c�X��
��4�V�a�e�o`�7�bp��W�[�/�8�� dY�Y3hd�kf�J���p`��Sȏp��$��*S��%>�!f��O�-��$�p�DE�O,Y���ԫ�R����t���N���J�9���L�v �~Ӆ_�Iy�w�<�}?���Vjňm6��ߦ��9]�w�*����A�Z�����
���w�oZ�֜��k(��57l� ��%��י}�?<��s-f���ГF!F�1�v�&�R��_=��kH��v���P��:��� �Q9E����ǭc�$z����������Lz-o�dǕ*ST��:�q`I��ڊ�^g���Sku�y�A����]>�SĺY��������0��Z�*�]�6o�1�|������c� E}2�W�ag��T��i�?+�I*Z&�Ǵ�o���x�|�sIu�N��j��I�h�qެ��z�Â���1Q�T�̔Ga�s����15O�pd�k�ڛ�N-�e@�{PEGKap���&���\)�^%���%5ل�{z3se�{D�&��F�QnǬ�>������hvED����R��kvx�jʫ�x!L���3����]�މ)� �>f+_($���笪�k���قE�*?c�g�.F�5�Hg��8��a���V�*Uv�9��k����Y���g�
Vm�0��"1Ɯ��u0n��VIO!��zh%�m 4��K���[�'��� ����8Z�9���K�C����'�h:
Ή��8u7��=r�_��d_��hy��N��$Mv;��)AQav�Y>ߎ����5dbH\-xzD�Mf�r��a����@{�������%W��<i�J�n&�F���rK~�,ms�Wh�\�$Oᝤ[��~˙\N�1�/LV�,�dPl(�?�l�+XΜT~��.ɽW6z�,�rn.��wN��|X����õ�.
�O��Sz8�ڀ�A3����#`i7X4�+e<j�0�q�Ci����X�ƃ�kL���ư���؝mkҢ�n�=�V4����/�.X�2d��H�]�r���Z�Y0V0n�]dw�Vt}���6`ɠ�_#8'Ox@��;���AQ�X����Ә������x)����]`nty�nx߹�І��_$_9?�-
���Aa���f�n�����1������6�E�h�Wĝld�W:�¾qt�8�O(:����?�4p�R!v�཰�s��mpE�QB)�@�pl�Qd�E7���U�J�a)���_�B�Nr�����,x�F�I;<�������=Qbv�L�>��Y�נWve�a
�p�~�[��]Kc�弚/�)������8�G�ou4w��������ZG�D�����u�M6c�EK�V�V(3�\/��P��9�����F5׷^?�z'����,˂M�����E߀Er���F1��c�	�
�}��B�����;���nH�z��J
�I��A���;h����zj�{3$�$'[��n��)�#ݰ������\����2����K-q5��N�\��Qv����>��[���.�=F���������S�l����,���S�b�4�7�u�lv�p�wm$0yn��ռ����5��rܫ����V+����g��cc����p?����Wugtz�1�^ҕH��S8t�5�6#��az.rОv�?A:�q�+�@���V{mG0�9�'>���,�y^�o�:sJg��y�t�"�6�tA�#l��R�jU�|�G��3��h��ѡԦ^jнgqO�}�ʕld89�ǖ�ZoX6�4s��ds�E*��&����zX�:3�m����DV�;�c�s�2O�wC���V�4�۪1X�S�7�����i�ݓ��� h��(�0A�A�^39�L�;������N^�x����,��Db����!8�>�4�q�E_��E�D���H�@htq�h��g<��4n���:{�R��!A�m� ES�a�������u4贂z�Sd�rq�Vݘ����P_�) IO��!����A� �[L{̖d7�G���;�)d.�ㄬ�*���D\�Edt��[3L���9E�aހJ������ �N�L�����(\=��+�Y��C�G�ಊ�u�&�����u��'��<k��a�!�!jڿ׺��[��0�r���z�z�K����� 2�`*YN1O�;��z��i���
�J[軣b��7�6j�!��8���f�� /ƚ��L�(l]�<�zKi��z<k��r�V����9�{�s�����M	t{h��`�k�m|�U
X�p�NK���+%^c_z�
���)�A7u?���$U�K�2v�Y�6@��*��Rh�0VO��8��}"iH��;�T����0*�7���=�l���ؕ!���Ԟ��x���4���&^Qm���[mdN��(��Ŷ�V��� ���_�Tq��L�m����60�+�T����44N�t��r�v�0��2��M��CE�>�v� tD����E�3�8�U�D[j5f�\�����cdxXRKA甩{>K>I6h�c9�[���-��X�VnE��k����W*��G����[;<�����&Ia��H�촰�V�'�?��iy�QS �k��	�w��a���O-�b��E's������Ai���uc���dZ|�	*�����]"�:�AƉU��z��8���{�0z9�nhe�X��$��ҳ�%���r
�rG�<��ߥ�����P�t�9L�`%b�Z��y3��;6m�:?�u����L>5E�x���̄Ժp�8�C���dzL���A5[�J�6x�Y���@tq���W��w� gE�$�DI��R��O�̲P�V,yy�o���c�T��_�P�I#��X�t)q�t�L|��?�kr��9���sy�z>���Lj�t�8�aVn�3P
dz8��|���f?��yT����Z����w,9�2U�9�E�*���۳;Ϛ��쯛ߨ �: L7p��{��9i���r�2S���܂,�b�p䅜qW%�#���OH�x�+H8��'MPZk�DeX��;e���a���-W�������_�E�%���3�v?㓺�%��a���2Ap��*�S;3�z�t��G�P�M�m@�;uox�"�t'���p�5ش^�{�5O2�qd���6T(s��8�=��|�� a��	�������������^$Q����T�j�w�ә֗���80.Y��M�����G�ߚ��9�Z���Q�H���6�n�i�[K��G�R&�K	D���;'�����7n[w�r��G�>��>'��1���CB�f�$A]��r� 5E^8r9���� VNV�c8�-�T�?�F�&�S�z��'�N,50�'�k�x�Q��S�E�kEoK��rk�������5|���=�S�1��\��;U�Q{��i#&��v�Iz�^e>]v�
�q����J6��'@s%ݍI��DS���\��U��Dt��b2�UX|=�� ��;�]�,���R'j�i߽�v��G$�O�I�E�>�=�o�~����wI���)�n��S�`H�n��8��;����ua��v�n[Q���( <:`��qY=�?�z��'�g�7jFDغ�ö�������^>��b`�s�ۋ�f�LKa!�ƀ*��Q�j���jQ"���c�7���U��n�_.�99Ƒ2�$�ǉ׷�{��fBq�,�6Q{f���5?���x���*�2ݓ��?��a˒�X�64���t��P,	dQ_�)��p�w�T�#8�&{�+��I�aW��>��"oC~0���x�����S�p��^�����b�?CzM�:�w&��E��K�H;��XZ��sN/{�|=�.��u|~E�)be�z�`4��E͈��p�����h��[�u.}s��(��əG��P�Z�оߓ����Cˉl\�?<5���;ǑWgV�.x+�HyVޗ��	�MQFVCbp�HZ��CD��;'�-#7�	u1��s��!XM:`�?�����xX5��C�7!�H��P��:�9�)Wə��M��DF��F��,N�`���5Q� %n	b�%$[���P���[���bw��2@+`�y�d>��3�d��[6�~�Y��x�$:��\G\�CC�h�n�XOM&98ӂ��z|}��Y0
�=�О^������{w	ʓ9Gۄ*Ù����%f�v��q(2`�l� a�j�(\�J��ϧ�~�i#^�p��`L�YfQ��y�B� /����t��:X�D�xB��}O����������m-3u�����?Er�\~�.�����w`� @�Sk2--��~��k*C���B�!�5��ț!���?��@�%�i
.]��*�E�s]��|��1�	pF�QN"�捾��#"W�؃�'���jG��M��0���K�L�������3��^eͥ�7nΓ+z<R��� {���甮��$n�����s��5Fˉy����g���������4%�
m�xx��|�� "[���i�ܽ%�:��_|2�k�X��{�N��$H��[�C_��-�������҂iy���$�Q�K�S��:�P��b�G�(�8b��Q��20��#�z"�$�����ڻٯ	��S����W?,�����k��WH�O�K��_0�j��h�Kx�W���벤��E�-�X���YG��|���yR�B�Pc�ldչ=�&�(/9^|~�S+vxO!9�����"�f#֯����i������0�ٻ��K�?+��q��*�;�ݍW߿,m���"�h�N�P2�$�hujĦ�匠$�+���'( �Y!���B=+H�ãJ�:/�	�D9	�:�PSG�p
�Jӽ�z�s���VQ���<�{&/��{�y�*a���x������#ِ���
��O�H�я,�Q�����95�3Q]U(�m:���?2	���2��G]i]&Ft���O�k����~ȁ^7�14Ƒ-���FY���%{�䝀����Ն�0��G��&�k�/7��T�34/���|�}�!(�Rof�4vʒ`��.8}���e�}`B�E ��|�s�L�ʀ�����6��Y��`�羽2��=�
c�:A��P���}W��;�s�D��[2q��um�	w�h���"�����3�f���/�90��R,����}?p�A��D�\�6�)�;T����W7`����f���)����9Ĕ܊m�i<�'�<��o����ءeW�{����4N;��
�^ؙ=��l>'6�����P}�t�*���ZI�¾]�p�������>�A���dr�<p�a�],��	�g�Z���KRR�[�+3�K����=z�M�+�(s���3D��(�(<�g��8q�LtJ1Ao����}S<J������d S�X��M�&����I�����OB����+\M�����{�I��0� �3�ՅSmJ8q��#O�43�1�!R0áUU��J3N�$"�f��?\@�#X���-����T����S��ȩ!(+`��!��^ldSC�S����������X��M[�8Ҽ��e�̠�CC��g@��MU��D���T�vX~O~�@�Q�`���cSC���?����P��S.$��|��˼qz�gl�������m�M����!�����w�ŧH�%�;� ������/X-<������b��Y�.c�{_=�8��&`v����J�oGK���,��G~z�M�/`��#MD������_rߤ�_��.��iZ���K��|*���J����:�����	Y���q��6�[E=٦P0B�SI�ά��5�/d�TtE\�%^���|#RAi-�U6��&�h�S�1b����"]T��<Jb��a����aD�R��J.&�c�'���P7g��P��4��L�=k	R|Lt�X�����譸SG�]��kux��
MUo�FO*�y��[gD���߰�p��6�_��sl�4��F�XܹR���<�8f$���1�&�$�>?��eXs��.�u\7<�����h)�H��8���E�ԃȈ�rf>(���$&�9�f�֟��m�H��	5Wr}y�*)��v�`Ƥ�E�R ������Ɨ��m��A�u��P��"�Ε����Ӗ�5��j:dp$�6�i�t��?�2Z��E?^�����ߕn���Z�I�
�f��a���u�/#C�?�v���oy�Oh�H�����]�Ӄr7���5rܾE�6N�c�;�S��J��r2˃�f�C�,��x��02/+`y����%�"1�*� gZ�<��C}p�](/����Z8����(��wV��>��_{b.Î���$��4��C�O�n�B�A0��-�m�N��i�.W(�oW�����Q?fu��M���r�o ��9�sgH��5��S'Y�>�kK��,Q(@,03��.�1P���k���䕆d2�YUB�;7Ֆ13d�(��R����0a(�e_�_!j�������T��8�a����.H=��/���1[dʉ$��ust�tk�'ɥm"@��U�q��*C��|�C�C��-v�n���x��Bu�*	޻Ѝ��\.��	r��
�9�M@��X�|i-�䀇��ڊX�N�'�$�xt���c�� �Ί ��_Dy��̴bu�W<t�����o,"�vlt���u"���:��`��i��(��t�5&ۀ��/>�Nr�;���%܉Ude}d���k��'���OP=�\�}w�I�<��1}��p2aq�G2�n<��VB�!�8e4�ZA�FbB�<؛��\�"E�&�c0KN�d�V��y���O!��"�"�m��|J��V���lmq"��w'�1�rt]LmG�tĂ���c��Z?yr���p�pw��`�]>�.,�U�Y��v�R�U5k\�ۨԜ���8�<׬��5�°!��*l@S����J�m��]/���`̲���� ��EO���Pk4X��r����o�P�? ��)nOym���|���
|�y]�wl�I2W9��;i�s�;[��8$��j�6b�X�>}��*I�X9'�c���c��]J����P�*��F!
��V��0�ZRKd����#��:����PW�B�S���K��c��U��`D���+&9�q�������lJc�C��,�n����y�Ԏ������U@g�JCa݌1K���`�36Yl�XzG?49'றh�p�lc����Yf펶E+�+�3Vl�%+]������8N4�8#W�v�}��4B숇<!M�>q�Ɩv ���������_�5
	<�&�s��j,�:n�P�?0�bp%���>��x��f:�kTʈᐮ�I���mv؝Ũ�4���R���X`��R�ԌV�DZQ�0�r�ӋG�j�,/QGZ�xn��Z��2o�K�J��[���{�R��(�'�⼀���J8�c��D��q���e��(����e�x&���t}E(�5ibѽ�+?�kW�1�K�o��Ú�?O��6'�\�^D��m��q�_�{`�4dNQ��i�u�����`1�ޞĞ���=&P���fzR[���2�E8��|��"8ŁKW�kc*/���l ��.��ٽ]�?��޹i���$1��I��b:���s�r�X�Nۇ��� ��3�"��K����TG���2�s�b�����.W��U��c�_�:�	b�����sF)f��jC���j��8��
��E!�r%�PV!�{��^��-Gݶ�8|�r����Of�黶����V�C���4������T�_�pR�������t��o�e���������2�"��̤W���r�Ш�:�@���GD!	;���7S�@�G�vk]ϩO��&�o�ꈾ)2��G_�"eW��o�1P�q2�<ں�3���⭫� D��nA�������A϶m����7#�!/��VT,t?E,?��b�`��x̾����`e��v����򁤬B���:�g�~���{�iô)��ǩ4}h��R>܂e�
�v�Qg�^�S.��<�eM�� ���1�罈w�Y�2˿����u��M��*�^n
�A��_����*� ]͹���n�ڐ�;bI��h��E��tijpYH��?������\&Y{���8�n�!�]`�'�¢xL�MX�cP�F�:�UamdM�=Jw�M��-TE�4Ԡ�VZqJ<t����i=���Z����J���̎�I��"�<��,�(�ə��=^b�ܶ A�d~��"��7���fV�Ҕ�{��n�X�շ�^� Ζ2�υn�0tL����V	ޓˤ�dB����f���"�	3���6=�����V��Ck&IpDܹ�����<�0r�kڸ����{9ǧ'T��9(��aԛN��L����RS9�*�y��?��|�]��0Ie^ߺ�!&�$�h5��
d1�b�7�.T���=4l�� ,>i������N�*(tm�p&�EC�A����_��/'�30��e������=��ʺ�,0պ]����F}޶��?!>Qا�q�����$N��0g���S���$f�e�k/8T���L0ÖY�� ��,��F�rֵ�$*Q��~��~!�rK��#�Uh�e-
�܏�r�U�Sg�,����Jk}̡�I��|M	��׫.�PB� �]���00���}r�i`{+G�������7	a�I3+�<p�wH�G���5�S|��r:�.�M�_�����!������
����>[*Q��dw�V�Y�s^ų�<��32�?�]��3I�m�X�RǲJ�ˉI�o��{4>���JpvUX�m�ۮ>��;�G7	��zů���Xُ�;碢MS�T9I�#6��)��旼L�?���tZ�1uo 澱u��{Ņ%h��%FH��f�5���M���;H��=Ѓ�\C� ��?9�,Ī�0X��8��c���t����*Z�C�eB��Q�H��yzV�|����N��V����Q�@9�t� A��9oUc֎�J�j���I�Q��"�~@c+UD^��U|��ā,j.�
H�����:�l��[*:�S,>���P
 y�	��u�{����g
N��Ǌ����'H�S�I|`���nD�����Y��m���J�U��	Tv���C�$��$R������%���q��/���*8����לL�8w�HWƾ)IQ��q��D7��Cer���m�,�XH��c>�pS��K��s:	J.&��IJٷ]�P�7�3אZ�g��	��٤y�W�N�j�;l�\�F�h ��%�p,TVT�j0���v�>B��5G)�c�� ��iwwv[y�_������KE�Z�[�4h���x��/�n�jYjH�>�C��H�ր�^Z%���4y�7S?����5r�)��>+>~��N��� �=��D���/V�D�*$�$�׳_Gf���-\F�-YJ�E�l�h*�fk2��������/���r�$X$`�`��|����1��������o��z��|"�χC{�8������d��&(�CH�k%Bx�&�7��M��9`�d��g����4�mJv��<F!(��ױCpN���	m%i���fcE�t�wHW��R��0����z�e�\�ew[��ƾr%�)�*����:@��e�PP�h@����GN�Re�w`�X]��0��yt����3TPh&#���._��S�(��-��r\k(K=���M/?\ ')I��pTƷ}�Ю�+y/	
�QI d���/��@�5Z���P�TgƯAz�zy��P�U,�O�v{�2��j����2�����Ɣ?�{:(�`��5��x��ȯ�#8�3.%2S%�e8}�k��/���+rw:Ҋ,�r���}�2n[�][�O�u��.�J�C��=Ӵ:��u��޸��BP�i�¢�����l����뼧T3�q 쌒��n�/a��K�$]˲N�w'�����p�z,q$!�D���P�aI���D�b1,�g���o˶�^����-��(��$f�B_l�^mtFp>\.�sS��8.�����ẟ�*w�'64����C��e��>]�5�H�7��F��}/����z��d�S�0�:v��p��.1?����P'h�� ~f�1��F0�Y^�"n��]�w/�ݗC�Y�@Q�x�48��l�|���W5�9>��tgD,�+l��3��縒o4+�|�q�hSF)�N�#wJo�7��qZ���+�������	;-��UsOL<K�8�#U�A`�E��+�0u'�
�la>Q�U��5��d80.�2*7�ۺ�/�}C7���ĕ���Ik��Zֶ��ES\O�0r�ZU�<��J�bv���AQ$�/�73��`<�l��g��D�Y��G�x�^hg+l�8��2����V�=n�~~��[L8Z�0Έg$�*V��R���b�_A��p,�̖t
1ͦ3�]�wtR��^���h�ڢ�G��s�_^,�Q~�=i����m��l�P�&	xhB����`��0��];�����z�P��3P�}.��F�ƘOr��qa��N#�iW&[�4S	�k�>��_b�F�M�����drJ*��$;G E8��F��(@R麾���5�nQk|��`����5�彂e$4V�7���ђ�Rp�y]��0#M	5�Kހ��G]eS+���('�{���ε��T���(^(��`a_X6��H��ƽ�y����܁u��A�f0���R���'��~dK2�Ϧ�P��Y��~����R��΂t:���P��iW�"k�N��L������V�6�$&�Md~D��:�?��?lV��8�ukv��FV]$:��'�̧j��Έ�Qg�[��wTXVZ��~�5�?�K��"�5�T�}M���o����
��4�쎤z��H�:1��c���M�bW�T섵���U_�6�o^�^Y=:6��en�R?�[�%�k����O^&��������洐9�,
�^i�.�gȑ�,D�(%��I~�@uP�Q���>�����=/�k
��;"���4�Ny�n2�DHb�e#���qQ�*���kJ�|\&��a�Uh��J��c6��RzV��v|��6r��|��]�V�����o�
`��8�޶� |U{��bM��#K	0N���JBO�p˟8F��+�)����	a��k
�"��8E�(����ǕH���QɎ�o���z�^ov�[���(숳�Z&��'�*x��)5eO����������dn����8��E�`Fܬ��|.�1��+�T�<[r.C��K�L��S�Ыd��Y�*97�V�C>�
w~���W�C����]��&�J��-��_�s&���)�G�{=S'���	v��<�	P}�s��7	}VXڅ���:�o���CH�d�{��p̿*�qe���Z�� �oKe�7�[�t<�G���1H@�5�b��Z2�L�X<�pr!|+}n
��)?�w�U�W�޳�?�S�#gF�{�9��k:���.��>��)U��^f#�q	�e�%qF�[��#�d����4�ݯIA�gc�B<���
kb��%�2��6#��G ��օ9/-@���VvV~i�:d�Eb=1�1<��(I�o��r�xe�r
�U{�+�+��Q��y��[W��'I<`��:�Wh� �h%�I�Y�3�/q��;��	Uڲo����D����e�&��N���Hy���ܶ�W�ZH4���,��T`�`��<�ӼG>�z��㓮*��llT�W[b5�ı"ӻ>F��6r��:f'�&��
�c�1�3��ё�l+S2�\M�d�B� ���_y�;a�78�KG�C`�B!���G���ʥO4�&%T�X"'��A���};OE�zԝN�c�D7�R܄. �B^d��6 `a�)�p��R�A+R~���S���E�=V9�H�t>#���HAu>{;W|?	�����Dz���=S�x�}�K�ث�\#�9?~��É��T��)M��,���&9��	���H ֥��{���aS9o�ˋ�.-[1]ql�y��"ґ��Jl�n����4�뼋YX�Y�K���"��5�
����-ܨW-e`X�L�".�#�f�l�JT$��5'�����g�I����Y(�ř)�'֠R��sSvZ�,'U�����&&��z��љ�%��3�fߐy+�y��J�Ky����(�~[a9X6�-$�葏�U%\��D�	�����1�D�����0u|8���W�q8U��ؼhs�"������ju��R=�"�@E�c�b��sS�4_�b/X|cY,����������6ݴ3ֲ��Q *�Z�`�a�&h�%(kA����!��R-��yP��ސݟ�pd�L���?@�X��l!�K���Z�,���ˣ*��}lu���λ�g�X�4��H�n��f(l����W}��y�/T|�lO�W �Gw<��ɖkH���~k'�`$���7�V7t�]��ؓ�ث��%�+�'V|�e��%oQWI��K,K��Ê���&�Z��+�F��r��W\��%E�(�_�%a���w��+���J��eL,ĳɺ�4��ܵ����W8U�q�?��d E���ެҥ�\��HP���Gb8�ya7V���ïjt��lYꞎaR���x�iUV�!�� �G�Zq[���o�p�2��	���}��L��~DDb����]`.�����������堫��Q�1�i�r ����]ɖ�\#3��A���AK����}`�Xzm�b�;�_�0� ���߽K��p���
����Ro ��V�tF��d�+�A�?��,�y �.t��h��L&�:C �&׸�
������c��_���S.��E���Ũƻ��%�����Fy"<���@"@�TC��->|�ub������p��Th)�� zm���xaMc�����b�뵑2;jʒC���ڄ���8?ک�Be��F�B̊�m����"?�q�	�3��,i�F�5�%>"�G�z�����X;	���QN6X�"QM��H����3���m}O�A�ҨC:9��B�"(�����}��'R��R��v��C�>V��r�����
��9����LS�1�EC�q�DYcyV���w�s�zn�!0@cp�l-M��
�V�tM�X�1���O�9��6U�"��ƞ�!� *����X��s�^�d�#Ǹ`������֕��qG�=�u��-� �M��?���U�|s7u_��Om�B�0����G�+P�nU��%�{N���֍s���
�wΑ-A���,�C�BP���>�u���$�5���<�V"z]p��z��Y���ĳ�4��>���j����g��T	Θ���� ����~yO�8X�:b*��|%;��iS��:aC��C��;���Nu���A�ӻ�.f\(v)-w�$���� ��ƄP�$ܡ^h�~��ۂBۊ7^_`F�EK���CǊ��䣼 #AϾ:���\��ih�)�J��5�H�	楥,�,Ul۸e�>f�?���t9`��,;mm��1;!�&�W�Q�e��~/�E&Dq��*_O�m�����|�C��Ǵv����������C8�ol3&O0�q��0M���v�&�"�}JY�BY��k���]~���ok�G���C7�iZW}d0n��z���k_a����$|A���$7��J<2X���"�����tzDf��8��L0T=P��	%��λ�ۚ������\�~)љ��:@k��'���b�i-���e�We��F��vD�d�hC����Tt��A��ֻi�]�Y0-9�|� p�`"�z�h���N�f��;�erOi��!A�9����;~$�fJM[	�]�:"r��
�������e��қ���8�X������_���F�Yv��5����K=аDS�^�\H(��sC�_��[�>��o5�+��:���v��M(Ǝ��h�+x~�Z�*�9�cV������J`�Ъ�4���:��� ,�e\��ʼv;�NQ2�L�-���b�
�qK��en�W}�˫y$��]�F�	�e6�l}�����$����Z�Z̑G�g�7�; ZG��V��4�OC�i#� 0�_qN��~���F`5��*�W{��{D��Cє�,���r	����G�0.�,������E�H��9�KLdb��b�B�٣�`x��m����H�h��g�p;�ۍ��N�f=�����H�(�I2^kE����X�uʒ�A��7-��'�߀xq��T�͵�G�N��D)[�ьn�.6�I����(�M�]~�a��ӿ+���~;��}@]��090}�����:��P��x�J�9���f�<�P��M�Ur�:��^���&FJuM-��W���PY���5�~Uk(�v5�NSf���^2�q4�Hx"G�q����{5��ͱ�b;�J�L�������[� $OKyyE�:�$� �	�`�o�]yk����	]��a��g�*���&�E�]ڢ�g���-���[���@���G I)�X�{���v �L��!��v�hX"J|�U\*B�~�@���9��Vlټ�8PI��B#Um�|���������Zўp��r<��d_�Az�p�.Q�e�vG�o��y,�G�N��>�n~u���}��d�B�e��;��s5�=M:G�������=Bx(��������3�fEʱ ���3����8�k���N��s��o<����N����Kw����܍5���1�<	Sa��:.}s��:��-z�`��<�䥬͆���&�H�ʩ�=x8.)�q��V��OxV���dG��w0�yd�{�����Ɛ/@2@��
��W�LIb/�&��+�&�T,��[���5��ݠ�����}��k�	�^_�T�_�4{1���t]F�����õ���C@�i��4d�%W�/�5�L
d�O�����y%�������#��t�$Q�;�_@�,Ĕ�֙IF��y$n��H1��Z$r�ω��;��837_��Z^2����:<D��޿��t�K�����,f�)�BHt���%�H�3݇�
{CM�X��1�+آ��م�����8�|ۊ���b4�����@�P�Τ*&��a��x��s�6({e@��-Sg���1#�����c��|�(���p�%U�ۘ5�u�g	�ֲ'��ii>ݣ#���1Ձ�Z���Ύ��4+� H^k�����Ú��R<>لI�mJ8u�_Nkd��n�%W��\�`�̳����ݒ����HMQK"��\e�����|W���la�[�)�!��-�'٩Vg��M��۬\
��:ʨB,�)s�N_:Ә�?�g@֎��-f�zO�p� ���(�m�~F��Ӡ([0���M�u�nT((%�'[��=Jڗ=?�7ūn���9,kb���3ce�y�A@��U �����az��tx���cZX��jK�<���ދ�מ�.�j9��Q�D��z������b��򦢓yZ�}���v�T�(��y�l��C��U׬wx�=�c�I���{I����k�Yhg�93�K���beL��n�3?N)>H+0'�H���h˖����ve�������C]�ɏ���z�~��
=��q���65�7lh��F6����Uy>�����3�x�t��u�'5�`���Ӝu*�t7�$U�t�- ��k(��5�[�!l�p��L���8�OZ�]&e�����nVn�~l�Ӑ��?/�Mz�D��܌Nv�Yh+���>�sն��Ś�8�n�� ��:w}>[Vm%��ы�����G�9��j��m��zФ} ������F3ziy۠Mǌ
��md*���涤V_�,;�{/�3�GltM5�5����?S$���E\<��Xy؜NP=;Zul�.�ϫ�'1�wJ��,Y>ǖ~U�	�o"��V@C�yzz�}��U�Z G;��!,�6~����GPŔZ}T�~�{�'��O���~3V�:�b�o�%<�G|ܨǵ`�jR0,�>W��֊�����6{���q|�>/}�dT�6�J;C������^�� tq�Ϟh�66$R.�桟�k�b�@�IB�k��q3���X(���f��%bAz)\���/��%uC��_�\)rC+���i��@��ʆVDBg�=f������m^��W������h\k���������l����3k�7wf�6�s]�dԩ�C��yv ˂�7z���VF4��s�����7$0������q������=,љ���n1Q<��Y��cS�t$��@P������ۦfQ����]���]��{~��BzA�R�����uX�q��_�2�V�� Z��R|~�IT-��90r.0R� Գ���F��C���j]P��D���M����!�5�l1��܌��s� Lg�x��ċXY�ug�ưd],�#�Z�2zU:$`��x3�V&�%�F�Z�k�,{��މ5:���C=p܇X��l;�j@��-RҘ�af5��0�(q7��ݨ#��V�&��'1���샱�����b
�"W5�d��k�>���Z�>2�/�j�z�Kc��{!�k���5�PJ����z<���R�΃A�TE��Wƌ�⏩ݏ�$��y���Y!g�4�(u�YC>��	ǡ�V���J��`���qsK��|�2Ҳ�ą�+z�r�*�h�!=��J��9���޵�E������)���7�ܻ� B�}?ͳ�/�~�������H)wT숦��Df者���3W���u�r�ҕ����!�z1�@�F�$�.8�d9�f>�_4�G�G���>��x7���l;{�V��;:��<�3�戃�J�s��g�g�Z����[\H�T^^�v��	{ X������}BxTa}�L� ?+lqI�e���7d:��4���O�}����#���h"���1��.�~~�@8�N�CT�;��r�0��)�n�B��*�P�zU"M2� �I֦iv>1[O��+���+�b����_ྉ^z0V�nJ���}�ڋN��C@��<�@���r+҈sFA�D���7����N��N������ٲʘ�!h�fݚE��v	���c݋JV�T�'��(�@�18��9�F����K'-_�R�}���]+�S�À0RCC��K/�4��z C�G�4��߁�CM�y-+(;W� ;�z�ٜ�/e��[������,Ҧa��)P.��� �_=φx���9��Ř!Ѐ�����ϜDh�l��V��G%�t5(<p��˜|���ٴV�`��H��3S�%	�s��N����P��%��-�̧�G�)��t�@+�Ҩe��RD�7�Q�f�j�|(�1�iuQ���[�v��&��U0)k�H2)��a�6�V�Y"��^�"ur��$Ø�	�QDg�wV����&�<D�y/�oa���C���\�]In"�}�K���9�{~2�&� ���a��ᲵXy�1zƯ$I�*)�@��z�&m�7�K�BG�UR��,�O���Q�l��-�D�H��]�i��Q��Y{�Q��AQn���sQ�0�!;D�O#�U�B���JJfq�A��{q�z1]F�M����+V�P\n��Y�[6�o�	��}����#
��s�ըt1��`l��d�g B�B�;��#ޘ�4T��&7�Ʋ�O�&��~��g��­��A��uP��ǹw[�hdx�� �~]�
S�����Z�Ș�8wb�{\L>�����l�t�9Q
)3�]��~w���\��Q4��W%��0�>��1�I�������<��
n&](|�K��@Ҕ��'T+���cd�b���= ��,�x�;���+�c�j��5W�9^���|��ƚ��^����u�2�KY��TT�HBz(8\��#�s�$up��Ad�yk�F'>j@�"ЫX���-�'f�/��9����l���"��? >A�8�)a��_��K[	�x�}.����qԡ_�M�\���Q-0y}��Yc��8��>&ݧ���)��R�\��ŵ�8LN�P�DrX��j���9F�6}ǆ�V8
��(���/C!����֦��M*�]�M�,|�$	v��Bh@$�*�;<K<ɰ��Dsd�l�*qP/�C�%vsTċE!��O`72��gU��S� ��I�RV���!��_��cg��ŕH�rH��Y��z���H속oW������w�����m�Ef�A#�������Nj9ʊ.
�����Z�x������6�Q��v{ؕ����&RH�f�^:{��޵���ϔ�F|dIw�p=��$Ԡ��S��9E@����rSm���
DU�y���;�g`y>`^%�1D�7�v"V����\��g����TH��{t��ź+���C��M����Vn�]7���Gr!i@H�N��,b6TxI�F�c[���H����v �I�	,���np)����B��?��ݦ9�u���Wc�F;�t� ���ߓ��s�K���э����Z�#[��儌��%3hϠ����q��Sm�Y_�����P��p\K`�J�D�"�z7��j
��������_���&Z�!�z�3�%�N3�è���	o�}�pC�K��4np,!�$)�{�����I'�r�	 ��Y�>�Z��m�|m��f�)��2$LT�'�N��nd����ꭐ��d�Z�����Vm��1��t� 7r��:c��D_�l�IpG��^{Z�`}Gs�y��3�S��Ϧ����+�F�*Ѡ<������L��f��W�U�Zn�7�,؅�����l�hsj��fӜ[%���e1��a�s_
ܞ�}}�/��t!�L�b �_�q� Z��I�f�&u���#�?ƯϿ-���4/)��2v�L�2����DS�`|_��ݐ��� I��Tav�'aL�b��3�Q�D�X����W���"o��ir,к�>I�����yːn��rw��W�l��)!�5k���M��+Q���	��2o$#�&�Q,��A7�����.Ə�Y�Fev�u,�������p}�r� j{N�M�������!��)�S�@��Y"Y���14�n��$��=�!�6THs�=�|H�%��A�� h� �L��J�FZT-gxxP?֫��)��#W�E����8�Zd��S��P�h�m��̠`U�Q�V��Np��۪y�`��IƁ��C�2�$1��cn�O��5@�4��u2m8��Kkޥ�Y�����7O�y/y5�h��ȤMP�8Ww5��IG�\_�sZE�
��GvQ	�t}����7LW�[��:)�����g-���>��k=�ӱ��D�2ϢtI=�l!;���Q2��\YI�<�J4'8�k_C�z�a��JpA�z�S�.Π��(�Œ^r�i���b���`�qw�0���D�|�o��� �P즼�� �C������+W�D�.D��I{�E�����uatD`"��X!S�blж�fjK:k )z�anŋ�Z�e�nHOқ8�R���h��_t���%
�86F�*u@XO�J��pa�����͓��v���?�P	��K�"�n�SD]o�d����0x�-ݰ�ޏ��O�ʷZӰ��)wgE�)*P捛����J�${+-_,�y��es$*��SB�³Y`�������Yڈ4v�.�Y�n%!b�D�!7:�;_�l���,fJ5��q2���gv��A�@a�6�w����8c74Q�,#A�ɲ�J��z�Q8����ç�0
���4�y��#�Rj�5�S�,$
��>���_Bx6 �mƛ���v�	�}���ˉ�e:�R` @v����G�bM��r#<&Gq� ֞1��H>\Fv�D�R��SI
Y��롢M��4^�8醮%��qҫ���9�.4�ۀ_�Hz۸'E7Y�+����������sw���ڐRD����o��<1���<�5��/Å��I��S$�0k���7hۨi.#�6���h�G	2B���1�Ca��%
��d���|ѭKȴ*��g�J
�Ez*���J��8ܡ+���)	��23!ūR��lF�	���^�0�� �p��e?ɝк>i?�:7�[~�D���"�,$v�ƴ�C��$����Ǎ�_�Z��-�نQ�U�s'�@&�*��L�I���
/e�nPo`u��ϒ�ҪeKj,h K7��	�V-��	�})d��|2�����A����YA�_�d�@��М�t��p,,��K������9g��į����81� �D�`�XJQ�nd��ۉ�����Ҧ��|�Z�Wl��-�L�n;p�4Ħ��eY�H[(������=�u���0q��-?_��"LFN�ORB��
1iF�����΄��Q���
�3_�M&Z�IъK>��{J��j��H��Sˎ<�:���c�-8Ң�m�Pm��9��Hd)������+ҏ[�%V�q�iZ;Bs�W��u0Ѧi������i�h������gEH���Ԥ�X^#��D���d�Կ�Je���ԯ���htʤ�8�zm�7p7 �~��{��1��� m�޷pi'[/��:�q�>*�����J�gh�0���cፌ�7!nT6C��5��+�|G��6J�e�Y�3`��n��b�l�_��.�tO�>6�@�d�)o�Ua��Y��ꑷܹ�]�k[_eD�5���q�ˤ�A�b`�]��`QP}ǵ�E���y����a'�<��o��(_�9��%�2h��z�v�v�&T'(��P�Aʁ��7�v�	|�@�{]�/��J{Gj�J����u����$7n4Eu�h	��z@�VB޿��ڍwG������'-�%�f�S_���#-��,���۹��8dz[f.w�.>�N:�+e7�1;���b�N&�����3��'��?&�=�Is�1aL��p����b+��w�ё}kr+g�q��
��ݢ�MM@"J����~:�ۀ�,f��m��s$W��Re�׵J�J�K6�u���_����RNL꬙�*�Q���*�F�"��G�c�&�Q�h=��$_�dp�x��`1��7�(��I�� �LkJ�Q�����H�y.�%��.�}���}7���~���y��-�UU/9��X�m(�v 7O:�'z/��O��v�����yEH
ܡG�ߪB��4W&ϴ����-<Rz{D}���S�a�ќ:0�=��JjȄ17+�ijdGJ��_��綸A�%49�� �Q�I��H7�� n_��J1x����"�?A=��ѵv�q,l{5�ݺ����k���!
��)���9$P��6�z�y-�����~�%�9�x��<۲�9�PU���ύm���͍�D(:�}�,��<��[_b�����P&�J���́c�E�]`��[�����*mQ�+�9�3(�þ��+h���0��<4�S�Uv,��T��}�E*�,/	��	�����J��'\�(���=d��ɇO��'�����c�Ә��k��c��?��3F��W�aw0���yB8�t�d����n�Ҏ=���1'>��s��~x���Z&<����j�Hi��Es��j�'���V��?��B�tf�;�K���E#}�k�X֡!�ɇ�� �UG�u4y�PM@�ƹe�h�+�q'P�,����S.b��?���f�w��GQ@lZ��n��49r���0Y ��|fE��������O$� �mO��ؾ������9Y� g�A��GOg��%���YD�g�������$Ljd���r(Z��
�1� G��C�0��%�ͼA�ٯ �����m�%i�9!<��YO�Iݩ�$�[T6�o��˾�4.O��l�wP/��v��+sv�PB/U w�Ȩf�.
"b5*(�/�8��e�s�>�����d��P���H�[}r��-E\���t��&?��x�A��#�_MH�p	X�?8��̅>C���G��8���V/s8Xi���υ�u���7��Y�����_�y�R�WScu��;���z�hXP������f�*_���F���!���xԤD��)�P��>�4���#�v�u��Ն�\���,`~c����D� 4/b ����X���-e{�bW�D<n��d�)s�0`�óO�
�Jƅ�<������+q�"���پ&qAa��"�J+e���kʕF��sQ�H�rb�各���s���6�Yʒswqp涠�&�����2i;U�+�
$�U���Zc���R%�:���f!��_�[���-^���^�:n��dH�揶/�}MX�5���1ˉ�၍��_䖞@DG젛�J������w������U����)�`u���*���9β���Då`~������Fs%�T%����B?a��zX&�	}�#�6��T��H9�ʔJ|D��2i����
'����

ٶ�������o�DM�v+"�ԝ�lY�j����P��e|��F���ʿ�� �5�!u"�N�_1�AM�����ޏ��r&�(7�D�H��'x��T�q㑶+�ß�}���ז $���!#h6�9���x\g�f^�� +% �[z�+�)�JbF���*!��*�y�_oI$���_��u8|re�i^+�:��sE� #�q��S-��r�~�mxZKy�v]\�<�����E'^�Ŭ��5���>E���Ȥ��Z�ձ�̣�=O��a��袹��!Ĵ��/q��9T�L���7GݸL�����ޚh�%ȱ�@A�L$9j��UrB�2��<����gvvM�8Oo���҅�����-_�@�e}�\�DT�pDŲupb~K�'�@W���;3a�rJ�˾�" ���"��j�[�V�����
���}%��99)޹�b�A��(05�L.k��#-��̈^�[���HJ*b΅�D��'�C.�a�\�լ�;�a��IiK8���E1���^�'���:h��\�!��0蒭E��]���aBA�8o\��_�XZj�6h�)/�U�&R��Dy-�E�Sp��Or�>��Li�з�PX�̋�6p�f|Fa1ԋ�!^���(��H&i0'ۨD�@�i���@�^����fCz����Wn/Y��ç�'KeaV���G�EL=�t���m�D�^N خ��WSK	�ά��eN~?�e��x��;�D���i䀯5d�Ei�Jde��`��p���КZ����a��j��y�> HoJ�ì�c�J�������Dp�}��I��r߉�:d�b��{Їx��$���M��L�)5��Ҡ^**�m�{*��g�e��Z汨�p��i9���;�,񼕺�#nۺ򲷬�D�{��}�� U��'k7n��7����� �:����I���n�>*��ӹ���բ#~���`[�����P�3e/�� ,N/��Z�\B�+�Ȓ?:��g��A�Ig!����=����Lcm���f��[��w���[��!�v\������&+m*��o��>��&�b f�zY��l�u��H�I�I���\�f�&�-�~$5�V����9���9hT\u���JL(?���R%|Z��*�?�J����[V�-Ny�e��:j,���p� 	��2a�KxU��r�;E�*�Q�h���������ZO��������Ӵ����fh?e� ã�$q:�	�5���f��v��ՙ��n+P�ѫ	)7�V��
�~`�=X��$�>��¢0I���3�]ڠr��T�y��2�MdbB�Q�
9me���c3b��!b��P����(��V��A7ʐ�u����4���<6���[c��&2i�ڧʌО@g�NIa
�~��߆�mL4�Ɋ���5���F��gϐ_:�Mcw��G�"�0,���B��Y�׬I�ʬ���"i>���2F�bٚvؿ��9��E�q�h�WRa��P�{} N��3�\[Т�� y�0{%wDbuSXeW���� >��%,�*a6�� �����  r�Sf=�x��IX�GYظŬ���2Y?hR�*�n_�2Vd��P�X�MP�x+W ��g�rȥ��eA\���K[l��f�a��~���ʽt~�j�A1 ഈ���m�f#⒯ɖ������'�6�ΛO�W+Z�a6�\�܊*~�ù+��m��Oښ�m��Ҿδ�0w2��|`dD��������������Nԫ7���T�x����j^����/�=�_��%�J��.E]�W��֊������	������Ӳ���>ifEj��}hd�A�����^z�qſ�W�WI����>M��LY��*�o�(܎ќ���K�*f*V.�v \V�֑���3���n��B����>�3��<���ciNEs�5
����z�@	�ȗ]��}�Cm��pqF
c/���[@m��I`��
42k]���{!���5R�@��p��!��%���&��e�w���7 ������/{q�򧸵���>-=��c|1���
�@���Bh[����t&:@'��:����z�.в�G�\@W�i���w<9�9 �OH�ڬ�8y�<���Y�M�!��f�0��P�a���&=��r(HbH�a� �m���.�`qt;P�
ß�L$��c�ϳ��3e�i���k��g,��O����M��L�4��d�� ���nz(�xO�^�^9c��Tu����Nx<�N�9��FX�>��A�/G��=|����S�QVM�ίB�I�۩ΊpY���Z�q�����J�,<�a�2wY�m%�b���Du�����
�V�*-&<i�E����E�C�$�}D :�jn���P���ع����R8	6�T��u�61k��6}���z�2���zL�1�5PTi��I����%`�5s,
�9��BVj���$� �g������XI-C������؃��H�@��+�.�
C}��s����/��i] \.��n�YN�����g����$�R��P�l���L@,�
p���\�����io�ѐ<g�H_���Y��~��Y���F_��+���4��8S��R�)56�$�9*S�ϵ�a
LX����,�lT�*�i�:����$˙�agU�ع"�_�4J�7�/��+������Xq���|W��a]fw��1ZBW�����SE�
Dc̹��wS���������E�~��u�BJ��Ub^WP��`�q���ŮUW����"Sj.]z �����s!k�I��5,v���t-'?�m�H)��H��	*�����a��8�-����f��(�2�-��zYG p�<H�7A�Chn�|	_e����hJ�Gi����k���kFD�/��=��!'�Ǆ�%YVӘzU�j�ॺ�������W&W����_���HI[�*�L����'8�X��=��>2�왻���=�GfY�^<���������</׽k�+�W����t��|����ä5}�*�&��mcm7Q���_�����������X����E�ׄđL�)P��Jj�e$�) Y�";����*�.���mi4'��;���m �CMTfs��D�(��T�g=��]�a����������H��섺�vo�[o <F��A}5�z ���#���H�C �(fG�I�j�']�XtA	z�͘P�� �����f��n��J! ��e���I�+,k��$��8�ش���QT�xw�;��؄�y���j�� (0����)����\����+a�F�Gi,�-�����a:�U]��D�F��/Y��Z#�K�z�j�g�"� a5��{�8����qA�=^��r@�A�!�x �FÏ�+m޼j}|Q�ı�G��
^k�Bt=�E�mSUI�)tdM�p�b��{pT$���/�͆nǙI)�֎�/@�b̬�d����[�R.�����qP��d�N�4��G^"qy�Sl�F�܅�`&���;��~�{��{0��%�ٕ*������7}�;���À�U����IO �6:�! ��w�r�� ù�}o����R��۾��Z�ĺ�_z&��P��y�ߜ�k��f���һ8Vu9�Yu���V%���2h�z*�3>k� �6Ѯ���KCu��Sf����S���羠�T�{�~σ���� �U�y�o���1br���@���;������)1br/>G��h���G)�_-d>�1�/S;���Uko���+u�w���`�T�ܵ�FS��Nz.7K��y؀x�K�ñT�ϕ¢���{/�����_
��>O5�k��h�G�;��h�r_��n��a"1�..>h��Nv�W�X�c�������m�c�e�$Gїb�t[H<lrW�n���LP�T���;5�����N6ez�Y�X6S*��a��m�6#�� ��&��2L�˦�ɜ��&Ie����w�I��3�^;Y; ���X|�8��d�|�akBQN��Ŷ9S#�Cs/v���2�rDy�Ɉ���5�0��O��\_�W�}e�p�x`=�PC�z�$%y�v�������n�/a���5��k,h� 7�7eAy�3�� $a��e��ߞh�=���F�t1K���2=k�x�y=������a�6� �nW�)�e�E�|,D��w�r ��5ž��>wd�Ӏ]_��ӿ~΃�!	�t�yQgo Npdql`���j�X��b%�n�M\���B37�A#�� �Ń���U�||�7ʴܿذ7D�jMg��kR��epi��c�@����	�K�Ma�C)~���(�GH��K�b3|@���Cے|�����T�>�ͬ�tJ�wk�̓�EER��k��S�H��O��5�	�3q#��`2��r]�}|��h݇f#}�f�C(�7�~�ȗ�V����X6�n�K�gR흝��!:�t0�MWq���������"����x�I�Y�	A#V��kks/;�%���&
�GɊ#��ƌ�=��'Q���6y7y��G+4����1�����=�x�S���`�t�Bҥ�W$_�4FK�Er���X0
��Q��d^�+��ې�H�	\����Г},�6���9^�jS'�F�칸]����
F�y�t��'S^�wDbL�CL0��=�;�C)�6����� V8����^�N�k�HJSF��3+�FC���5����Y"im�C����H�Ͻ�wo�8�7����u]_�a�l�+>������*/1��&q~�L0U"J��w��/R1.�*N�}ApB��Oe����C&�;6aÒ�YF��1��f-l�Ŀ���.S,kv8I'nN�f<L��y��%��06��S�Ħ�cؖa��;y�;��\Y�]�G��Q��p1W�Oq��ǐO�ݧ���u��$�`#����ɴ}���6�aD�eо�˚Ū&{�ǅ��%���f����/ �!���>�����,�D��(E�4�\�^�n�I��%� ���"o.ĉ�R�򅱷|�-���Sb��U�g!影:�����+�q�=z�c|�R J��R�s��R�4=Dgm��`��q��t[��M�t&&�nU�+��2Į���a�Ғn�wW�7͚��0��;p$���n�3u_��Ѵf�D��$��)�X������hd������j"q�
i܅I��7�Q���,cs����vx�>������6f�*��$GQ�>��|��o�3�{�Rׯ@��.��C�;��eQg$�%t�~��ß.�55/��a'vRC�Hh^�d ����lof&M��3ș�\�r�ϥ����頡�sq+�R�p&D���[ғ�JK"a����;^fxb`�v�%�[o�v6�Ԑgk�L�a�
��U�IF�Opv�����?������\UH��+���3Pab�	�+�7ELu��/����W*��
m�ak5B�+��	G��+F�h��H�z�A�T�Q�������s�g���%i-7xp��ꏽ�۫҆f��*e�\J�4���"%Me$N�E:�6G�S�^��/,��݄�	��ڄ˷���}���"OM��O:W~͕Z�r�+I�ۭ�*����]H#��-"6�a�g�@!�
8Gت��*���EDc�}dB5Τ�ȁ+}I���n�}��D?�8�D��s2i��h�s�K�Fyzե��ܫ~�k�|wH׺[�S�z�@(�¦��}�.}K1CjR���f���8D�S�<[3�G}f����%�!_(�a�V���;,�_��ץ�����}ߩ�����$�j�}�Ix�'�ܧx\`#�`��R� ꃀw\ /��W"�
sV x{x)N/p"?F�ǚ���&��%Lْb�H��gh�8�6)�2�_^�̄P�Z��5�Q��պ���f��,v�%9���#�\�c�����Ԝ��� N2p�V�<'�]/@���I$��2�@/�*Л�U�:.�A�w�$��C��#PJ�NSZQZ�n��!��N�ڏ�Ś�}Z>ɰ�{,z@�0�L�1��r��~��a٧�����"�b�w���J1����V���\f�\g����u���+I��B��4-�12� c��]� ��Y1�������6W�@+��&��m0ՑM܇(2M�6�m��}!���B��H�D�$Z��5u^�/���g�(38��U�,<w�}�7�&�)��4�̀K-�;�*��"�����nv-2ޙ�C�?8�Ib-��D�<���Z�v��g�E��j��+��IY5��>J�/`a&�Q���`U��.?*_ �o,
�v�Xq3���%l���2x����&��\S �βkS��^�f�kt�?��:��cΧ�G�4�o�T>v����hH\��C#�2t�qX��n��E�$ �l��<�a��@r�Ԩ�P#)�������+3�}��Y���M'[�H��J�L��HD����"��u��s��}~t�+M[g�X��oV/��v�1tl��r�n�n���$涏�+^�u��+��P��B{���Ĩ��(�ݸi얥� � �pj�]��;U\"�K�go�<_�S����&KOS0����������n�ޱ&�Z�����d����A����|�� r0�'ܚ��m�ʂt��:�Ĵ��A&r%��6�{�����	:���;D�ȹM��K� >��|�Г�W�h{\�}Be�Fs�����Qbeb��WC6��La����	��D��:�%�rz��N7sy�O;Fhj~����Qn��%*
�t4�`\�Y����Z1��B�psT�M�8R	�k���V��_���������0���$�э�z7ʮ�4�w��\I���}�P0_��ָn�W������۸����n����F��T2�|�>�j���rs&K��ʫ	8q:xO�M�p���L��;0�rgM�A&��e���G���F��D,��%�ن�p
@I�.E��}���K�bX~�K�����B��ս��$xF�M�j?�*��M��2j����H	vlm�%�����=�J�A��Ej�ޓZ���OV���kI�W�N�H&�����Xs彷2e><G=j��ק���.�S�������+^�ؚ��Q���i���
 �BH��=L�\)�ٚ���0��q؅�HM2]��r���rYJZ�L�17���e� ��d�`W6G><=���C5릸����|jb��K��y��Y�p��2d����DV�����.�t�Й����d2���h"ۖ��qk�Ĭ�Ng���	7؀���V���owN�|���x�lU&Gm�"�^�xR��թ�S~�~��CYH�ܣ�G�d�R�Lc����~�(�Js��`�l��<}&<XZ`&�(�V~�pk��Ɗq���n*���$�NSeň�ޖD��8��`P�<����^�O}��*;�T�ê^~�#��~�CO>����u�������b����E�ߺ\HQ4���0&N�e�<���nj������R�c���9	�n�`�fNE��.����x[���4;���)ȑ�1.jK�����nғ�=�����v`��W�?/3�H��#G��;�Y����94���^��5�J}7�U��@�Шv�w$.d�I��j�3~2;R�i@�*7�憍������>��A�G�\0<��K�����=��=0[%�̾
�k���s�I��r��_AҺT⿯�[�j�pZ�Gxh"�ڻ6��yZzj�jPe�L�OC�o�dp%��.l�C���u|CA&�����uV�P&����,�UȰ&�Ǔ�a�K��5���=$"�B�G	�<a�@��`u��(�����t|���B]���U�k�)3���c��!祕���p�j���m��"ެHp)��'�o�00�w��ϴb��C݋�#j��a�2 %�Mo��͉�
(;���,��QD���=�Sq��ؘ��u��*�ӂΪAZ��vL��a\}�*~±�q���eA����(��b�A<�Ƴ�6J��Y�B�-b���X���	���5�E�G<!���H�g�^�U��K!ݭ}`�*��F�d�wc���8*G�æ�ͦE��;�����s�`<9D�R��зhuQ0Ţ��&� �)�&yR��8]�������7q��IP�]��]m'w8�ȲQ��=R�@���uhԄ��{n�p� iJ�g1e*&�?#��B+7|&��Β{�"`X�'g�uc��Q��8�M�t�k�U����c��Yqeq/§�~t���������	��8ԫ��4R	1��x8�����*MB��Q^��[�fe.��(�TA#��CZ����TSc��� FR1f��{?�sc���Yȗ�����&
��M{����>�'E&�ʯ��J��/�7�([��܅��'�H'5#-�(�-#�xY�9*�t��N{X	:�k�� Tq���r�D}����wvO���8�1�Ȏ���˕��X��+xB-1;�m����$i8/��#�!�4��V�5�[��(���&@�v1ف����k4^���V0-y���}5����jnTF���ȧ��?�1&�c�����B���@vs?����)�o���d����=V�1��3?l����#%����S���1x��{9Ռ�xɘ�V�5�U*��+|[����NU����x$��[�Z颺b0�E��}�t�A���\����۱R�*�/������9��eW�,��`��J��۳��^�O�&�h���twPC�$���@�He\�*rJ	|��h�z%��^(��B��l5�����c��c;�'�"7,�G�I�^����g�\\��\�%{ Ýɕ�,��Yq��K={���1��1D!��nN��t��6v�_�,�G��<�ta���b6��;^�y;�?��kz0H��X{�h&I�%���W�6b�po;Y�P�\J^�}_�J��32W)XrP,�O���_iGh���Ш�=1�R:3�l��t}�^�V�[8�؀���֘�{��K ����q:A��fk��`�s�������w�-xQ�+��_�[,�l/�0��%Pv̯p����ť���Cd�U[~ۄ��Y���9)��#�(��E<�gX��*�HͿt�^�����i���2q��ѫS���]�K����d8-�m"S����;>%e��5�T̚��͉���U���t�=+h��cJw�^uN�?)��<�lPY��Հ?L&� v`J��7y���}*�B��Q��N�"��.&E⟿�9�n��e�'�q�㉶ 2�9�������W�ΔО�y�v�S�w�	�7Y` ����%?���j5ql2,����0��j;��{1��q��l����z�|Dw�z��d�#]�6b�+�P�:ĲRɜ�-�ݯ��q*SU��z�����~�m|ςf~g����	��6a#������/X'��C��]�7F�5m��]����Oj�p�M���~�[oUؚ���ɂ�}�$��nB������!93HoY� {�K��cG��F;�X7����~�����Qل��BP�_�|�8�h̜R˒�1Ƅ����0��	t��s�Z�բ��|�|�����!��@�<ްb8���b����W����:�f:��p_/���c<�_}�8%�|��N7�pKg��3-'p ���5�r������X*�s���gkN�ViW8�n���5a�-:��U{bs��Wz��m ����[�m��)~�Sz�8��j-�xa����ԞL�ͥ��D�Z	�iPPWo>���`�\g��a�9BI>+5���:.���E�7 ��-�q�҆[h�2�x�~Q�$�}�<��I�x���<,�sL��'��_��_˝��>�j8ʵk���8��;<W����V��)����F&x%��}�L�{�K��~t���20�PO����� TK���tي�����7}�p�B������9���i)�N�i��6Vt�
b)�y�����x�錀�}��g=�,�н�kbҴ靕rjxe���>39����T(��T��PC^Fu�*(�9�6����>a���]fN[%�Z��,e!��8��ݐ�N�`��T$���a���x��V�M$��!V2p�]/k�6����]�mvU�k�b�q߸�����o����MY�7k�^+cu����W'c�Qv�P Է�N�r?����N��[�������Z;�
���w_2���a���ׅ���$8�議L=%��T
��G���8:�4��Hޙd���'l;�R)�U2g��P�/��w>98Ub<78���I��݆Z�S�_Œ����z�bW��Ћ��c8����ў�����z뤪?����Oz�3�wVN�����i_��П,�*"qo�sK�����R�:o&�X�D��l�U0Ŀ�q���|k|��g#.ؓ��}oV*��b�*�P"�?�dޛ�&4�Iۆ6��T�D濴�_�=�(6��e�@*5t4-�1&��[�Z'Y�-�<���[�����x�A�Ja="v)u���	�( Ǔ�vP�Lq�(@Z�)�m6c��T����"����,k�����.�x��'i��rִ�vv���cN�[C`��B,��
�]�c�������=f���m�eK�{.�0����%�ְ�_ӝz��U��Y4P|%F��P6ɪ��T�z9��������Hp=�h�������Kn�}
e�Y��d��칗�pv�0!Z���:E2�,][�ur�&<�.%��+A���'N8@�j��Sq���Y.��}���|��#�ԙI��z�ā��8�rl���ᡌ�����f������ק�Ad�c���ƿ��(�fTꝇ{����^�t����yM����]��M@Ӛ"�hi�NR��N �0�2��)�7�`��K��>�3�.��S����Lӧ����X.W�vX6l�&���XW�X��r���,�2�D��&JS��7j
�7�]��Y,��
u���	�p+�f��� ��g�$L�Rѫ�4�.�(�g��h�g�O�K�)�^߿�Āc,25S��9�zn)���ja��?3/�d:%5��!�O����f��J�!�nJm��J��-Ѯ���x�j`����FU}� �0$~ܐ�AI��*Ee*�\��"`[0�<~��M�R搢���.mo>�4�E�d���zv#t���\ ��ϫ���(��""��u�K�{�t���`7}* ��-W��/<�5$/�_oQ��"��#4~��&����(6�Pzс�X��?�S�#V� �<�2� �����+�sq�^�+��I�5�fY�8��n�� �3w�����1��I;��Q�v9v;@�uEE�O�ԏ�P��mK(���{���*uR`�q�nX�����t�,�2����+E�3zq���$ּ���&էGh��ul�x�B.�В�!��I�@�@D�R/G�Ȃs�X�[?vB���?[���&b
�Ej̚��VLH�	�������c��H���W���6�.$�y;�;>�����&�׌���=���d��
,���ZqJݘ�=��Ik2G�6<	�Į��X�۱��L����@E~�'
r8�V�����欷1��$�����g�`d��G�����2�@�_��?4�\IF �ٴ1̐gi8����NRP'픭��JLp]a�'��}J���3Zۧ����8>8n>�S�c���/ z�薸_�;�E�~�]bh`�w\�����G�vg��>�ǂ�|��A6_}Y��h�H���ά�6�?���bj�㼗G�)�2bD0�*�	I���Q^YU�R[qYi�"�`��a��\�	�mq7.^ >EŁWt�`�G�P�	�[ �4)��1�ޭW|p�	�Q ���/��$m㜂�U�j��|N�H1{Cz\�S���9��b7 �ȼe��N�z.
�t����L����j!g��g5W�C��v��ܨА˴i�A�!���X^�Q��N������6���g ��D6R��7պ��С�N^�[�I����NG�A�Af@��B R,�G��l��/�zm�cJ��w��G��������ګ���L�5�!�'w&�G�<��i��_h!�`3��^+��������M^�ڀ���v���9�6rK;�bo��0�)b�Ƅ��s.��\Q��N�� �l�������;�.g1�K�?���F5i��ْ}v�˟P�I�^�.������m��6�7߅g��0�,z{��S(kn�z��@�M����h����Z���D8;Em#ɀL����S�mv< �a1�v����dh.?���ȃ_�v{Ź�(ƒdT��u�?����as�*]�>)�;"{�y(���{�=NPe�lTɟmK
�oA�c�ߚԒ�r=�/��܏=d闊��|����=� >�J�RǮ��v���R�+�RK�@9t�ZɎ�C *�e\����k;ݰ�̭���� ~�v>�N�QH5��բ�ψu��@=O�6|��gK�i�"K���)�2�H�~09�w�����6Ó�Kݒ�x|)6asL{��C�P*m��"�*IB�~2F5�<�,��(ԉ��p��x�4��6#8�aWq9 A��� �ɜ�-:o��/*����˼T_NN�%̀*�'"d]T��L5M�a\2<�J"!0@��m`�w�s��;���P��h�_�ח����YP%w���iUn�bk�g��|:(�]6I�$�5�Y�-@ ����+kر����[�\�a`wfu�a"BB�@]i�X��;9�Ȑa�6��+w�ݘ�Rp]���*��˖�ʽ��!||Q�Jy�K�Ӯ+���
�|��M=���ѯ)u�R��Cr:PGga���ó~��y���I�� �[�@��$���Ow懞A�AaW;�$��g�{�m�"�B���^N{�����fq�#�"!�/�U�nZ����C/����ɪrX{�6˲�`��ld.�~9D�<��c����Z%_mj{^�||��[թJ�u����/5DG��P��ÆWBvz��fMrL�h� _q�;����[�\8���lr?��Ej�ǃOR��[P���������A'cV�~ι]gO��G����2�NԠ���k5{���"7P�ScwR��@�L �%��]z�o4k�j�]2k̗sεrq慾�J�8���3]���C�~�^�ڗYmj���\	 �o��5a�y��y��-M��<��)e&N6��{�!H;�v~Ҭ����H��"��of�( Y:R<Z�;���w<G��[��4��K��lTv��q���\���55�@<?\��������ˍ@�3��wꕬ]<���\Kei�G�^������x�V�N̆���x텫� dD,ˢ�x��ӑT�k;D���p�~�!�޴]���$*��G1�ٌ6�&{�Oɶ}�j���9tU��. dP"�#��C8�bB�,C���S���|���C��"���d�hyߌ��IS:)�������/�Z�Y���m%R8
H�L��$6�u����1}��a��Dkne�&𼮦d/���B[�Ӹak�hmH?�i ���~C0�F�X�C6A	����T��%�۹�u���b@
��\�~���h9eC6�����qY�j���� 5
�V���{@�&*NR��wD�P&�֡c���� �e<\L�+k�*k���>�Y��Zu�
]^�	2�K`ha�Fb�,YUI��X�C`-�Т���eUי�H��G��N�ZJ�����-�A�9lfwk��� Nb�B���P���)}C�,��I�&�د��l�, |�qP�rt�g� ���&6�q�߂��K��.K@�rʪ����:L4{�V���"��n����wR7�t��0��_,����S�}.��u� ����Q��=P"�<\�!S&�����w0!I}O�����u��Lٽ�����\Z< ����~�/y�F}����:C����n�.^ ��g@�}V6�/���c���)��,	^�N�1��|c.�8���jמ���?�p�Y.����h����O_�j�8Sg��0ޤ����mU���ݫB��10s?�!�i\>������O����|!�9VFy0EԼ��w�,\�PL�����J�a>&8��*gq�O������q
#x����Ci�����Eݪ�|8�]l��@$U���G �wW7�P�=������رw�H��r�12�Ά�-;-���b���pR�}x�"Kg!���	'�T6MĊ!�pU��w%%�9��C��>�/j���Y
'(U�)qq�har`��Y�3��宬dT �[Қ�}פecuQ��X������>?&K��'p�/�_-�o8H u��Z�(Mp1G��xK95��L��(��U������G�~�y&L��y�����)8{�w$�古ҵZ�����6�)C�`FHR�xn|����"I%Cc�.LE�n�d1�L���� t,4��7�2���P�n�Y���>�(��Ym���YR,>,:�aN�N8�����2�;�ng�I ����S�H��^���:Vd��p ��t��u]���#r͹����9�^#�� �TIE��!�ײ�36~8���>HC��;B�����o�����_��k-�\��nO�^�||���N�:L�q��	�B.tVW�HH�r�F�ⵖ�"ʍ��o��.n��^�#S��X��$7�-<,57��E�Ł/�3Rŕ�#z��+� Ɏ�e]~*���J�Ҋ�(�e�',����&wF�*A`(��
�'����Qx�-��H�I?[ۼ�o>�~��$6,=R����O�Kc��*��v^s,������fD��N>����=o�G�;�@�3.&2���'<�T���H*Y�E�KyN{�/�r]b^���; H��Zv�fT���3��?���h�f��z?�}��Zd��0d�ĥz����^��,��)��5"��b>���9Ŕ����\�����2���6|������l�M{���\˭�AH���@�HP�����2zi%�](��F�/��C@�!>�LY1��{���!q�)�u1�Z���@��4v�)ݰB��p�&#K
��%k�����JJ��M�T�8or��Q��g\����vI\�$T e2��ჵ���\sĜTb���P=�}T��宊���6�x�*aZ
?]7Dʻ�"NX9>j7�>'����;��#��?o붍ol��{ۙ�0,�o.p���{���f=�#y̙&3�b�c�J�� ��ٰQ;� r�J��x.h�1"V���@�}�!�7�Zgy�*�|*9�)�e�^u,f�靘�d�W�h����S��(�Ӵpj�ܖ�Y�(�g�x_ǐ#�Hc���iOڷl�s �E$V�~��t�T�]�cR������Q�W�JΖT��y�\���G@f�/#��D���C�$j�8�j;'�4'h�7n�Q�r,,�-��D��G2��/���k_�a%kh�K���T$ҒpW1�L.��:�f3�X`�ҤM���|���T��5~I"�����G�'�݈f߫��N�<�^;���e+L�_�})�V$�*J�]![v����}�@�� �a��~�F�뫬+������0��u�7p6���!��ӂ$�n�S\W,@'Qj.�����lW��IP�d'�v(Q���TVG��R�E�`��P~�]^��S�C �����}G�D�v�!���R�A�l�K�������l���3����^x�D^���tC�6��D���|p[p?�{��cz�L@��+�<����ݧ�ŧm��N������P>�5+ީf10P[Zpyx~j?~��4¬MN|��jˌ��3jH9�~*͕��)��\�쯿�h�у�O�i( yN/�O���%ĉ��&���06�h����`�{Mzp�#���I}"��}0È�$i��}Q�.Gb�e�\�^ ��P�r���Xň�`�2	(�]��&��D��y&��`���n�嫂�G4H��hyV���yGR�G�b�n�����w 84�n2���qw�g`�� ���d/��7�#^,)�N�cU�FB2�(=i���7x�M�;J�J(���O�1��^T��l-W���U�ƻ�<Eo]h:HQ��Φ�/T��/�`�z|-���	I��j"ۓC�&n+-D�h�s�*c��rK"[���:9�ڂtS����Nڹ���5�)TP���F���lZcަoSO�|��n�vcj2�A1���9���>�� ]b]�!�T��r�> *VD�.��ӑ�O�j���y�@�PT�`��� �mon5���,<7`��zEG�?O�ѯ�V�o3y��xط_�Z�1��EH� ��K�5VH`z�z��cS��3�)��$ ���i;�;ґI��IZ`V/=���W`Ha���1>�ց_���.)_c��
`�v���껛pj�N��|�-ߜ��Y��_���޸�d�g�>b�%{
	�{����W*Y���B_���R�վ��S�3SR����h�բ�Q.
<F�;�����]�U<�*��<�v��a��$�N��F���tI�����!K�G��B��S"(�O�8lP,�M��eb��B$�P�F���ekI��j�餍t��4�(���+O=�!c�Sg�B&n6�\�Aw��&��J�`��B��⃲��Ѻ�JyB�2Z��ŝ=.>�e�S�r~ߝt�C��&�wCJ����x*��ۖ�^���/t�F,��︷Ħ;�11���pgǰ���+��Q���!&��f��_ȱ9<4]����� �d���{&�pom�W��&�G���@��é�I�f��"e�L����7�]�j�έ,bKs^e�ڂ>������H�I� �XR"����#�z�G%�4^�4W˪��g7C<��L���q�z���[�7����	c�����G�ȿ�iSJ�q�S�" ieQQ�Y�h'oڀpl)Zo<��^����Y�����ߋ�5y��nj�����@����~GU<�~�B�Ը����_�ř	�$sinu���z��f2��q�+n��U�9�����ֲL�W�̞�UF�5#��:)[~#y�����iCA_5�����u��#{��`�A���u�EK��'|��5eb:Cw?G�^��r��,`%��w�l��( ��-������"/"\���H�x�Ee8nY�9�X��=��"&K6�w.r���;�.���y��!�x�A.���I�%I�wuɢ� ]ف$�F��J	?�e�*>䜜S3ǘ�H�:f4�����rʙ��9B#t���@d�͌�����`�E�����!���,�9�}�%���}�M�^���¶bjj�t|�cCB<PF�=����F� �ok�I.��H���7�X�.�qE�!�d��wmז���%5@�ݑ��H�2��5�L ��ܽU�85Dޠψ�z���w���A<�����.h���1�e~�E:���NP�N�|����*�`Йdk���}�� .�UIRw��
��Db��0m^cI�4�4ĩ���r�]��^ŏ��Y:B�T*����v�g\k
:���d�e�[���,����Z�D�
�$!r/q�X��WkR��R������"�?��P��c���5�y6w̓�����MX
DJN����\�����\���ʏ�G�ce�3S|�L����Δ0�����eV�MIz��M�L���"�6�J~�,N"�G�ROZ��ȿ�P�F�0w�7꽣u.��A4c�[��)Ʒ߯e�I�h�:��ੰٜ�feN�qL	�NGΟDf.�I�o�����fx�o�G*kL�uN�����p�]?�QFw<q<coC.1�@QW�o�O���8��.Z�%
i�jH���,�q�'f�g�FԌb�,Ta�Eu�=s�o	a��'�1$f�����n��Έ+�,MJ�8�/{�pTYcZ��=�*��VX2�+�A��(��;��[�"�s�Q7>�Y�v�x����TzIF
�š(��5-�_��H(ZhKH/`0�}s���>�4G�NEj���i�=����,�#*��n��_�W_%���xd���>X�		����HT�����%��H�9�,)�"���*��j� ��=(t�aCIʙ7�����e#�R��$E��wa��'��+�<��_��)���A
�-z��(�����s*��!LAܹ��g_����f�c�(>� Z���2��췀r9�3������bHS�����L�p��j_�0;/c�B�[K�
4��F�����?u��(�����]^�H��L��̱�W�9���gП���3��r�\넄�����X��"8�`t���-2Ljs���ixP��p���y����t���`I�Z�qc.N���6_
��ۛ:��bO��� �`�D��~$��ͼ�]9�yM)�^��G���q�������r���W{�\j�H�C�'2��B�m[��J�mG� :�NPDNQ��r��wR���D�1�ۍ�D�ev>��e�z�?��a���U�ŘdN��-ǿ�Ed�&S�
����⵼�1|��)e�P�h]�.(���D��}��؇DjH#�M�U1�T2��*�T�0�V���:�A�7�����a:����ء�&�G΍"�~a�/"��:*��5q��h%f4�*	��]� txVА*���mP�����1C5E�wG˙�d���:��b���1m&�Fm<��d��H��$�$ �tr.ė؟��TU���/>/:�<.��Z��`h�R�b�z���q������	�5`蜢Y�6�tPM|[�q������(��t��(�<��ޜC?h���ˡ�fq?g�B�u�m�p߻O+G����u.�X<�[�¨�E7k{�$[�yruc��=9;X#o�F��!;���?*!�~[/���CܲEZB�v-�ovy_�4�v�[m^�����%,M��쏒ĈV�pjʐ�N-�L��*Z�������@�Qc'K=���k��*�z�Z��W���w9�[	��A:Y�r����>�����5�)���w>�nlDݪ�f�-�H(*h���s�F��y�H�� �>,tk�h�i�J�]j�N ֗��{��$�	���;�{����&�+�]�5PE{��+k�*UG�`"؅��~+����_�#z�i��:3l�2���U�Q7����V����2`�D��u�H��|�`t��f����t�� gBD��1��U�̐���&8�0׏�iݠ�S�P����x��G�kR%:b���I��W4!۠�%�S$6-���A),߂c��V!- ���/��u1�1�T�p�l*�E��v�I�jN�R�>�|��-&��;y�I��������$ �tP]�2��η;y� &Z(B�̪�Z�wEJj ����+�TF,:��Tε��$�BPVa.���}���ai Y����=�#���y�)֯ q�l�@m����w�{����Z�'�T�j��љH�oQ<PS�דw�߲�V���9vL��9X��r���K�T���|4�Ihx�W���ZX�@"!�sر�w+��9�5���?�d��Z̚�VR\�U��h��iaTA:�au�%#��Y�,�OLY�S�	*YS�^�4s��h��U� ������𸐅��tp�ޟTր2� 9{㾿�� u`��WpE0�:�8�7T��?Of�PTfT2B%����c4C�M�QE��:�z%0����ղ��vK����� ���4MO�ۈt�-6����'��x�����	ԏ���>����뻰��u��'W�Wc�LZ�{�r�CL���P�k�+r��VYߦ��}�^+BWt�>�ŵ|�5v�U`�6V�U�L;��U���S4��+���ћ��i�܁��FW�+�i�3&��yd�k�$�Ŋ&{�%b�����4/�n�,dfj}`ȿ$d���9����o� �gc��1���YI�.�AdC�\�{�C��Be���r3�2���]Y�]����x�%��E.�@��i��!�ث�y��O-H��<��uϭ���ܣv�R�ǻ�%jႍg��{��G�K)�0��8���p�&Ya�6�>~4P��d�yG����wVM�C�L�@(O/���Bg<5x�p�k4+���D*�{^7���L<X�&��k1���3-v��M�/ʵe�yܪsS�-�N���"�"j�A�k�/���9��P��&��d���J���=kZ�]C�H-\m�fM _S��BM�)�Hh��&4��Q�z�riyS&��r<>�/sT�����36�<vFll?@*�ا��~�t��p�5;�O�D��T�c�Zm�0��Q^�p5�������XB(h�����..��G���Y/N�n�AeL@��.A�ʹ���^t�Qʆ���)p�1�	K��<���{^9��3B�ZRG�S�d�Bnqإ�嫦��A��?���\kʻ%{�'���L��7+�����3]E�~��8x�"K!����k7�-W��Z�i���b�*QI��v�zz�
:�0ͩ37=���Ky�z��O�#Ӈ1y�Ԉ7l�@ M:`'�B"����6l�p1��H������y�a�v$P��׏�D���"�@l�KL��4�ܠ3�?E������
�F����̪�FuQ�o1���7�N����7Ė ��I��27�@�Y{	���]�7]�먽��]]�� OF�������ó0X�P�F���0�-$C����F��6zP�!.��1�::@�>{*�� b�w��2�~��r��v��3D�3��P�W�嬅�ự��M���y�h�v�NE}�k��V;�I�����0�
ma�lw�!,���S���j������h5��^�+�}5�����ٖ	P"P�L�j(���$m�@�J1%�:�ҷ ɏK�<�e ��{��4V��ם)�MO�r�2}��J�t���`�]$Ćs�k�<��?-[�:$��(H���m�>�ą] ��
��`�wJ����U���aZVo�24��\y�W�OO ��$�������=s���t���4�׍�T�8g<q����bY�__G����'\�y��D�,i���v|ҁP$��[�uȜ	���"X4q �����O�#Td���H��������@��Z�� �F�H�c[gJD�>=:I_��\�?�����vj"y"MU�ƂI�iW�1I��z��i����x��~�>Q��N:�]�*����p�/X�W�h��D*WRl�zl�w=2c���Z�[�c�P��jq���8]�fU�+2��¨l��0�����i�o*@������s��$ݛQEEm����D.olS�U�a%��H/� W�|�Y(C�v"�pr�9�j��g��{�S�oj[p��,���L���	V���+�Fʕ{Q�H�/��4%���8�匢j���UY�R0u)��ۧ�fڈ� ���P��?�n�[�t'��DK/�����Q�/>�Q{�	p�nߡ���% �w2��N�>_a�O��7�Qn�@�!�#42�����KLx6/�+�gx[f4��/X;6S�ֈzA=�%���c�[�����[4C��B��B��s��u�Bg�@|SG��VeA�hņ2k�M+N!`�-�9��V �r@4�(y?��vZ�B8�}}N�`f�ezc�h��j���t���b<q����8�yl���C@;=��I�W���7����1�T���W� �Tϳ[J���W֟���[�%���l��Ҙ��@챘i��������=>t�.���^U����@��~]��J�@e(ڱ���M���u�53v ��85|�I����l<����N���)�ʲG�<�����EN>�
e�]L������ʇP�8 )ӚZ��0�4� ��ґ|�}Ȁe��<'��"Â���j����r4��yrv�׃�����n�sހ���r�TF���;������7��v$eLk���o�IΊz_����(B�׌���Ƌ4���ڼw:�NW�	�3×/X\��g�9&nP�*�U�M�����JjH[s��Ǔ������k��{g�,�{*t��q0��q2ȫw�Ua��d��g�@;����O��� D8�".�(��M�/���3�.#:�]u\���f�W3!���G�0�ڝ^�7F�h�0���D;�@/�d�[.�e��P!��5� I�R�E��]�L����;/u��F��oi��%���r�I��aJ���.�����g�9�����)�B��Ɍ1>���Mg"��R
����3~�%��[i��?$y�
 �.҃��8!P5	$�Vȑ+�o�P����������1���e6���s�h��ύ�ʱ��{�m�r5�L�ĕ�P�?󜦷����	��s����0���AԒY��\��>��h�B��W6]p	,}���k.�p�bZ���r�/�����W����ds�EZ��\L{{��`�^���6���Q���5��Λ\s`ݝŠ��S�*�����e�2��G�*MR�/�xxe�_ޖc���dz ϡ���ZlsnQwU2��?�o�U(T#�Q�(��4ߕ��,b}�v5�ϖ?}�v����m�E#j�
���lVAW[O��Ia�����`N�/\����=c�0�x���i^^ �z�ǒ��UcDS�,�q�ח��e@M`���v�%�>0����Y89��s/)��$�#�7ٰʴ�4�=��m��;��墙F<�8}x�\�o\�+��K?V����x�G�Y�:�9��|��]C��6T>�Ĝ,�F������B�
��+a��&�ese�N2}=�:�&xGDnU^f�����9�p�[K�䯱�[k��bT~��*=7+�~�sff!�X�C]�O�AT���V���i@��^]�)���¡���?������Ba�o�wXĖ�1}�bfg�#x EQϿ*��i�{cg%� 2)�X��`��#����N6�늰+��*v�"\���:�h�uO3�&��ԝ� X(E�b���څ�;�`�Y7/ ?��lg������/KW les~I��-
�(���8ED�P�qqRr{�;mC�t�?���q�盭Y�2�j�"�#|u�*����?2~�D�W���� ���Ɠ88�S;�5����$6����ĭ�qq�%x��M�։�c�$�iYN��t�\i9n�>����a5)j6�%���T�i���w�<1Ù��Wm������u�Ԗګ�;��1,K(K�2r�}��z
rM6_� ����;c|F���{n�PY�e���;%��~۝>[�T���
E)�\9���r�����~��	C�^TG�$Bj�e�z�ɷ5�v���Q7�B1���&�`�Y�p*ڡ,���f�
��1$L��s��wBH� �T�A�db�ҥ=��c���3A�
J�	���l��꡶��8Fۋ��h	���*��n�q��=Y튺��}���������.�Bl����X����U*��-��هtZ�Ƀ�Q�{F��rͶp��`1�ҍ���I��+vG6g>';��]&r����:bpV��Lدٺ���,����e�R'��V͘�̇��w^����Qf��ek��:��y#�m:����* ��]8|A��p!S���y��\܋�=�t��u�"�d&�4�z����"�q�u�WC�t>��q��^p�k�\4Y�I�{O��-ʹѿԙ���
��+���.�=8�H������$Կ12ؙm���/��Ģs$�F/���~����[��?���	p�'��..�ͮi���ݍg"�F�->��E����=kyOc�c$���x3x��`F�!g�Z|P>��Db?��f���s��L�.g�oY�cE|Z&���T�h�p1��Ң�B�E~C2_���.���9��;��q-o���R5�Z�l�.��J�:�Iv��Ѝ��G��?d�K�;O)��a�횀Q*�nQg���C##Z��ᣒZ�ӌYa'���E�%k{1�	�I��?�Uac����b^�S�����+͍�5��ߤ3�^3�Rܛ��3R���͉�2љ���5�4��D�R=���1��0%�}��&���02���c��?Kk.xr�j06kzH�u$�RW	eL$I)�_�����	�<VS�-������_dw�^Ơ�?\5Z�-ƣ�:����H�"ӑ�w�e��֣�H��.���ϝ9��z:㞖�ń؎�0%4�<����X��-A�!/1�T5E�;�S��`�ƛ&�x�^����dI�^����<�3��~�Sa�;UKѭ��)y������;�I�N`��#�.:#�����D�]��M�q}���-!�|9���1tz�XPL��wR����˸j>�3��wk�]�m
=��S�kV8gX2���<Y��/7}}�K?͙Ŗ�ӻ��r�c���Z�:v��_�Q��8Nh*�(�����Z}�F�2X��"N�@R�5E�WUG 9$J@���\*�}-Y��iR�k�Bv�9�b!��ڦ���E������ܓ��N�R:�(NR��/Nw�Z��喒�w�t�H��y�ׯ,�R��(9�ضЧ�6wv{��f�����u� �^#Z9��������=�AmZ����6hO�X�V��^>-���4�'G?�BR��{1����G$��laܩ�(P��$;?���ā�F�`�Jy��;ٍ�hG�Kf	��-��-������/}����4�2�f�+���%��i�tԌ�l��OB�X�`b�X�4,�r>�7r"����`�rT�$PR��7�Z71��IR�:�U�e����N��ゎsY����1-X>ҁ� Y��}v��/���z�%���q�ra���r�:b#�C�Q`�]u�OI(��FH}��/��--q�sV��U7.�������g�����֜��Е�}ɋ�3��=���S.�� \
�)�����ȉLfW�nۀ"��y�3w���\\�����c�b*c���#�i>ًxU� 뒮�u@���������������U��J���/����{^��B'�̀���,�R1��G���<#{�=��N$�$��	@�d+4TK����}�҇��W&t*+SG�z��'Z)L�bb�z��y���:�1�nPnc49���\N���]Y"�u��֒��{
�������G�%�Ɔ�֏���Sm[ >b�}[o��Ϣ5fqB*#��t�\Q{���҄��8ҝbڔֽJ�_�h 	8��>�1�����^����Z ����z���qC֑w%,�?���W}�Qt4}�>�\$�����=��;y���!~��J7��(`Ѿ�u<���]x��F2��!�@��mano�:.w쓒�	��1��t���!�"�.����u����CB���K��G��-�tPD�qڹ�]U���dU��
����I�sΒ�6��Z��^��]a�fJ� �}�l�4|������T��
��z쁊��8"��W�L�qg	�.g�M��&�_����CG�H�S��~r��dL�X	&�'	�^��jE�
��.��q}��/L.q��CV�_�Go��XW����<6WB7{����8j��C�v�[�/�����<RF"T>N�|,O_���dȒef��;��K$[�^�N��@b����h�;ϥ�F8��">����Sٮ��� "�/wl�TI�u��	P�Z���M?���b�F�A�{�I�u�U�ۻ"&���:�V|����3xg�]��agϦ8�i�;go/��l��E�$@ ����iy~[�T�>D�K��+�X�Y�G��1�Ѡ����:�}��+)�F���a�|V�5zw���<k��"�㢧G���X�AC;SͶ���P�Ur\����O�q�t&d�t/ś�����;�U�9x� |�}տz�/pyƟ3�]]JZ�e��W�IYei,���_���+�b_}i�d���o��"
�:~��y�I�{,�����{�CY����PxOm�_��ʯ�/�F �y^⪍xA��3L/��*�Ixʁ�Ib�����>7���~�u���s ���i�4�/3��v�*sU<B!���4���S�o�>vs��h&BIy�>���
KI����Y�o���?�T����Bv�@;Ã:������3���H-��L�C)˶�8{e��$#���04��j0⦶��dF?�j~��Q}�U�i8dʐ|3�,�f�N�nf(=��j�ݬ���8�t!t��@GP۠��.������������Y�om�7=�r<8�r��iBǵ[dݚ��9��&�Ro)�r����u�suk"#[=����c��JF�V[<.�H�P'���+B��N���0*���Ģ�`>�~��h�B�1p�}��^t�]�F�}���5���Q-�|�	��=z���;���Z�^�5�^��@�^��S���3#DK=+����Y��*�h�B8I�����Ov�:��N�G�T������8����m}Rئ�G\���T��|'��X���S��.��F�����D#ݪ�Z^�����$�J9��k�zI�"D;�o��2/f/ �ȷ��}�.�����fކ�n��u�ф5Z1�l6�\'f֣��4����hK�o �A�y#p2��.��N�+��_;?h�;��0l@����R� �Hp�G� g�R�����m���kf�����@�y$�	nƥ�+���@S7@��*}zmJ�659w��m����m�j�IY����y��>�W�ֈH�4#��CC ��Hf������4���.��bB��cIɂ_*��[S3�Ҫ��}դ�8J��N�<p&��,#⼰	����	�Y��"����{�6�+���Q���)/J?���������B����ҳ�����w�&S ��u��T0Q�y
3Iz�DI�]�dXWx�����3�$�Ů G[�cA{#��:M�u�T��������$��9M�nO�,%Fd���\�{�:����s��_��d	D�g�"��g�j�U��	K���	�tJD�^����栃�ᤢ�g���C�7�/�&���̋J�`��������޽!�:�R׮��oj>ՙ�GqE�R���(L�K�*`|���Ǝǃ���=�E ���:�儊�J*R k"��||U���m��t%^H�:T�ӭ�M,En ���ҧ�7�gbB�쯂"�l�u�֬;��HJ�^��.�c$^8�Ð� ����C��$F�GE���[����
r�|��8�����%3س��t�a���h_K��Ez>|��az%��V����9��oL�>����q��][v��K�,%���?'<��3�r�`���u)�&���<�fL8(��N\fM��Ng��\��4����x8ѐ�z�t�s_���$Q��
���S����"rwL?�R�������mɏ(�<~���~�q�����Cz�۸����S2" �b���}���&Lځe����3 ���}r-�����Ws��	n3� M�$� X���p�����k���԰$Ef�w�Ȣ���K��!	M��A���j����_H,��h���þ>m�c�{h�c����b�D�(��5x5����Y���hz�z�?��V�O��]6CZ�kvѨF���41��#�� �<)����Lxg��GVUS0�5X�����D�އ�Q��v��(}%D�݈�PQ����ǳt���F�uRv�ٯ�N�w���7��c�?���|�P�B��SR�Nf	�}�
�#8��ֆ4��5����)L�?B���XA�d�	�u���}�P��=�N��k��a���v���L$0�/k6ƛW�6��S�L��������G��7l*	��1��z�<`'����e]��@�b��[������ o�q`��W�Q�V��_�W���$0j�j����hں�ET,����S,�>�U"���7����*Ud�`���4�xM�c��r'^���Z7D�LZ�5˓>*c��I��4���)VRZѳ�b7�wӈo��p���5����z����|۰����N�=��u��͊��+��p�,Ù4���gڱ_b2^��Ѫb�iG�}�'�����!ea��v/~�gܞ<-�U�^�b�za'�CU�c�bc oI�_�
��q4�p�ҧ�Հk�]s *����#��}�U5*]�{�sd���4l;�{���D�W�j��;1p���<��?��ׂ�2�=����%Ͻ>�pB����͢1���u(�;��H�Y�v��Tw��C	��G��8�n�.Ӄ�#4	�
4�i۔�H-r�8(�]����x,W�������T/l{�G	E�!��o+��3K���ަ�R׷�2U^t�گ0J��۬Z���J�d�C9�J��u����̈����\�¦b��;�|�Q��ô����:#�����D}8IЮ3j��C?�ڸ���q��;B��흎fMF�~4jٜ�c�6�N��z:Ed��E�=ԇ�jD��W=fp�5~�$f�~8_:���o�Ӷ1���e!���
��a�b�0��n���t�*��u��d�����������q����rkl�QN���:������p>Џ�H�7�^�e02kn�%�~>���>|9�:���ra4�|�}3:�V35�x�.}��^gpC�Z�Q+� GV&�e3'�%d��ŲF��Nb�fF�R��ϒ�%"P]PQN7h�E=lKnw��(Mr�d���6�C9�ɔP-Èf!X"�G���yE��C�}�(4�� V�u�P\/q�� �����(0%�~Ax����^^ݷ��1�Wƃ�|��G�`���N�y�l<Q3��l����q�7�:v�G��Wsލ��~oh�Ά�?���&��u�Tr�3�V=̗���v�d� w/m�i����>� �K��ײ���t�m�kP3!#�s������S��*c�=jEJĵ�+��>�.�`���d� ��>H�"�6
���u���͓�ј�¶�7{�[�ù\��-K�����hc�ԯM����_U��-Ȑ0LV�!�c�P����0���3C�8p�V�t��sUӯy�U�j������3�nfY\Yz��_��)ZDca�D8&f�Z�`���^�7���g{���V���jнԽ���#���M�w;،6��
�c�v���E�]�k<�����#WA��O�	3�J�����2B�'��>�g�7�%L����QZڃ�b�uc�!��(ͱ�-ϟv�� �5$�s;�	�'�9�!b)H�I����V\�4҈��>�d2�*.���y�4�.������rj��QoK�ݚ,w_v��]���wO#���$�&�����6�i�K�zʐ�?¬w��p�ޓ�r4Q:95�Q�7�ɶ�#3�z�M&⼘ӡC���Q�aR��i����8������R��n�����j�P�(瞆��Z1��+�94g)�M�d�;���7��hy���B�1�sȝ��-��4"��505?F��~m��W��9<k�@^���u��ŀNŜ'y�J���̸?lJf�Ϯ�o�37â�qܻ�*�X��>)V�|H��	�TcJz70�5Y����m�_8x���;\~�G�L�_��3t�~��*�2���(*ţ/Q�B=��Tא��}�^�9����b 3���-�������;*��AlI�q������ZU 7��C�e�W���p!F��H�_|�@:�>�@�����@��>�a�څ�(�	��7�~`&���6���	�V@T��[8^��8�|���ߚ��w�	���:��wO�UO`z8�}��~����4C׊cj77Qsuɺk�+-�7�~S�)NW=�<�9��׏�41W^�2cBEc~��f:ǝY]�ͫ3K���%�z%��y�,�gH��%�Er��Ew�����x�i&ı���^��</�;��|��.���2O��2OmQ�, 1[+�_�a���5��h͹c�c��&!���1_
.������ n���s���Q��}�Fv�����9��a,�w�I#!�H<S�,�_�#����ւdoykeV*$ 4��NQ�=yFb1��a����/a_Hk(�P��{�'~�]rŅ�����Nϒ��/�A;������yw^4о�C�ɔR��e6�9-�+���EO
�M�%@�G��*�!=D2,`J�Md�$i˼�,v��1SL������U"��} C��}W��W��(�y��O���3�KZʄ_ɝ�f�}����@v�l��M1�'��X2���uw�;Kc�]�qy�[�Ӛ�IB��l_��y��M�$&��^ۖ"���$�h���9B-������uT93�6yem��2�C��6��u��	�}�X_�����G�^Qxտ��d��"��@�q���B�Oˠ)���b��d���O��Kv�c�lhg��G��<�"҇�C�tJ����!�<���5|H��j'�9�����Z�1}������SՙA��8q�e�R�`<S��,�f���9�o3x�P�
[��óS�wU�!Q5����g�<����Mb���Eш�~�=5���YXJ���S�X� �lT��ǻ����_; �t�N�]~��!�U䴜'��nB��)�Y��Z���3�Y�Kp�O	�Ğ[)P�pŉp.ǀ�Cl4���j��L�-6����\;v�!F�=�d� �R�׹���3C�jM�V�l}G���M2�X;�>}	�����?
�&Tn5��@�~�n�J[�"j�RPz��H��Ǒ?&�`n�^��2��'��ֱ:�l�U�k�:և�W�H��WdT	�"���z���(|r�G�T�^��^B"�J��"�9$�'h�ҋ<�,S*!P9�za���Zk9�2
:�0�u�gӌ�:��\@`��"Z��?��״B���{U��,�1#��I�tZ�qZ��2c�^� �?h��^�,4`����a��hd���H��̇���]:R�`{V��I$�Km�3�+ԉ���b�=~? ������6���̿��@ �Qі�qM�#U-xs�Ⱦ�dÐ�C5D��\SB���X��M�7U4˼S����9x�h^��BŰ��x�qE@�0s���W�6�@�k�m��*i�L�#�Ra�'���2�6�*�����!�"Q��s%kٍ�V:�T��� b+�G��L���3�_�*�*at��G-8�{
�@���[�Iea.W�!�����3#e�,��!�A�0=��HҼ��z[�e��{X�b����3(����w0�ò86�N2F���mYg�;v���Qi~2w�k�iR�G�_2�:�4����Aٱ�J���cw��������ól2��<�j���+0��Z�}E���,\�8�a;Nm�bfv�P�g����t|\����K�Rh�V];5s� ���T��t/���h�u�bY�v4NHJB����Ip�D�!���<#T��:���)�O�ԗ:]��S�t�>7�4����i%�LF���8,ZD� I ��K�����:n���qVG
T���r��xӸ���L�W<�Q��%|�L��!y�p=��������H-F�ã3��X�_��2�i������[�2��'��Y�[��Zb�o��d?[W�GQ�8��v��:��sAWt����<�G�Q�FG�}%c��gw���~�DzD�sY@�K�%tC�lx�H��-0�l�f��")���uH�v���g��&�yr5}Ͼ?M��"f���7��X�� ��T��x�(�-����z�R�T�V�1|���1&\4�?1���z�3�Mu�f%Q������4@9v}hz?�3a��6��e��fzn�Q5c���-�c�`(}jvR���*��	i�Ȅ���`NrX6�׈J]�����_gy��]�pb�U�dv�a%}�=oT�tw���6&�q|eX�$ �m'ז��� �_��M��6^:Z�4�=�W�OSv'���~���] ��=2g�`�v����*#�����ך^�3Tog;������ukQ<Q�	�K����M9'6�ZO����R�:J�W��e?B6"�/?R�[N�2*IT�� 4'H]�f8�92��f�9��p�f�-������k��ӖI���d�����R��B����K�u��c^EZ#��.���H�~[��<���+�;�
~�љFR�(���}T��,`�<�SQ=$�/L��U��� ;&
{���q�/���7�Wj��.l�u]�l��w3$ԣ��Pu�O氚�6��r�R�4*�;�`�ʽ�$<(��|`�U�(�wl�O�@�]5Q��:�Փ�?e<�#S�"�ظ��3*N["v4S@0�'��~*�Y&0�u��{�fS�>7�O��g�ғ�����L����P�V��iV����(!8{P6B	@��C�U���/�i�K����� 0���%���٧Rp{�	���0��n��QL�'1�����?���$N�2�{�L;[3�dy�eA 82#,6���ѽ���Ղ˞�V+��_̌�O�%T��zI6&���Qe/�L2{DB��f������dA��}����,����s=;�Q�ܐ�����+M� ��wۑXm���y��T=v�֓��D����]������ ?G��_�W�D�8��%�7	��B��x�}�2��N
�}7�������6i3��6�=�kB��k%at[��o��
(`�x~�MPR�H�m�r,�?�xi�]Q4aBU�'$vJ,Qv��:������BY�F���M�>c�ry�������:K��AX_�2�e��o���u�E�; �1���4ͥ���ܶ&�ҕN��}}p�P&��9�T�jb�
��G��`�J�9up� �}_>�b\o����ů��� |�b=A���fǲ�\DtP?�k_��(-�h�c1*��χg�ᖎuk��i"�g
���6f�t2� 9�A�!E�v��E��5O��*UF�V�*�Q���9���(q��;ڇ:����q�����''���;��$��tV�Rт���&�Ղ����m���I�L����\)h�:R:��ӿIK�>׋�|�{��$�/y9���C{�z�QA�ఞNpwӎ�u9����V\��mЌ���j��_������Q����3m�B3��׼��p�s���	£� r�̵���R��P�b?Q\���܆��y��c���uY���U�|��C �p�X֔d6�&�!��3\|�0XTƭ�t��#�#(��ED��_o�̸֪Q
�O���XM�� !�Zj��ܜ��R/q��?�!���qR;�y+��d�'*E-ʎ��:�,���Zl�%e�zؔbWVV�90R�v}.!56�$K
��ڂ�� �c�@j$�ZR4��������g��o��Fo�B�BE$��w�dn��Q�.��ѱ3�+}n`w]�Y!�x��u�R���.��X�����X}Dwe�6X��m�q�C�����{z�K7��}b;r�8m֓�D�P��� /�Eo�(��2|�_�B�H�8��5�M� ��6�=�=w���A<���&�/gt���[������Ѕ!�-0z��7�0���n��@P��U:�d�ғV��~��-mr���-�+�Ի�D�q��������#Sa$�8/���.��nbr�1Xy�*�dbMa��X0���z뾀<���2r^x��m�� !6���Ltf�\���9V5��PPS@�$�1�q�{�d��� ���ʓTY�f.}�#�W��S�bǆ�v��a���T�Թw|����}7���R1��{]0*�ą�]��[4._� x���o�@2v(9@�?�%%oN����}0�q����+,| {VY|20��0C.?G����]�H��[to�A�o)YJ�u�Tu���c��Ƽ�J�A���q��+�_h���ؘ0�r�N�0-�|�;Sw����2�w��o��T(l"���oG7�,Z���@�3��os�<�ej6'����q���.Ygް����4c��x�O�S�xQ�Gu���󮦵O�� u
�c)����um��nYQ�8�h�c���6Gr����*v��@����Fa`�U�[��m3���(�E	���>�P�(�H��Ξƻ(���U�Y��K1��￸V�~A�Y�ł��Mޢ���E���]�B�A�}PQT�F��L�~p����ˮ ��oS�ev��`c&?��d�xJ?:���}������SD�.�7A���E1��Gw=�1{�\@v:�^w~始T��9E���BވU�1����	��c�$]1���=4�c�Q�&�e�4hJ���3����.&��!���"lZ��7W��[g���+����vq�����c����B���u��a��~�4��1�`�;R=�F]ۜe�N����D�� g�8=��/a�å��#��t��i
|�Sr��?���p���~3A� �E��ѩ���C���z�(� �~�MN�e�x��p��q�
{O��!�]�M0S�j\w/�F^���XO�����qfK2�'�&l��{_��4"!�&��A�K1�a�Z�N�k9��ޜ���Q�j�\J�I�\)󟉜�ͥ��Z��Q���$���JZ='w_FC��X�P��z�� ��_ $�wD�.%㑚�`����9J!j�����{Nr�Hs�N�a��vhW��.�v����)���}�x2;��8��Q�5' �9T��_�`�|'$�o�tۜB�{8�6�xE�vw�ȿ���
kEq�Xt���]�:��:�ᝧ|br��ł�6�E�WA���9��i9���L����hA"a��ކ��$�"(�E��pze jD�����䃩t�Ɇ�H L�
�En>f�;U�0Dq{����d_�v���-X,�Y{����&���=4|�}q5�Ͼ1�����d��.�#Xxʀ���m�P�CP��zD�oW|m۔x���Y��T���X�eʾe��'�+���lu*9z���MP�f�iV:�g�q�O��5y�-T�	1�Z^��~���N��fm�[(پz	!o����z3��<��LuI���"7HO�n�;���0^�4M��ҍ���P�B4�;����H!�~��F|=\_ZR���q�!�f�V�� k[>B��d�`��j�Hl��T�G<�Qn����qS��g�@B�hRxO�3�F ����d����6n�Ե͜%:tP\�Q��q@77y�[�l4+�>{aj�x�.��%Y�~���4_A�4�2�N��l`ߵ�a�����ǟ����}GC^���LpBm
�p�O�A���{��ؼ�Q����C&����(��TU���6�*ߐ0P��	NFv�/��ͼr�F��^L�7���8��뉠*�����؊�jwʁ�L5Ի~ 즷Pp�88+�)�������G�W���8Mյ;j-U�����\��R�2��F��Y	==jkH���,�`�N))����4K���r ��x*�{%���H=�˲���+��<���&{xRU����Ͷ\K�-����B��-ߜC���DF�9)��[|Z8̐q����3���z먵Ǧ��R���\�&^�sY$��x�p'�(�%3�O�`���J�J��Ӑq�h\֐��5�A7�W�<{J
�H��C�Ս�P��>��K)H{Ny�Z�72�]�K3�G4��:��	���I�V��aX�'Ӽ7rXKPxDu���ңI��?����괿���F�0�g���Dv�Tf�NH�����8Ք԰Q�7&�J�u �{�g�(25�s����K�ش�Ƣ�����ڌxV����H�
�U����mFf�Nc�|"7P�V]��"d"��B,&�vh��+,�:��Ey���̓+��Q�9�;�`6k�U���˲�P�#+I�Y�aܪ��ս�x�)��ʎ���$)6|��o�޿��޹��ۛ��.�\	���l�7(d/,���8o�e�m�OLǮ�mNw���Q��9M.�"PxĔ_Tt��d$-��%T���֠��t�]�=N7J���x����d1ux{@Y2��1=�L��}�!jʟ�23�O�������'��+O&�U�G��/e6�'�5v��6?��H��p���~p�3����O�z�_��F��.'Z��6cZ�&��j:W�M���,�$���a-��'廫?1�wqj�Ű� G�g��Z�8�
?_DXʮ��ڋ�r��Uphگ�^ś;#��K����������S�ͮ�-f��_���CH�|>��W'���	�6h��m�AA����8H���B�'�O;���
'��CӬ�|i6���K��V�$/�q�
�n �I3�:!.���r~o�hd��*LD�*0�Wpn	�*~��$��!�X�V]�w��ס]��OY��5A�l�^F��g�E�:�9j��ی�b�zFy����SQ�㥈��ۖMҢ��Sb	��]��+�:��y7��sh-p�zp"���-`��٣��
��s"��1Pm7�'������3�����2�(��j6��͒���#U�^L���f�CV�(��6�E����c�wIݢ{�]^7�E^34WZf?��1+�_�S�<`�V�Y�#�c�����D���7�������l��)���k�IF9�N���w��C��zlN VNH�o��W��?O�!�-Q�"{6"�Q�-��Ŕ�m��&����b���(���n��J�P����������xVb6׹1P���tm MY�,��d�� ��սF3D^�zġ�}�6K�V���I��x�&2��~T��ah�y\�/�1.W���mx��Y׈=9�z���I+���.���;�\���R�G���KL_��8��/ �~����)!U�c��k��x�ɚ9�8	A�z��xМ�2.BeJ:Ҳ��Z�<H��燢�����&��I�E�"7/�,XҠB�۬�½$ۡ�� P�?E��6���x����Ÿ���ٻ����c�x��9B$.ߛ��G	��`g��r.3%SJ�t,��2�5�@�0�.�O���IR8�`���t���2�_����1���HK�|~,C����S�a8�@׏(�^������R$��K��	������Tr[�^zoL�/��:����/���^֦�^m;��,R� 	sk��7�Q���<}uȩ�	II�ȡv�\:�^:�e�I�g��
0$2D�<�-�{�Q�zS����8�hA�6�'UAޒ���`�`J �[E�?��/� �Ӌ��+P��u9���:���GM���l=�m/�B���m�s�M΅�>�	�/�ηC������&��|�B�u�I4�M]����|�'��'B�����9$ts��
?@I�Yrp�Q���\����}�5�1X����˓-oG��T)9^���ZGZ�QK���9�3��8����ҷ��H|;u���Ð�nb>ǜ�`/kwOHh���QЅ�1��z��-�t@ɰ��]�V��,���B�E"ak�]����-�*_�KftOHB��r�:�B��+<ʑ���>���ٓ��g��� ~��&�iA{h�p��`mD�
�%�@�@z�q�-ǲ��je9h�M�Q��lM�K��v�2���`�^Y�����Q���pk����y���_�O�0A୭�� �� u���"�0>��E�������1�#&
C��E���[��ki�ͧ�K�i������	>��2�U�!�g�0[k��k]�T|*D��eAD��%[�iT&���\P�"�m�_񅻞%�{��q\.B���9�1ÑH�����rm%�������_9?�ctnk��Bt��ڮ<�'<K����>�Q� vht|O+�D�r�Y��oHU&/ٸ�g���r1�-x)��P�To9���+8�����1�d���:\�w�����"QĖ���R����@g���?ɳ�_23e/���n`4!�o���`��#/��H�X7[d��-n��ז�.p�@b)P�a��hF7x����l�7j��*��ѓ�{�樐Ma���R:�p~Uy6�0��m�A��������Qx��`��J����ר�"<���4�}�ڽ�f�6��/��͵=o�@l�T�Pc�M�l��޹�B�B���<��<��d�㝍�����W;5U8a�Q?
�~B��j�"��3*�=ڌ
� �U�	�&1�	uh�d1t�ו˄e8,W���y�*���M�Kы�.5wQߋ$J6���e���VC�k@
 05CT�F��k��:����! t�8�1t�n	1��~a�H��'7���Xc.� �i.W����y�N�R��6֍�^Σ(I��=��B�f������i��#}�"m$w�g
�^D�A�x���FIH/<���s7u�D`B��LRe��#ֻ�g3��1�ѷ����O`�0�>�J
م��s��-?[���Q�g�-q�l̴���ͧG�\qz�e�;���=6�y�H�"�-"�����/MP����If}�!eEը8�z���y�KX#9��RIh�`�FX<c˫H(�/�4��C}fY,�\E���0�3����Z��$R���t���D[T���$���I[�L�΁���kPZܳ.8�w�{_����U�FpPt�t�:^ �4oY��������WWSʙ�z΋��{s#�����*{�؛��������H|͝�w�VO� ��.���趹*�"�ڞ�SV���/���#������VK\O
^�7|�P�8�|L��^���RZ��7 �V�;h���ZJ��^�K#.�Y,�?�庲
���z�=C)E�c���Q"��&�|��
1\O}���-��iE�6�&]7'WRZ*i ��]�
����-s�S��&�R-����b��G�z�q/���&k�NhR��&�۹:*��Տ���P���a�����n�%R:_��&Q'�1�W	> ""�$�a��Z������=n�^j|jtM�D��7��Un�\1�'�Ѹp��]��5M��m}7Q%�GI��'��ݍ�&��(�a����\���jH�>i�Gk��FܸP��3��t�y�-�%�ޮT��b$&=d|�A��)�f�$�ܿ��ҼR�S�W!�56������;��*+����^8�~�5�^+����
g�؃jrxq������i�GV����~OBΛ�V�u�E`�4<#���CeM�9�[��)Z/�dX�����Č�#H���X���O�?UT_l�g;1�u��j�FS�6��t;T��po��m0X�;�u;�F���V^P���+�a é !	�op<ID�5w�8����� 	���S
����G�y���}]�Q������E���4!��T�0�	Mt[������&���-B���&]���p{���q.5k���$9QF��ď��/�H�i����96.�r!�P���+��^�$�,��>�T�Lo�v�	r_�K;�	��Z8�T���ȕ6����%c�E &�z����{�0�iF����0��~��lRd�lDB@P̝�X ����+�ϊaL���C���#���L(|v)x��i{��A�+�>7�������qSF����!S�ۇ"bxq;!������t�t2�$��j3M�W�$���\�4����4�tua���he-��J��)�?���aE�7����/H��"�w�k�vv2/�����5���9agTCR̡�@ ����ĉ�E��dR����c�e�#{qձ����MU�@�n���u��:Է۩,�8�B)+:��z��d���
���K5B$�B�i@C���Qq���
��h���v��Gt�\Cld�u߾ṭ|��w9��)S.�	HMҟ�J���ݽ�C�`�A �?��`R���g�5���������!�ЯXWJ��O6788�& }Tq�#��!��}��U��[`O}�
��|#@��ېb߉�H��^�Cu��I��6Y��k��0�{A��+�-�ߝ�ӭ�}B�&�e�#��jXk��-�GA�y�PC�W���W�����B�&b Ot�b���΅Ґ�US�a_!���7�ݙ��ԣa �
��+;�0$A����:�P��<�%�Hm������
I)Z	���-��,��v	��kzfx�t'`����¾z�d��q t{�9 2�d�~��cJ	�|�����Z����.���R����W�J�_
�D#�S��n܌f�sb)��Ow�����&}%/�N�?e&:uF���z�$p�רF|�),N���j}��չ����h��'c܄���(�+��u�$��-|r��=�Ss'�W'^�XH%�������+�$��\M?&�޳;���}q�r
K�L\ƈ����Fo�o
#x��_7s��x&~09:�Ĵ\V6����#FȚ��V�k/��"�����s�qY���"��h�V�Q���L1z�����M�@�k���Qr��GA�d�N+@��m�HD��D�k8��4i��Aa!��Ʌ1$�KS��h���n�[��7�Ȟ8us�s�\���;@	�ڟhD�M�0Z�~#�bb�8�ZBQ�������2�=iMK�W����w�_����F���]���XN���_*��&�~;xz����b���v>-�/En����]@U�B�����2U���P"��YZO��=^U��N�c� �E{m2���)>�Fe;mQ;W�Hyr]�6�"HC Yߏ��9�Ǉ�(9�Αl�����VY�2�y��4������� ����]KK�����-|S�^�)硫 ��Ҽ�#�-�3.���퓐*�J4������CsS;ݿ��n�D�Tf�;?�.8�1�ӌ�[��ǋ4, �្?NL�I��c��Rh��hGDR�n�����f�b�d~hY���GD셗tO����?��,K��4�V�#S������z�;�;QiW ����Re׺S1�I&zw ����i��%�-�j�P��`�j�&�#u������ī�#$�&8o�AA%�]ل����b]�w��z�J'�]K�`&Z��:��(V����޼�?J7��G+yw��)<���N�7��%
�Mǂ��Z��A�3�#�C$X����Ƥ���^����Є�+�祚����~��SԘO]���v����Ӄ.���n��zt��混0JMF�)��|,L�`L��5�4`ֽ�N�AX�i�R%�QL�AܓE/���(��Y;���O-�<�2��k��*!�B� �yXq����ԹR}���D�"R("����B���c�X�W%toX�bt7�:�ȗhDw�V>��;��TSr�]\gQT
F/R������nҸ��4I��g��SC��T��އӂ;�r�T��ebH�P�M�xK�1��W�x"� KF��i�?�̃�.KJ_L&���S�h��W�1��w>��G�0��h=�#�JhR%jߛ�1������xNNZ�#<e����4���'���*_�	R%5�M�,+�E�Rȡ,Br)u���o����&��w��e�bu�D�p2���6\�۵��T����ݤl�I-�u^�x�`Еd�\�C�2�Ԯӧ���m�&����c�G������{��"�K�"|�&$8R�N�ѹ�N�<X��?Eb/��"�Έ����I����i���S��L.�.�g��=_�t```l���f��bE�wOYhyΜ��S\+Ye�]��_�{LT�I
}.����GՅj��M�'P\!����k�gw�w8����D�f���u$���6=�\�)��S���؄$+��d�H':sH��|t���E9P[���5��.f��5�Q����"��J(R2�/x��1�Y�CE�񭑕X���j���>�'��DX���z*c���nN� ���jŌ��v�Т�~�+�j]`T n�14���󯥧s^v�Ő9��G`����;��  c�GSm�wدZ�s�����	�#��7��B�������qe�G���~�p�p�F7�
�+�mw1�����C��!Pe�ۈR6@� K�G�.G�o���Pa8Pt ?WFZnXd�`���H(��G�!��Q:� _k�1���BS�o��s|`R��l��}T�qĝM�G�!9;M�v��W�'�-i"Vh�c{��.�1dt�T/��x�.��+ƛp�W�<p�9,E���,���8�J�fy�Y\f�W�1���OÄmc�z�3
)<�2��K=ux� �0�V�q�=P�w�SFb۠zwl�(���܄�-���)��>�������Qoj� ʈ7 �g��q�{a���*��=6!ʉy�z}N���}^�M>�+��4Ƀ�Yu(v��1��y��Ț*�������ZY����Ѳy���O&�`��=�	�*P�ay��Js�\���[!8Tp	���UE_���$Q� �ГJF�
����Ȧ�ڦ-Rys���9��/�=�_#��Y�6�v��p(_�_W�:�6�a)��v~B�b�'XR�S9��$}��qhܸTN~��:o2�����gs@u�@l%,�.���j�^�B?����~<�^;���w�s�x�gX�}�������(=�ɼS��1zA��Zz��A��1z�j�����z�'+��mzg�* �=ګ�����u�WBt*p�y?�+[�%yR��ƀ�1��Dr�V�Y�Fф�y�źlw���
.ٮ2����Dc��u��}��&$
�x[y��[ <n/����gp�_&���ͺ���Dʱ4$u�X�E$����d�;v��+}L��P�1l� c/Ȧ�@SF*�*� L��K�lC�`1��{"s�\��h����kyH�օ�!�|am��X��6ȍ���b�>�cN����n{ ����?�?Bf����BŖ@�E�,z�p �Y�H$$��1l�_>wk�&�9hdƗ�<�J?x�r��[�o��%���)�=7������tt
��'l7(+۠����XN�e��*.�R�=�8�k�ֱ��ɿ��� �H	��v���<
1
����&�u�×���w�#�g�$+��ǻR -2�N�]�5x�]=�<��e���)`�a��P�"E�H����ʎn�4�Pr:�� ���ɠ��&Y�Hnn_�b7�@ ˗�f��jZB�r{�\J����8f�xWZ����̜iCϠ��,K�	$���Aͧ��s�Mc���G&�ژ���s�6�Y�N_��>���JAMQ�ʝ.��o7�N`	M��Z��"hXF�H��-�c����T��#�i���@�4�p���̨k�z��e�x�K���y���+w��^d�*�ֹ�i��ަ�c�|�T�;�%yk�ڕ��ߚ��'���b�ᩍ[��OV�X�+�2�/ƻ8������obS5[X`l^�kO��fJ��6��Y��ȝ�Pr����S_�-ޛ�Gm 9�����<x�W 1��_z<��!╞���[�D��4��ň�����_�=�>؈U-p����h�@��I�S�_�vc�/�^���
B���t���
$��*�;�E����~Y��Kp��qK��~�f��˗��ԧ�c�4l~�}�0&_/��R��9�Y�ݭq��0{un�����B2�|�+*��e�,��K&�j����+�¨̃-�.��2QԽ��k@�j>6��u�D�N�.jA�${��J}����1������1(��n(3�����ئ���K����?�:�1�,
g�P�Q�ŉ��i���⃓�q��da��(
Bs�\9=5��l�(jS{��fY�E�6����е�uW�:v�9u��4�L����2RF�%�D���R��0wJ\�����Ԧ@��J���7�Nh���K�v4������	�8�Xu���8���1�=�w���"�� w�c�nu�#�1Iz�D}�^���?���� ˲Jl�	xO�dN��/|����9;i�Y� ��6�^��b���ǜ���5�����/>JXt� /�ul���YhC�b�K�!����[[Z9�OQ俐^hU��;��{��͇��LáX�̛��9[{ؖ��`Jd�z�˰El���/j�u�����-_������(/��e�E�rc!����i1(=)hV�-�`��#=Nʾ-\��/��aü*��\8��:A;<���՞�7ٮ��)Tʈ�g�����*fӱ�2Ό~��*��/
pO�WQ�+�~WB��/�d�z)�h�oO�ـ1����5W|=*CLp";k)���=x�X���ĭ��Z��ȧ4d���Xa|��K{.�B��W���%��t�����΃�'�E�^�ª]4�	�d�"����7�ܸf�[ w7���(^W���r�c�I�fU�_�����I��֔�O3�c��XNWl801�x�n�lliq��v������Y��!k?x�Wرc��C^6&����D���M�m]�}b����t(U�g:ar?P42G��Fo�_���N�UTl������cBowe��Z >W�5����o#�~hY��%(�f�O�0z����<�u����6�tEO\�,��r@a�;j?A��)�M�9Tpl�&��Ч�=T�Os�c�!�;_u��"����F��,Y`?�q"�\/bQ�� P��$�������b)���q��,�p�z�cO�h����G)l�䉓��K�����AO�B����&�� �S�����#H��H�DPT�'���]�`x"-ZLYF�i�2�6�É��E$5���|�W�7z����^���.�E| v
��b��;K�Uz2�ۺ�%�t�]f��+H��y���\�i;��_��hsp�o�?�͝�P�+���fY2�ő7F��8��ϯ�YxLhD��y�E�a��V�@���~�bQ���JI���o߯�:D�^��#r\v"u���[̼�JЄD����F�� ���
rݑ������*jb��c�j���.���We=H����i���L�\-ߘZ2"5t����ǁ�IY2�m��yL�ѫ;�#�M�q�_�+�j���&��6l�p`�S�"����[a�4lO�"�� �dv4S�o!%�pk�E���.r��d7N]߫=�`�"���2M�ԂW�����3��j�u��@�3��y?-;I��ǎX������|YH?���tW�=�#���S����&�����j?����T�%kЏ�� �!��'�p"��X^.�80����U�s+}Q����ё!
������d��F����Ǥ�����G��u,�b�4�=����F�o�2��W�n�������@�x��(#0,�F�IG��K��l�M�d�cʭ�K�}jnw����a��I�ޙO@�j��8E�N��ԇfY�
�r�m�j��.��j)��|$��q��!q鴇)l�A���Ò�n�q�D�E�#ly�ol�zg{&���X��}�eҩ��R��n��eU��.'�
j9c��c:X�T�1�\����\�"��lU���a�@_֒ �sjF��*��D������&�I��k�茷���+�"�k�K��C�r��x��M�{};l���OgE8��,��Z7t~�\�Nf**%�3.�e)�7����S�P�Vh$%�	��VϬItz� &�5�b�U�:P�׃;a�f�P��)�|���혌���$(j5Oj� ������2I"&�� ,�q�J�ܓ��hd�CP�" ��i�pV��zs?�P�8W�Řgpp��c=vh,@������N`����/��&u�y>��u=.y\��2h��*53@Ȋ��0�u�6�����7����(S|��_gҙ]��{��k�@�֤��@�6���m��iԚB���X�۟(z���i�.�o
����L�d��G�M^��)ђbz`�c���zi�D#P�Y�S+y��\��"���j6��R�Q'���L�KO����B&',N�~۳�C�����w��1b��A�����������X��y�KZ�Wj<_�RlB1����x����]%*�	�n�8� ����|%)�i��((�|ERvX�%��t�~rKXn�-)���8����P��IӀ���;��w�\P(FK�.v�P ����b�b�3d̎g-^/�HчǴ�=5ۓ��F�-�fĩ����W
�cEI����/�ڪ��vy�^�װl�?�Xb'�=�%ED����T�Mr	����
4��h���������ϧc��KX��i�$��x���/&���乘 �3�:�ˍ�ʍL�;�[|Ql§L��g�X�k��jY���ٽ�9D��e�4�	q�m�ɿٸ��_�:OV4ݝ��?Lr;s{�j���5���Ytm�� J��ػ��6�UFB��?�h\�R���U�o�vmR2�Ԑ=.���m�+�̈́�^�Wi�Vg+��L�ai��:{}�����ǌ�N8�,E�JO�Wή�C�ve���&�h�SS��I���#��죃��\,�xM84@�L�Ө޴笢\�����~&�g�A�����]��`4�W�v�j�t.�KE7��Ok5"I��GHf���7����A��Fk8a����We���s�`
���E+~:�:�l;E���t=q��۱�Od��Cm�4�G�AW�vI��jg�Gtj&�r5�r��7_�4$?z�1N	X͢8�Ql	_���aĸw?��ؚ���&�p�u�q��S�f�����V��L�ϛ_;�һM��B�ͦ�WL��}��T�!ȫ2�J���}�b*~�!�޴�V�UkgC��!<�J�x�����jP��Vlۖ;�HB��$�����*{oĢ$��#�[^��|��_皝��Mi^�7�I�n�0Pg�N�l�^FRJ��W]�H�k(>b}4�����n�r`ա=s�\��+��a^�(��E��H=\��czb.]Q�K�5�� Ы�5C���x�
�a9�+����@��G/D�U���u=��=��z���ht˳��h���k�7!ߝ0۳% gT 6q@k<�8�J[����*���{�~;��b<��ҷ ��ұ���>D�٪�BY6HU\�C<L.^�_޴��v��aP*�M�zHH�x�n�t�`�"��S]ۨWCR�2L��[�0��`��ل�>�3"�fȟ��`\����a%��p�P��ϑ ���F7�`����CN��?��$yw�x�������z��'k�"ɹ��֞�+A���pT!����$�����9Z���wE�'��ͅb�L���4!��݌�
���p��pD���w�k��?�0������诇/��6Q�Ұ�U�b��2r=�'/u��7F���9w��fAl�h�V����7�osi-ܢ��LS�z��"�I~ϴ�9p,���e~
���a���KxYtDI)G��uFv��
�'��Oo�{|C��7�2r�	�sz�ۅ��"��6��=��a�N�ѣ�rr��,���&p j�����~��c�	s�x�D-�4��z�RT�gϲ�~۔��,�ݸ�v�JKy�����4/�dЂ�|Ȭ�m�?�,�qP{dxAI��(*h��w�a5zέ����L�>[�I5l����N�j��u���[�WY�g�p��Y<�7�&������Ur@f�������&��N3;��~��&�h��O�X�M��=�|��>Ѥ�82,�*�%��@�/��ԫM�/g���O�7:%�q��:]�7�g�R���`Brl��G㶓�����ܙg�D�HW��<��,�!��c�ݣA�a�TbD���d[��}�YruHV��_���:w�!>��/mo<0,�i]X����d�:���|Z��#�x�k��_�fW[Qe��J��k��X��Bn!4ߏ��( ��X^��]�|��	^Q|��	0���Ȱ"c��@a��]thy�1dKi�������~��[ʈ������K�����Z����n>;���?W%�nաLq)a\��:�Äu%̧qb[�^���&���t���l
h���Mn{.�X8�Y}Q��s/�Kȧ����e�,9K���$%Zh!U~�lyZ�0����<#��E���C7<��g�h�hR�f]Wѝ���A!A�3���<����l��{9��ih���1�a��ȓY�8$���i�(0g����R��D�aEɧmͺ���mt_ߩz� �S�g�z����W����վ�G���w����o�`���z�dc�IK�A��63�u���Hn���t�T��qa�i��k'���V"��b�-���$�)��f�h�^�~r�HMCR$g���Jg��w�Cy�_�K���-�Κ�~���N��2,��� ��n����m#$����wGt�N����q�$+���HE�2�*+#�Z��k�w� ��x� ��q����'7:Fk��y�������u�Ā2B�DwiЬ�΢�L���I�:�̊��g.���/��W5/�8-)��^];Z,�=�wc�*,�yJHy`�$�QC��P���e7apۭQ�����[0�s0:(a%���j��L(y[$`q�p��z��u?	�.�x�K�<����4�V�����b�ޭ�(��Ԋ�͐C�"�X�r��g�� x��,��,#f%��O]1��20��4jd:2�(Cg�6Zh����{���O]k�	@�I6c�<zbP�����\%�� ǫ�|�c�ᠿ�]8��O���[ܽ��m*  %��w������lA�q'�W,Սg)�G͟��<�zH�kI:k�C�8�-�q������<�]|���ec������j���#j��s��q޳>�˼G�,�4	$�x�Ѷ��(���4bM$�ϩ��R�g)��fڅ��=5�Ň�_f�vn�&!����=�U>^ruf�<"�hs0ؐ��'�o�~ەq^5�,���#��W��=A8xD���ſ�$?ےv�j�Tz�)^��k���0��Z���.�ң�R�_!,O�kYz�4�L�g��$O��Y�[���>���d��J�#�ѐ*<��}�R!h�'CO\ ���_@w"Gz���4�S�x�'9��l�7����؞4��*�!�Ӽ�%�B.��>`��vsk��3u�������	=�A��N^�(���e�0.ew���J�ٲF�$�<�q��#�$9�ϟ��hkZI�������"�;�!��x�$/��+ ���+:��b<��O<NK5�S��
P��n
l�d�	��XX�j�ed2�J��-H�ugE4eD`e��v<*��0!�u'�z�/n�9���{�cn1�G{qqښ�|i���5��4=�7�Mg�|�$Y�a�h�d��Q�`�;���4=R�m���#ȭ�pJ�a�w7�gI����Q͓$έ�O^����X�C^��k0I7J�^@~�`
e��,�*� ���x�1��a�;I�@�(+�F���tٰ	�{�p����w����8�do�f�',��6~�h$��J�:�^���,�ڿm�.�YI�=�K�G�����#
���J�yv��q���������SsLU�)�{��,�[^�j��<,Rs�-�Y���&��"����u*p�Z��*Wr�
q}58��j	#�o1")��<$�he�uB�:;�!�o���_}g��E����������W����;�Dλ��32�4�&�v��mt��X����E[�}�xW~&<���H���R1%(,��<r1Y�uɪ�
.f�g��f�n7�"����F����9F�3�bAD��2�B�]p?d���x������5�0k}�3'p;����\I��)y�'o��/�"$�D��1��r�Dgkra��"y�Tu>��u����9��y�H���Է\$�ߛIA�K�v��8Ճ���#S;�E�n���n�󄱰!!S�H\��b=~c%[�$��ۮ<{���<��eBe�<4�ܕ�<������w�SbX<�Ju�gW#BW`/C��s�DYb6)c��B���%��3��i{�J�q2A��{����u7����(�#r�3ݨ�tv̌|���+��-�7DMjk?_�ڬ�>7�bUuȸ��BR�0�Q0�����������␍vpV� �R���;���&t�l�bѝ��J�YK^h̛�����7�Ӵ]�oJ쎾D@KԪO+�ߦ5�^��ZwVh����5��?\]����}T�M�W�����Ȫ���%�H�h �:�fE�T�#Du�F]���{.�a����Z6�]R%|i5�Ѱ�!��D�O0e��<D�ls���x3_/���~ �m��y�ъo,��:u����kc�1�����ᆾ�ݒ�"�	۠3�-���%b�&B eܷ� w!{���Q��C�`{#�����e�;8����,�C�����-���#&����IG�і�V�FOxa&��@���W�T�����,�\4HB,�١���JU����بE"?}��jjnH���j�S�l
	��w(G�O�э�p��y����Q�4K��G�;�t?��t�����q	.�.�U;֢5��	�5��,'��\�n#3��O�����܇�G�9�$o�:ſfoD��bԛ�#)+H>�7��m�x��꥖ZVDKG��;��UO:�/���ؤ*8�v�yB����}���Q�]��ۯ�s��{�t����b�a\������Ry�ho��n��1 n�4���6�;����X��wI��������j�J9��k��y�u������1�RD�׻�\���9����A�Z���-vY�����ͥ��sT�U#H��D/Q�5�z%ec�׬�c@Ex�
5@Ú�QmH�~��zK��&�L�����D����M���֟���ͻ"� ��g3=�(��9P� �5�K<%F�B2&�a�OU۩�:N#��q�IV~#T�%2�����4CfӸJ�/CO��4O��m�fu�)��e�2�bS\��6 �y�t�ne)k0+@��ŧuG�I���$��"nӀ&uL�9齪�3#C?�x(�ʬ�3"�,�a�ǻth�������>8^,F��@��u1�G�g�-�q5��'�7��j.t����^����Aܱ���Ǥ��]  j�BXXm�et6}�Z�ii[b
\���D���^��W%�e��H�nF��,Ld#�+I��N�q�{+k˲���������KT�)�	�e���apN�Of	H���<e�I����D�D�Zx���P0���nk>��ܹ��4�vL��0���#��Tk�f;��������Z`��o�M��@��,�[5@z����񣷬�x�W�����ܯİ}yh��b�G�p&h�a��3*���T�j �)��k�HK��Mr*�\7��J�צ��˦F�H�Q��4�˪P` Ɔ0t{ʩW���n�9
��*.#�3#�DU�K��OF��7�Q�uV��O�Q�xǙg��z]�h���K�}�J�76 �%;yw�n��M�	c-���~"�;��AO"�a���th[�olpH$�/r��KK���V泞��XCh���l!?2��PDEe�όbSj��`ۓ���3څ}����3��(C����ړ5X�X J�@�=��o$l�k�ɶ�$3ܕW�d[��.��߶FM��z��C?�3'��/��,6N�D���1d%���q=�GM�5��J� �}�kfTT��wj$�%�hI�j���VtD��o/�3K"��EU��~����@���w���w )���7�V�Q+������l)�ʕ��b��W��<Ɖm�p���]�t�u���|�(`���a�>ѫ����@�s{���\K켝�\��e�/_�yXa d����y*���6xci^a�}���[���,t�*Dr$
t˂��]b�o(Θ�UF�՛sB��'_�Q�JO�c������a�Q%Q�*(S3Mw������f����f��I<�nHo��Z�V��f���%��8��`����*^�YC�K��%̌���'<�.	��4�e9�ڶ���؋2=�%��:��?J?ƴ��	�p671r�bh�<g�!�%���l�&Hn7�&#h]]O�\c�υR����0Xk4�^���GҦ	�Q�>�I(^5�2�/�V�wg��On;T�#�Ѝy��6��'�s�2�4�b	���B�_�94/X#��Q(2��ټpRUSZ;�l(¶�_�C�#���z?��`���Zy��]�tM�����}_//.���]��j޸�X���#?4����#B%.��6fz��0���k)�f�w����a����`WG�O���K��X=ē��z���0���c�)rT$�ϒ ߕ����jB�v�qw :5Z�K�����)�E`KDEUh*��n��aAw�h���oz�sYܶ1R�P��s�R|���&�o�휭qH����|[,���=�'�N�kB�:�/ơg�Q�QND��(h�Om����5�qJ/4����7]�8��J�V��OJ�rc���`-빷s':\qk��t��D���-�
t�c�L����2�Ak"nn�I��r������Pe�����)�q8v����̦m�C$o�Q���>������!��}�>�?a�~��]V����D�������(��2�~e��9�=��*5��&��ăl@�T�8r�Ԗ����as'&
m�q�Q\����j������(m��GsF"�sKX���NG����]�'Q����׻6�!����wqІ�,#�`�U���{8�"s��{o�Ҽ����������d.6��_�9�=���o����¡�� ������q��Z�ND^�nD��"B����xQ8 �F\T�9��y�|�g��Up�`�x��!K���[�tt��&g?��g��0�/#�|	�C� ۉ�#�{L-i� 1�5R��w��`��TV>�P���E\\��9`7v���u�I�s:3�r�X\f�@ܞ3�V��7Ό
�u��ƥ�z�q�t����d�hs���5t(:��4�#�#�k�Zm��ծ>|W<�5_���df��/څ��r�Mr�k� ���֧`��Լ���ʧ��m�O`��P�����y��1�-��sm�!�+½r����u+G[A��5��A�Y��Xp F�~��L}�Ҍml��*B'<{�?���ǧ��vN�K�T�݀`,��*�����<��;�9�+��%�5I^୙)q}!(���n��w�%<HxdAX�nP��i%>���� �g"���L1���_��ޙ����}IW�O�2 J
<�\��+�������h,������u�H���޷��7�1S���@Zxf𙋔���=��"է�7f�&4�w=���x�E���Y�;Q���T�^?���v���	���Ìn��QT�U�)�1A���Dۜ+���^�Z,w�D�.nR�֝m.��×=1����q��ż���1஛�a�2�����Y�)Ls�SvΨf�D
�:n����?ci���vo�Q�nחN��@���#��NTg\�t釞c�8�ny�Z{@ZxD�l*'j�Z���+n_�?��o>L%沘l���b���P �3����y��'����4�'O�8�����
"A��3�UI��v�7�RS�*�:"{�_�M�>:]�4SqtG�	@��;2�W�%8C�@�BN�d�CU���97L�M���dP�0�L�wU�=�a�ٙ���
�j��	�����ǖ$#��y�A\�l��@▛�=A���%�9��Ķig�Ŧ^��F��Z��_J)���-{���G�{o���"�[&K�\D��jxB�@r�p��&.���t��+��A�49��ީ� ��*��f;(��F����:��@x����fy��qY��y���Z���R�� 0�"q�j|Ś�vZM����J��n�N=�
�C���Ck�AND]���I�V�`��<a��M>
1)��r��_�c�CH��l)9P�S&���9�6�^�A�AS�A���!����j�6��^�E�I��xv�}��l;���Sq��O���Iv�`)�\��M�Ze����Z�J�c�V���S����D�S"Q��(���"2��9��l�j�B%����.[(�Ṡnq�k��G�b� �i{�4�`?�Y�����;}�p`;e"��u�I��j8z��ݻ����l��V9��;�z�]�A�2�mF���5�g��s81�I��`�yg�{"G�^�s�HVl}9l����7�jd{�Q-�.D�*|�9���=�񤀕���<4h�]Ho$B�����*#۸պ�������ۤ���B�]� ��4u�Vx��2[*���1��>OFI�����5�߿)���h��T�3q���i9/0O��{��%��~�]���g6,2S�V�׃Gg,tFSr��N�]%����9�xF0�0D�8��16���]���Ys�=B����a�����N�s>�α��/u|��/�b3�s�r��x������'�X��T1u������8�荪/n����x��w6Y}�b�#%L��Z�J�&�"�o*��d6z�G��H�=3�� "�%�8"���M����G�7ʛ�XKC�k:�Οd\ƌ9��ʮ��S����4�_i��J�cZ��*�	�.�ا��;C���؇܅Z�~�� �
Q�X�`�����;�)ā 珣oỹ����l'ڒ��*�L�~v���d	�������	M'�]��M�j�B���W4��" ��0 �%�)�{5GL��1�.j��C˅9�ܰ�EH��;~�(��@�s�>�<�e
&v�N�o�=諱�e��\��ui�����'W�^A�-�]2�ߺ�w9�׈��:3^�$�*�BUƂ|CX,�N�-k}�P��T����+�����t`�wӋd̀#�%_�)c�7�����*���֢� ��k�E�#�Z�Z���,���i�ЁN/i��4��܇�FA��WQ����,�D������� %I	R�^����8��vpϗ�-���hM�Ş)�=|M|�bd-�,,����7g�0�T�o�`6E70���z��.N�}�e�2_���d���F1q�n���k��AI:E���@��A�O��FB��h2V�S��^��4kAsT�t9�`��XMf_�D7j'U=D�vG��-�f�D����_�4C^���u5���N�v���`��!�����bG�t"����tS��_����f^f��Fwر&|F�:�.� Z�~�ZnLhwLOSKPY�.����O�	��u�GS��Nz�ix*�!�i��n���jg�3MF@Ji3���|9�����`��	����	mJ}�P�L�@i�
���c���˽�p1�W^x*�\��3g
Vܧo���}�>i�Z�N�jx�\NM�����y�L����7"6_F��_�*�b-F:��Ƈ���iǎad����|��-�@{�~g��P�~���N묔����CH��PH���83��M��.���׆� p����hN/��q��6���3�]{O1!"8)4�#�|	L�I�&��)S�h>ؐn5����ӏ�P�R)��Q��#��,k8�=��ã�3�@��;���dV,M�,:�{Z�'�#��ڠ����6���!̹���̇�k9%j�'L}~�y�n���@Ӿ�S�~@��@���)<|��	0zZ���at Ò�r������Ec�x�]X�Zr<�xn�~�q��:�cP�	!c��d`��g
���u<!
mY��D�pt+�|�T�GI�8���Y����C���j����bK�!�����LEu�<��_�^.a`���U�zBW%H����������Q}�Vgs�{�Ͼ�D��{7�����97�?X��m����������Xj<�"P�������G�C�Ą�Qe#�T�a�L��%�{B�$icT51�%b�s��A����ݽ�Ï:%��T�؞���d��*�Ң��֧�q��L1Z�*�!�1?���e�/��tu�}��&C���9�Y���A����mщ�|O��%F&�(�l|��_5�&M/#Ҙ�Y��V!�B4�)�-��=�l����\ː ,��=�sS;�z���܍�E4��������k���#S���؁X�@�*W:�8�l����4��H1-�kX���B�$��+����'��Y�tO�v��6��]s�u��CӉ�ԍʊ���~;j9.�FqnS���|���GxK&Sv����K� �D�zw�z�"c袶�@�0���+�������
`�!)�;@u�W9�w����B�
[�v���_u�����D!��=������}�
ˠN�B�#��W�?�Z����"L���r�6�$���x�V�H�/��~��*ƣ� 5=�@�R8Jun9�Q����ۡ�
r�AR�!F�bp1�gmr%gW�3l�ȁK�v����VԸ�J��[��d�%�����)�!��h�e�1Ϟ�V�_�v)��k���d��L���f�n�3�L�e�},�C��vv��%<�F3X�����8��|`��\�h�r��`����3Y���# � B�'�y�X����}���A���O��]-b�dmg ?u�;�9��(E���X�T���B{���UXԌ�oð�yW]+I�-���l��.�|�I���t��i�X��i��w<��$��nݷ@:���`�Cd��֯�e���J��UR�=��B!QwүQ��$Y��a��ɂ�Ыrv+[�����H������F�b4K����)Voz��F,jc�`qֲl�>xnF44�"s��h������
r��
ƚ�M���
��o.�Hn\��w}�H��+)�Z��!JD���^�2��d,T�5�m�f[J�2�zf֗�{���st��\dG)����̀?��{��&�G�e���x��c*�Lu+'�@L���K1�y}$��8�w���n���ܥ��R�8���/�vi�nߧƲ��"�(l��a��x0b_�^A�F�B[�s[�G�>un��j��'���:0T^f���B��T\R:C#�#q�eFg+#���DY�B��s��ǿlz.����(p�/��L%{��/U��%���%vk�Zc6��i����*�I�驋ё!��^����y�q!�Qf ��7�P���H=����G�.u}v�F�C-xΉׁ"����uP���7�|~J�j���oO��v�hap֖�'g�|�+W���M
ֿ?���Z.1�	G`���\������'T�5AFj�rs)nB�)]f{:Tnxbf��V8�aV{KMx��GL+�I$�o��)k�;PV���z�����~O]h]� �"����&����p��hT߂+��8/Z����O��g֬%c'\%1?2�#*;�=}���3�I�	�ܰn���؎/�������ŅG���Vi8�B7�:��Bc$�|?��/8��ұ����)��_`s�b)=Ds�o��s�B��T��z�N��G�VV��3C�؃���[���!�Ċ�g�����7��Vj�!��{[o+��Y���������p����wğa	r*�Z�Z>g�r� ��3������r�F� m߅;1�V�e�3K����.\nu�:�´�H�����D��pT v��m�����:�(q��`hj=c}4K�"�����_gN[ŉv�LR��
+��H����$�3��|������H���*���<��i ��"����=�WF4����m�L�Iq<r�A&@ǠŋFS�K����+�[��|7��q��![V���.�4i��(s�����E!{hۨ��&�Gp	�����tP�.r��zv�,0��_�߫BO�cGeva,���߷lM�V�8醰���;�q����p+Sא��c~�E���4�C�n�	5��w�!��p���PkC�٭}�(�_ٕ���B�(�o�ѹ�n�7���.P�8�~���ǔ]9��e�-�a�rMo�-v	�7t����2���|�D?j��5�y9�#ь�H6��5%�t"��BɲG$�O�+�T��j��M"|�Eo|@;S�њ�!���E���͓K�V�|i̜\�(�Ԇ4�س_�NN����X0�9�V`�̍@��,���'x�\2��b�I���O�J�>�%Iv��.¾ &_tT���9�
S�f�s�$��x6ʈ�]��E�b9�� ��dO_�Bw���X d�����4st�����|�|y�r{{mu]��C�8��|WR���9�me'��]-��=B�!0-�*�i���*�O;��g<5���V�Z�V��y"�q�v+���+'��x���ŷ��4�R�q�E����:��`n{am�^�{�Vٓ#�zzG�{~0�1��4�ܽ��L�&Nd��-�����;\������$̀0��A�E �P���d����#���ߋ5E��J��P�E3�}�i����!��Ģ�4A}�b�V�Qs����861@��;��>����3)�!�������͠���[`�(5ʐ�_�#-�0n^�A��ky�3�y<}u�8(!��5�W��>�9�`���m�ۺ�A�֖b@̠]<T`ij<�GH�:�70;��rz�{�?p�G
�=_�C������@�������#9|~f$@;�9Sˤ����}`��Me�jm�*�#��5�q��&;�:~؛-��~�V��s�=�����:'���QFE(BI�вHu����+��t���]ȔKc	}�B{�:��F��G9#@=,��S�}`�|O��(@��Ԅ�����7d�z_iל��D^�����,3;�]��f�
����J$��F��Z&!?��8��_�&�@I�O�F���6�ܦ����r��	�ܭ�'���=�1E��(��(
'��|�<_�� {�&�M��);=2Y���T�����@-�f\�"4�N#¨�n�`�� /�����(���NaK����g�b���[�����<���%��i��{K��'ܵ�D���6�Yn���A��"��G����DO�PѠqd�����R���Ht���g�dL�踩��T���5�q���x���p5W�V9��N �	,�rw"�ؤ m�!㕿y6b�t�Rt>�Gbr��`V��6�n$c�
U���z>�_��)%O)��sԈ��5�W#��|�01b����l7[����}[��q�#m�2��3f�v�8^�H�l�� /�������7�w�$�0�f9#�	�#��]��3�p.׈���!�g_.�^6Q���@9dz��\6�����ap {�"��B;e��G����:�����m�z� �_�����a��[̛�][�]�_hÄ���&����5�:נh~$u�����N0}��ե�>���0�����t��¨�ӊ�e�@d������K �)!�H�	.(n�E��Z��vK
����9&{" �b�Չ�
.�O�>��g%X$�/����k�9rkV ���\ X^zE׮��BH�)�70�L�÷5��)�]2eMmw+�q�2��X
7{�B'Y����v�O�%�z�Ew�m���nhH���w��N Q$�u&/Y�xi�j�ڠ�^�Ap*OR	LE�����0	5b?���͑y�<zA:A��������%�A<��o��V����͝u��G���Y����w�bSӥƬ[�W�t�Z�4�ۭ�w[U��W�V�o�E�����M���*���j�I,�Neܢ�튲P�M��F��7����Ȝ�̃ue���%r�����я�L�r�z~�ݩ�p@m��xN���wU�D>x�JL=��_F7�(����m�u���v��Ԇ x�/,j��8��}k�=�����JR�I{���0��.mo�;?�H���D��|@������#�~%�k��eX<1� `��N�`Nió���-��R&;��E��-S�wØ[m1�'��&T$��������MC�W�<rc�l V�	�љ�
est����GV��hH����@��%��Ql��[��
�:`B�Kl���¾u������,ρ�N}*�g(	�����+<��B��q�0di�P�����g8:�g~�d��_\�Udww�hfl6��1/w�d�L����4�&F�v��D��jp���� p�D����2���>�q�s�G�U����ށ�Z�>y��wUn����/����#rO����p�'��CD}����R�7�Gz�P#9F�g��U�-����({�~ ������L�v<t(�V��S����Y��<������m͂s���}ReW�=�eM5�4#_[�f�5e[�vP�Ir\s�a�V���3�\����ԏ��P0��Y�[�Z)9�Y�i����[F�9(�Ҫ�f'�����^ݒz��e|�^Ћ9D�����)0�)��%18���?��go$oM;`1�6�8�j�D9V[�������	R{X�ɹ*&���_��Z��<y���\�qfw�o��N�,E�q�\M�O^S�O�]Ē�Q���b����<�g[HOn½)�{?RX���j:�,��}��$��ծ�DTǜ����v�,+>U��ʲ��������I��Е�h�lT�^'o��I��\���w{F�#�)\���66S�b=��Q<lק2��N��D^�D虠��a�v~����ޜ��/erk̨�~=F����~]�?F'	�����+h��҄O�`�0`Kf�_��z���&��Y�
���U����V"EX��6�\̥�X�����z<��(�5��V��Y��i��������¸Z�Up��'($�*�C6�<���G�:�ǰ�)�"yE�<��h��.�MY7�3�u��iJ��� д�X�DhP���_Ou�N�f��sG.�s@�-RMȗ���;���~�U7�-n���a�C�dWV��zö߈�E���^p�J�q
�U���,}���2����8�������q�n�)0�P�� ���؉���'A�6L�2��E&,�y���L��eq�ה���w =7<���42�v�����^��i "L���0JU��9 �H�[��X"�Ԏ��2�GB7s׋�pML�P� �\��F�Y?�0��5-,O��(�|�Y����pә��F��]˾�����QE�j]j�8>�/�:���Nf��.Q����:�\)��,����U���eh�B'h�rMm
�����Ib.N�՛"��c��&������Or"�zQ�h�m��Y�ʶ�Ǽ?�C~���D�e���󯟭'&gE������NvQ�o��_n�Y]��5�.芦�r^�Cq$*Z.��!���N�G<T8;�"O�"1Љ�~�+�F,~��� ���T�؆��n�l�ǻq���7T��u�n�{�W��bIK��e1�b �o���$|�褢�y�c9��Ps�l��-W���u!"����]�Weϰe�I=ho3��c�GS+�T�� �Ҝo�'�c�=��p�r���wq�x��Ǝ�ʣդ�p��Ʊ,D�s��	��y��Q�!"��n;�E�dj�W�+_�[�n�;Əzվ];W��,7�UL����������CǍ(���i��Ӕ�s���-S3Q�U�ӱm��W�.$zn��߆!R�v>r��1߱����2���m!O(3de,S���4U�|� �]0�7eC%���H������1��q�����)��I�����6�h��aW��m��)E�\>�ADU���^z�z�zuc�l/SQ��s/ ����M.�$aiNd��������w_J�^1�g3���Z�k��K1CLf=ѳ4tVd7�SzNe�VY�J�`YT�i��ʹ@��n�tS�k"h��P�'�O�<u!*������I�D5��u,VT��Z����L����Jh��t�n�Ƶ�X� =bv�g����9pd�ly��!Nt�90z!� 9`��Ħhv�{��tP���?6)�6 �b�fSf|�A8e��c�rD��K��~1�҉�7���};�Y����":>��s���;�^g𱪜��-\U�t:屓Ӥg��Z�sO�h��]�/�q��f��-��̮�d�s���.~�[�FVl����0�������ZIP*���3���s_�B_�k�<�Ii���n[�ZX�ڭ���w 
!Y2�~�/T���vԬ�Z�,5����A��Q�k�.�5A.�Q�?ZZ�S2=�a��(|$e)w֙�����ZP��
�q�ce���)"�B��-���8�B���Ʊ�7�O�7��|h_��C\��KPi\��ޚU�R�'��V8�C��Ѥ��6M ]�	^|�U" �6BC?%��B�{|��*
�n@�q���6{8��Ҹ~'�F���Ki��MSՙ9p�A)y���[z|ԔK�)e��K3�_%*�/}���'�a��@m���9#�FKf(�o(�E��¬�j�J�W���;p�@벑���eEg"�1�Ti�Z����/���DD&8�����8��mtň��*䟀^�]����bd�����ݵ�1,̪���ߐ�1a�w�P�6Iexj_�>�fG����_'ŲX�@���hP���C�� ,d`!�����~�e�U�,��KB%ޣDs��xA[���5{��q�V�}WOU���	T��z����J\I��C�v<���TN�9�F���X�hzS���IF���#�}�ۡsz�kh^4#�5�,�RK�v;�'���f�Fl��Ǯ#k�����'��3��cN~�+�)ց�Z���Gc�V�el��f����(n���hK^�4c�'׽��j�I�� T g
�!���j\�tv/^�OyԋD{n���� �u7f� �?��LS���&M��3<�{���y��o�'�mc���+S�_���N��?�w��p�k^�SK>)�!�A�nH����.����0�XJ!�Tf��.��v��A8?{�U���)�ZU�ё�3�}�Z
ET=���ğ���?�q�1{���uF�f�Y�$'OM����yL��e6��
~�#/�N��)��?�$�Z� �����@C�j�1WLis�e�z�ce1n�?����n��"/�k'�*�)l�<Yom�N��iA��{��`�Nɇ���)E�����+ �$���#�[�s�G�y��d�)�S�0[x�sSC,�)xA��\�Y��0J��B0�g�)H4s��-ϧE���[�cׁ�HN舷�%��e���"�}qT��z:=?�+5U	̍)פ��t;���c5�\�r:�b}[Q���� O����+]B (9��
m,��x��V��y���\d�=U����jeOM��1�����~W�^>��c��
l�0$��mA6�kT0�u�	��:۷�&i�$¥M��d3�̜M�=2)s�7�Џ�����S/�6e{ ��H�u�L�Ɣ������V�2@��;Q�n��5X�+���YD�֤�M�;Gˀ�H�2�����\z�z'AN�O`���cM�p�.L�se�ba ��s����S�&��L�5���$C�������u;�I`ǥ��8Q����Em��N#�����Vn�ߤ8�f�y+���~k�V���v������s��iq���^d��\�#*B)�܋��Ǹyఒ��]�U�.�ֽ�Y���*�_4X^�Y�b�be�i|ڤ��;���������%�ݵ`w�h���Z�V����\  ���%-�y��r1vk�CX���'����yJ��L��&q�>!�4��>�~�.ߡ�?$�>��==���}�r�"U�d������:7�[Y�3K	��};��E�{Q�������$�"���;*мg`��c�"�C#*�������!����/���;�a%s>UKr���	��+P�:�ň|X{6X�q#��#5�2������� �4B�9���K�
�	��o;�ק�Eh(�3��@��.X�d=6w��0q)�^<��,���fzp),ls�� ��p0�I�ot���$Gu�T���U�Ӄ�X����<A��h�6Ǝ�MD��
�$St�G�}��Ӻ�N��%��]��A�7�)��!
�~AD���/1г�F��dL1ٙDr�� ����0i%�+_��$��[Н�����5oM9=?`~�_�I���R�ԡ7�2�a��L)sX�f{-�@����k�ITr1�H�ƴ8����v%���V�u��k{�=���y�Kƻ�H�#�FC��C�"s&���O<f���8����r�N;�P�w�V��t�!��8h群<�2�1�	��}<ͯ� ��l"Ba�EaDk��e�
� >~3�̿���<p&Cs,)��k��!��e�Q��ܷK�oڐ��ЮzRe#�1S0���9��H��	a�`�XC)﮾����Q��c1��	Ufy�MCx�8)���e��Q��K����Z,$���;��Z/�nk���ay3��}5�nK.P��{ʹ�TZ�Q��P��v�i�6�ӆ��,D��!M�Pwd�zy�P9��r��-�%�HnϨ8F1M�Re��~��4�t�Xɽ!`���|v $J^���Q�K�m���=)?p �mϱ�0~��-��4C�p��<Gb����E�4��`ň��1� �!�Z�a�`�ѓ����ĚM]3>�g3�����I� �ʓ��8^=��u�����˶-�s��,��@S��E/�f^%�Z,�N�
���-�T��JEVY2<�xa����N�O�U�
�N�ovO�e.��-c|K�*�޷*}�V���#T��a�SY��f�Ő�����"�&�>3;ʑ#�.���*zkp����^��<�[���g�����q����)Us0�!����/��<�ퟷ�V�t�(\�Ӣ�����gǡ�'�}W��4�߳��J��$�<�X����Gkἓ���k��awG2;1��̤��瘆���}��L��a����
���O$x�Q~Za��}����ѵe2���vG�>�Jl��"��#9f`IRA�D�zU(c(pӊ���ko]|��ׅ�W����U�	y2LL�)�_�鮴�`Q>MPyS!�j�F���K�J���tu9��_��/�|�+�i %�c���7˧�i��&��H�s����8�X
�Me~cYvJ�w��1G����R{)6�I��9�w��g	X.��Ia�,�bQ'9�e�������r�X��K��lǇ�S;Qg��7F����]�mx�����%�h�a����S���u�ậ���O��(�?�/S*�9䫈��rNc�_�k��_bn�g~�*�ks���q����.oGM��@��% �!�Ƃ8%&C�կ/T0#cN}$��(��;0�[��8�i��:D~oܕX�B�!���jJ��h�˛��4ߥ�G��?hW�<-�>�\g�������2�ON��1T$2� Y
<6������kt0�Ma���@�ա�B�L���,e��q�Tn"��'�	�����(�����&҂>^M@f��0k��K�N4�+�g�>N���sCB*>�V�mUY�Ly-�_�(�ֶd)��
Z�ڇ �cLhkG_��U��U	n[�r|�e���WM���B6��M#�a(5k���|�o�Is�Wvk������K�o%�I��*㓬����:�zV�,4fc�������׮�C%
"�,S����nx�^H�Z*��X�ӄh��m,���I.Zp��^X��[
��6D>/ׄd�뿕�,?�W$MU��Wv�!���kM�����V_g���G��ƽ��B]�"��	E��6������|�4�:�,GZ�g���<s��T2��3������ڕ�p)w�V��{�B�舁;�W�[���틃~�zwKʨ�o�'���A��UG���h[Zσ<�
���X�b���Lv�΅�}-
��F����|5e��=tf�ٝh�=Y��Ɯ��rC!u�8Nf�á��U7�;�Csj/di�n���0�?��m��鵛؏�[�g�h�S��ȯ��!����Ԁ����)n��C�j��(w_�Oh���H�	���d,]�&���q%��FC��3���5�� i�d���S��䪞�J�T��#BN�	�#2�-���>|2r�7��I3,o��䘷�\���3b���?c>�����4 �w�0�+����6���7v��u�Z[]�A��R�	����hZ���e@;/E���D����8�}��ӊ�	� �_���<o��
�w^s�yn0VqO�OP@�����8��'~����
�O��Pjt���:�s�͑ˇ[`8��\�Ӆ(�XȅVY0V�`����F���[�9��g	Ї,�Hs���o	�iC���V)���H��SǶ�D��g��j�8%4��7+�#��7/�}��Rι�����k�@�0Q*�g�R���`ӵ�RF�H6�c�(�©{)�6��o6��'R~1�������ʁb�Ɠ�`�]�9x�#HS�U� �/a�L����b���G��%�ll
Q����*�M�ļ�����Q N~�g4X2�"Z� oO1M?�pE85*z�L���-:p�(FS��.�iI�S�1�/4�c�V� ]`Z6�p��J����������[���1J��Mr�4�{�����X'����P���� �&<�Ŝ��@�@��#���?�,"_�I&�Y�oZ���
�"n_����� �uD�!��l�����z^�{�������)3� �疈B��c���o��*��O���Rv�^˻+�����ݸ���F|���g�2.:+�����6x�<E�඲���]�ah�`]�Bf��^��:Z�����1��H���t�Kz��&s�{i���'�#��fB�,�t=� ���@�o�j�?�BB�����8��o$>�(�|2��A��:�D���.�~������hя�)�B*���/D�_�%���3]�`��q�������F���1�b��Bb��%}�2_ �˵mk�6���(&yVx��}x	1�9R4t�_�qHH��&iEӴ��|��ZD�N��.9V���v?�����R@�[_��$�VM����ʣkM�	��Z-<L�c�����a�8��%�(j�P��T.��o�3�����yQJ�m駬;A(���Lh)|Gdk�' M��&��\����37���ĮȐ��6��&E[�@�r��������}�MȀ�%vJd��Q�x:�k��g�R7W�ƀԾ�� 7\]ܯ�T]В �(�؝�$R��t)��� 늗�^��C���!E�]���{�0��fy�1�c�ǱX��N��\k��� e�u��~�!�a�	Q�_3�)�eN�Ϙ2�%�OL�������0��z+���N��*V>�s*�,�-�1�M��O�:�s�\p���ft�Th����i~�"�w�ȴ��I��ű�0k.(�	-&���`eWaTDL�&�]-�J&��&6�D���P��{79�/��b������_���Oki���i_��(}j�qσ���Y �"~'���}�6�\D�`i���ʲ�דg̺�J��C�u{'���DG�M[��*#��q ��LR��r�[iّW�gJ�ܳȏ���'�͠}�d�t���g
�ǡr�T�������G���C"]6}��R0b��F��S:�F�LM����S/��1�)D3T'��$m�6�1��})� ��h���<��9���+?�Sj�	���Ϫ�2����o��9�JOã�@����5]pH��wr�.��"�����}}[cpY;j�ˋa�Z�t��v�G��7��M�w�L�����l޷({�����i�A5�(�2�:��a�$v��'�}͊�";�cw5�'�8�à�"+P��UIp�0����ێ!mc��U`۝{Ƣ�(�G)�u}�Jr亯�ꪱoQ�����c��u��״,��?���F4<T��e�[�q����đ!�����Q��"<J+���.eYS8�CN�ɯ�0����43h]��g5�� �S�l����ruV�hq>�\W�8˚]��͛�1-<���1@G��e���:x� ����x��� b�F�����R{h�n]��1ά ����*�o����x(�1��"037��)V�#�Rr��o��������{������}g��ʍ�L_u8�X�	/��d�\r1�L����7�i��xv��P0,z�o����F0�m�0��h�}:X��$
����eq��Ud�i�Z2H"�
Q���Q��_��GC�o�4n�s�v�{�+ǥ8�o�qDǩ���sN��_����k0@_e\R/M�H30䡏����B(mwx��ɠA\�:�/�@��{]f�����g��u���e�38F�;����L� ��.\	C��C1JZ��jO�$����ט���#:��Ȃ�Ur���r�!n�����Y(�g[Qs��C��_�埐�@��j��5ߗ��F_���}���0��T�����`a���"R�j��7S��-�y"Hݲj�
%Ll�%�VL��5���zܐ��� �����Ga��M#O�P����/�K�W��YԸ�nb�����}�kbg��1,�F�+ʐ�F*��+h�]�>�q���H�L�5y��x)M����>���S�kb��2��ix�@�v�ܸ��n�"�̔ݑ|>�x�e��x�S��S�K�xNS)w ��
�o��	�ŕ���׬f>�%��% 8T��:W�S�to�hh�M�̴����U��|c��{�c�a��=�k�?{<��=����k�5�R���!zRk:�V���S�:]<m�Ҡd�3���u6G�7������X�� 4��iSϹ��K���y�� ��R��*k��	2�Y/�c�R
_BB�hO�0�@�s��Њ5G�7�)	}z|Ӥ35x��X��+���RbGjs�"�2w}��2M,����p��:�}a��+f3 �Rr̴/5M����6�h4n���o�H�O70�ΕX���ԲZ�8[��$�Zѵ�PE���bx�_+����	M\�%�45LF��3��$�zb�g��������m����ox��̄��_��G����$5�;��u��h��U�0����J�y�E�Mt��(ί���&Yr�qw��N�<k@��Λ>���$�b��u {O�����^ˇ{��/&��!�����5"�@����;�Ua�3�UKE�}��݆n���|BB5���*���v�����/;٩�/�m�_h;!�CE� �)I�eG_H��9[����pY��5cS:������jo=�9������4ٻ��=�N�޾�,��(J��V����w����qfZ�ģ}s�u�)~^�\JyM���d�ρA�2�؛\���VᕶI��H�a��H�&b�I0�h�7L�}}���q9}-��@&Ο!��'-�H1ҿ}i�(������M��!�LXi~n3���1���_̑��1�5��=�e
	�ۙ�4��TQ���}�x@�K$J�'�(�D*��
����#�9Kb���X�荥U>ܯp���NZ:bU��qE`��s���C�Ѩ��dM������n:5�k�C����������2�E�7�kLc���v�����l���8�����X���P�2~��[tb��Gbq�����1
��ta�C���E�M�s<�c?���~{Y���AM�D�����k�ca�U� ����� ��r _̉��:�����E�/3RA݆��fZecg�ԃ �S���Ӹ��~�d%�T��1�i�V�I�~8´�?#b�(��(iL�
��:/;�om8较���z")Pk���b�}�j�֛�Ze��m�#���\{Rb!���*mY�I����n9O�l� _��Uͯ���Ϋ�Hp4���P���]l��~N1��J7,4�&���e݈�*�O�����U�Ј�FU&%k��7��T�Y	�S5��9�)kO����沫Q�-�!Q��u��Au�=O���Z�����52$�	��6�:�u�*J �5ź�>�
>�0�!?��IT
��W� ��O'����oUߴ/#�zBU��2�v�MN~x]�b	���+�*�����l�OeLU�S"��V��������5Ѻ|o��`�~^��|p�Υ�G�:徙6Y��瑪b�&͖�s��>}�{�%[�h|����EڝX�d���I�������T!�W��|@��!�
b&{ܰF�R)D�хD1�q����+��UrC�6zH%ǜ�$�ۢ�M�Q7��@�&�~ϣ�^6݉8�,���"ڟ��)� 2\B�1m�H'�N?h��8J;�*Y̍�I�4�)�+r8�+H��{���0rsQ���W�A=j
\�K���R���|χVb>��'���uL�����Y��Dm�+Y,r��L��{�G� -<�eJ^�S�>�)��-�Lqw��.z�Y_w�YJ<8���ؽ�����tc����l��ĕ\-<gL0uٞ{?��so.2�6P�L�3�!���:j�:|�e��[��\�9��q�%�W�h�oL�@�Ƈ��n�u�fX����A��M�J���.B�@�vۄ�]�8���<�$��ߪў��LR�E�7�?�v�B�;%J9n�5��T��k�t�� <2=AƂ`#E�~4���W�T��u1��n�o�����J��ф��P����;Xn-6*E*�;�xx��|]�T+�<K�c��圆t�����BQ�����
�V$�+>j:$f �K����������X�8:'ݡ@=��c&�]-�x��G�"�`N��A��#X����JZО�/��b��Q�ʃa�j1�bܥ��аh)�`�s�B��V�܍p�*��"�ѷ�qD�����b�����%����@�?ܢ��y���ŝ�����н���.[��<&R�"����.�^>eL��M[����Q���$�M���b���V���ØL�wW��k���6㤟�ҀP� ��x9�Gv��[A������F8��(����39�4.M���ʾ��bc��թ"h���t]R�����t�R[�\�/�^M���V��>BwlY���wsO�x�����ur�;ْ*8J�친������B�͉�CqaP
Uf���#WK.Y��/�C;�^E������UP�b���@,��mʆ�ڶ�r��87��%�ns���f�K�)i{�)�Tki�]�s~��
�L#jDAԴB�/���G;%��G��#����Ĕ8vӤ��-��u���L��kZ�q���j�[~2_��`�id�˗JY1F�ދ�Z.uc[T%~)U*�
��O/Ќ�V�E\��i-��D�s���uDgGz��Da������}Yl�~�ˤe Lt��N)r���mߣd ��R�qʆ�qu(�tRk�pL�RzE I��#s �����ȶ^g��x�D$\�O�(9�G�ޝf"��F�̺������� 7�g�=1���XgP�'NX0\�=�c����١�v{�E�!胻jj���R9�G#O��9G�>Bg�K�T�U�]�5-!&� �]
�zY��.
�ށ</�H+[�J���'�2����E�n� ��xKe*AY�o����Ǹ�`!=�<�ݖq�e��N�8��׹�p7J��=�W��{��w�	�W�߲G0�OZX� �g�����&n�y��H��Q?��I6�ŏTJ3��?�#ƥLSby�Re��<���<L�e���s�l�����R�=�R)� h�v�&l��0�1�תb�Vz��=)��X=��aH�@������6�@%:paR���?Z�/y�E�6��#,?�]��8&]��Co�L�jّD&!�R�����m��M$��jSS��PF����|�53�VK1�c��#2q>�v���t�� }�ȖB[Gj�a�~r���pj�%_{g�L�~�����V��<"�V㞄<�����~H͡tpx��~m��I��F�;��szT��8�rɡA>��H߻�|����1�X��/�Dּ������mxg�����ZeU�����q|�����`Hb�]�7ɯ8��������E�Fءz���n>r2c�����5��_�A��e��"]������B?lF�l�z��Sïc\����HHg��P*PgrK��}}wN2j�\�B���Ib�t�HaC�/�&k`w�f��5��;�<30B	5O�y��0�)f]�
A����
�c�{��e�;;8�4��'XհQ4�Q�@��6�!��<�J��7L�̹F �� �ߨ�{�*�z�k��;��.��Y*B	ৎGL&���'S�q��y�	�4�B^<nfN�'�[�^0XV��Yg��Z�@��'Y��(��<p�h��"Y����W�D��6��Jw��*��#�y�0�E�6�w������e�1�E-~f �I��E�4�_,n�ީ��w*�g��=v�<u��e�������=eJ����ȴ�W�e������D�EA A��iE��ո��okY锅�f��|�u�l�o2(�X�C�C>��a0{i9F�N3����'̿"�-o;a��]�$תL����A�V\T@'z�
h<��o�gY�VM��re�]g�Q�Ljd��].��ox�p��#�;9�A
��0%C}�����EwtE��e��*g��,�R���@�
\�y'Z(��zm�[�?���7[�=(�q��teq:a 5'v�[mG�������>��P&��?L��(��oX�p��߳�WBv��J!!����U3��v����zC���׀X�Uִ�Y �&X�|�b��M�a"wN@7�+A���+���NpK� ͗Wh7������`�2ь{��#ꮁ;�Vub�f�2ƫ��^*�!G�ja{�*O�A��a���stɯ1�z��n4��� F��43nb��(j�
y��?fk&�D߬.Q;����iy>w4*�AD�g{��k������LfYPKL��3�TsR�,�]�ή�܄I����r7�>�ɋ��%��y��S�>}�8`"�j7�X8K�h��̢���9i^��~��oh57�3��Ş���o0-H��sz_Gi�[UN�̜�Z1 h������ײ)S�%�<1n��?��Hi~���z��$��(�T�f 4�����/�,$�j�[W�"��IW��/�t#�Pd@EN>x/�-?u�5�f�o�B��K��Aƽ��U�h���0L6*:Y���[Y����ML�1�M^y�`���4�{�3�ɵDGܱ ��E;6�հ��S��l٥�/���P���[e�׻�8�Z5_�:j���Ü�(?M�e_����q�o��>@(�	��E�&�S���ȁ'���Z\�_���<��)��`�+<nTy�hoz!-[�<��O;q�Zq>��5u}�أ�jD�xx���N�<ۚ�~�(SxÎ:Sv/���Oq_�Zp~ ^U�������󂙔�J��W����hY"�,8��͔�>sPP�$�,Յ�P�LQ8���:��o(H������]���C�vn[�Ҏq5���t�d	?��lؘ\�$�ս.�g<�&��ly�R-�{�ˀ�e?m�m_pA��+ƾ���^V�?D��5���$��,F���ZZ�Tꢣʠ�@Ϧ[��5���#��?�kʊ�QCpe�5`5~�Z+[W��Q5e���R��֨��S���릻b��M��y�H�����,��ɯԾu׷-�Ŵ�g���戁r5�L�}����j��-�`���^�G"��dJ�*��~���I�@?i�;�"�N��!�9�M��9�W{����U*\���t��b�7�8�l�o�Į{u#�������
�b@�u`��í�Xͣ'+�8:��{�[��|TL��1�e��Fl�$����3���Q_k�����F�U���q�ϱc�S��d�q�A�N���{KA�X�����d����Z��M@{�P.t�6�^ �"��9�W�r��[G7@�b�o��N��L|.gL���C�;�s-��V����R9P�0tg��i�rQ�b8�	������*g{�J�#@�f�^��JO��OP��5IK�([x�����2�tۓ�B����U�\rYYeVV���Vp[�	̜nk�D{d�@Z���ll���:��5���?K�=���M�ND��
���r��q���k�Jߺ�%�Ì2\�'���ކ�E w�ђ��k`���gID�Ϣ���Fs¹��>�����S���W�&�BFH���'�N��x�^�%@��]��Gs7�يP�:7��b��0��(���N���!���V��(�� �1�����u�����o�p�l��������'<2K���=�T��v(4�}>.E�D�����j�D��;/������o�5���>�.���8��S,J�yÀ��S �K��j
4��'	�ow3��5yh��ͨ�n�2�{�Ge+������ؤ�Τ
_]:�+�E���d&{=��N"�ko��b��W._��Ew&��T�F�o��_*�#�t5�:wKZ9������h��_q����1X2��o����v�,<G�Re8��y��y���v�	/[��w\��p��k( 1��;��lo��1]G�7�M?�/_!��[�{_W���f�ǥ��d��_�+:P���LEq*��՜����F��{|S9p���B,��޼��E!��w�÷��Q3����bn�#$Dֶ
&�1��(O˄���'<K>������]7ɻ��%;��J��vb(���ϠZ@�e���hK�2�6?=�^� ".�H6%^$&ܟ�8|_��!��*֑�~�4wr��_T�F��km�8R�k�
�E��FU(9װ�� f���O )ʥ����?FW�x^J�N��ֻ����D�/�O�,7L	F܍b3 ��F�E�)fYSc7,,f�&���@������W˫ث�ݔ�vX$[�uNc�R��j���(��@�U$o��hia��?�PF1[g-����~Hsp4�m��BE`��xZ����'d���V ����oW�`� �(q�Kk��<1�)��A��J��'L���Զ��YC�.B]�B��n�JX��0��
F�e��Â�WM��Z`�cs4���x��_�I|���� ���A?�(f$�,'G'7��vSLO��w�*C©��kA*|�E���X4E�"���ܧz���8�*�����&g��e/E�Hj���>CR9����k��53ǥ�5u����M%�l9[�ֆ|�Q��"g�k�XRo� �=��Ì���^��Z�
����O��>v���lدsU}��,�"�B�>=s��ܬ�|�DS5�?�&5�C�����^�T�^���n+�o!iU�PV��[����_@_���ܚ����	lg0��*�Tޅ��y����*�F���0����oU�gor��7_�nާd$'M�I*=7�<�۸�{��~�n�B�ɻ ��T�i��͏�p�������}����c�6O�Y�$*��"� ��4���%Ӂ�l7?6a�`�R�6�"��Y§�QW��tyOɡi����Q��-)A��RI5_)[>R5ʌh���M8.��4������Iu~��AY�f�D�o�_[���kJ�~��RpF��lb��[�d�^n�U���PV&q���SP w��"3�{h��FLJ��b%� n���6;����_K��iوð���D6j����gKB��Va 
�z�]aH���^[~�,s��o���LEq㱣�<V�Y����O�N+&���{q�
J��,��ܱ�!������ "���U�{��2�I
��r��M�W��Mq�}��A�f>h�{M� �
��T�~.�̼ �njA�v�9NO�PZ<�a:Fm�-��ݽҦYB>����¨��?�ω���WQN����d�^/ц���i��H���p���ׄ� ��D�-=B}tw9wA�O�i�qD�4�&�T�hvd�e�D`w}����N��L�m}��8�\��p��^��ͫXb�Kq�@WޅجG	���'�u߻l�!y)���=N���$��j�%���԰� �p�V��$@�e�f���5�W��������HG �9�N�z"J��r^3���V�@C#��Ѣ�9P�v�_�v�3��|A�O���(
d��R`�dBR%VAYA�Hk�':&=Ș��9M�2g ���~��>�����m��K�,/@�EZT$X�Zs݂���</��Cz�5w�a�gј����ɱhy�s'ٳ�(���F�����6�~�� ��<CR�����ǹ���V�Z��
ڇC����;����Si^�P=-	�:��tՇ���%�-e&�A7�%�{�/ˌ/�2(��:�+<<0IK��`/����<�Z���DmQ����&N*��.5�P#S@��1d�e���i�R���N4�8ٻ�/��/1mɑ;|{ �C��\�O2��Ų{>Y��{����W�(K��Ǩ���<��I�� �t2���eqX���l?�=RWy
M4d@�:L�6�{ԧê#�N���3Q>���v�hj���BiǭT�;f�s��B3�B�/fg���j��������#�;�R9���4=�kp��Ӽ�
��2���<&�s�_7����cT5�Є��\��[�Y��y�����PV�`�}��b���+[S�4	?L���_���_�$���!�w+r�-����j�(-s�^��,/g៶ϧU[[ؓ����]e ?9��2�����7N�{�EO���p�'+���B��ʢ{v+?ҌgD��k>r} �Ô:��7\~E\�������'r>��Q�p���S%������!:���R[�67{�t����������d�:<�N��ޮ}�
]n-��K�XF�j#I߰n����L��=�	��ԁ��b�Z	���ƍ-!`�L�4Dv��O%�AѦ�l�RE��z�B��7L��=�%JRf`��]��:1�Q���9-qYMLc��p�?���XT�'�踴W�.�_��s�1V�p]�h�]�~C�P��<�J�JJf�C	k��+Ջ�%kVq�$���w۠ٽ����0�������]��eR�ѧ
�-+CsCK[e �&��'7��j������c�,�+x�3��aA�������W+��Ӕt���.=-
��ς}��7)Y���b��}�y�r�Z q�4L͚@V'��-٢@�J�m��!]0/J͠%��9\n�����4(	E��hU�HWeԸ���,�Ո�5}{t��_��7��ť9�X�D��F���22  �}U�³R.uΎ��erӝ����s�_T���l�l��t����3[�W���f0���gX+�K9#ԡ�I����5�F�t��ʀ�T��� =^2��>��
R�+�$�>�5�E����HL^CF�B֑r��{�Q��O���}"k��E7bch��.">�2���"����_>|���1,�q'K��#l��Ž�$L�~o�D����hzMf��J�)\_deU�Y��fZ'<*-���r��a��^�;�4�8��jټ,��]�R*JIJv">��R�\��Ό6����mZz����h��J�V�h�j�C(�W�d�
6�j~�j��B�ɠ����C�R���p.ݑG��~=�Z�R0�)�9�m1�����;���į��@H��\z�Q�"p�!Xj�(u[v@��o!�.U���rd����ci7���L�� +�{�M�s�TKK��"���58�.��E����aJ�>�҅�&U!��P������<!-e<�T_Ng�)�?gh�odU�(袍���00N����0Ɩ5'�ŋӋ.���+SM)�^ۿ��vu�C`�tέ۵��TM,ƧB��	H@�5JKCon����&L[����(��
h5�f�'T^nMqU .�OssX�8[W�A�{m7v����֞R8����z���tlXc��>C�]0�iB�R�Q���.�_=�-[%��pٯ��K$�C�Ր�@���˧��Ç�k�`@�v�� ����H��qǷ�]m�W�.}ﳦ�.��M���Z�m�敿lE�2Y$7�_H���m-i�~n��0*syM���ɻ�vl��F�-p	����p��HVU/�/a³..n��F�;�{
7�a[�YUY��.�P������������=ת��.���۸W��N/�t�y�z*�	R����Ȉ��b�������1y�܏�EA�g�G��dx��'��#[n�^~i���0���)J2��  ݵ$��Aт�K4$��a@�8!֌�S6�=~:q����D�������c��H��h8�2=�}`�b'+	�6�l
D�r��%S-��.{��q��	�]�Z�c�ٿ��&�G�a�5��g}Òs�/�gs�l@�kr���̪N����l�+6��4��T/f��c���  �U�k�++�0L��0Mp���f����I��PR9N�km6.���sD/�'�/�F�#i���	�����h�;P�!�yX�N�=�<��j
<݋mw�����::Z���v�t���5a�s;�X��5���<��#�,^L��XG��Dg�.թT��YK�F
O�W������e�xXo���J}�
��Ko�jyM-n=��M�n�o5F�{h	$܊O���Y36pm�P�T�Xg���r,���|�F���b9,�@�H<��=���^��]Y]!Gx��N������4�:8���X���2��Ma�-y��آ�g��:�h�ح�-<FH�84�89�Q���a԰_a��5\3(W8Ŋ|[��,�I��U2��D	�Ϫ,�r�qR��Y��+�KW��PO>������F�<�"�ո0J�eY&�I~��7�V�1(�m($"��z��X���@�K"0T�Ck�c(�Zd_n2�l���tg�9j�&�==�����?!
�y�g���.��wF��.�F+7]M�ڽ���_� �5�XO�(�Ϋg�d;hx�,�lX"t���L�`3XMeaϲ���P�0��eZ$�����M־��������B%�t/S�ؼ�Mg�~���o-�#ڗY:�{L�v~�Yq��ݙ�&sL�����%*ՠV�&��oV%Aؘ�­Z��Y��H�q\�y�!������v���ŏ�*��,x�F��ZnS��� �����ڄ3_�o���I[�ln������٭��H�D�X)�����,�Ѝ�=�C���!?*��o0�[]5�?6�^.d՚���E�f�!��F
� �/����s�/�M)�6~�

�٧x���-`�&������6i�&`5Z%t���N��3`$c���ۥOz��	���KG�B�݊����9X�&C��W`��c�2��MY�,��	���ݓK1�>NS�+��tϵE�*KSk9��T�>$�QO"s���$�?��'�q�`+��6�F�k!c%��Dj/�~ˎ�T��bw�AX�qJ��`�D�!B����H鷢�FSDz!A�߹H��7�k���PDWS�6��v��A���b>3�SR����wdKM����믊���� �8�aGɝ�M��=�*ê������T�s�=�l9e��c�_NxIv�Y{D�f�uL�{�=����U-(CX��+;4r���_���=%jM���!����A��n47c���X��B%x�!������f��^�2�&������#��;󵫁W�{г������&{xϫ|th�U�a&��%�Z��o���uί��ved��iA��JJ��A��?�;�q�;��ո�c0�UOa�Cئ�3�mMɭ���}Z�SOSML�;��\˞�P佀���[y��0Ռ��A����J<��R��C%E��E3`��J	뙛���H�j1�NC(��4�͐���ަ��^�PJL$�@��;
s繃YT4G?W���af�M�L��%(EKwkǳ@gn�G4�"������Dv(��o���<��]܆��]�T��T�����S�#n�Ȓ{u2���;@nʓB�+4���0����d�5���v��dE��өd*�O#�0@����?S; ��� J��
���*�az%�x����VG��B#��P�Ff��h�����T"0i�
�O9T���no� �D����;r�3��J�z]\A.�)1�wt'��Q���I�w�_�O���}�Y����g����_\����vw��ѥ�6����7�����Jh��يK�A� �����z���q���'9r�Z��vp�@��(v���)�h6h������}�z�l0������SN��e��N<z�g�5mqD/\1h��aHw6��+MI�4 ��@�zfk�?v�fJ���i#|�?���Fg���]�Z�"jc�o3w, ͢�:��Uqk��	{��`C�'��M�9�Oq:��~#%��θ�J�����7��R���JXt�1�����:�<�Q��ݮ�<�	9