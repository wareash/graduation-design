��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|8���e5�I��d8<�⚰�#���!���ҍv/�R �A�0�w�}%>��� Ɉ*OV���|	�zw�ݻ����9y��B�KҕmO���2+$��&��g��c�zة�X�FJ�|.�Cx��Jr� �٬�dF+@~�!_��P1�fF�3Dk,��BX��
���r�P�K����M�N�X�H���� J���lJ�Z�|����K|�&��?��_?B^@�L�U�tK���:/���tVeu�3a�m����hx����/8zm��_XhxBzM&^��M��k��;,�>��עۿi�����v��Ux��%�-�W���N��_^UDަ�h�%W��C �Z'3◩���B��6)�㼆��hl+L}&+������54����mq�@}�ն��Xg�]��0��˹�Ĕ�N�LPv`�R#���'_�ǩ��'י�^��QgIA�ƕ���u������V�"���IrI��)�tB�4���Bk;�C�e3�
"�)k>�#�:^ô����b��.�8S����Q��+��G��#�]�$֛�ʩ%I~��clW�������wQ�"���LYIlH,/ ��,�hVd�.��A�0+�?��ZIG^��u8�2~��_�qوR��ǡ�3��%y�NܣF��iAo��/�{r;�(�>e���=q��a�������S��?��)a�I��;9�����1'�
��M��ިl`� �`�x���L�L i�쨫Aw�e>�'(Á��k{��hBE&B��a&�o@w�$aNwu��T@�w��Ul
|g�1���p&nkד#@���/���2T��$�1	�v��'+��i�J4�7{\8�R�:��ISz= ����t3�eA��C���8~��T�=hQ.�n�\���cpT�R��`�H� Q�QB�j�B��� �l�)w'Q��±�c���`z�A�3?L~�a��z��ao�P�C�����D��4gk�N�`�4���I}$+�֖3x�}�1���:��%��r��!E,��+
����ubhs��!���A?P�c!F��0�N�2�lO�d̴�|	}$�مPŢ&F��YF���(髟����5^6��U�&g)�__*��f=�Z��,�0I�Ǩ*WN���h��>)p�&�}��f�a�UH�}��q��4%���Q�o�6��Ҏ�}��IQ,��h+� 2�RgXY���|��Z�Kq�����֍\yE9���ܱ��S`7]IOWE`t2�����1����8�à��gD �Ze�'�dlgܣ��O	\�N��֥����n�HP"�l5ڔ��r���fHx�����w�xE<�;hK�6���~�	Z�u1��ͧR��{�x゠P���r�i^�,�g���J�Z����ɯ�k+C����	�Y��.ɿ�D	�eP�8��W]0�;fv�G��rD�]��R�K���!��pM�:� ���4�u�ڪ��H��#)}\�Q�ƺ����H��5 {�s��m�ũ�H[8��'A��m��H�9�����Y7���Pc�m���K-�B�:�w6{�	��4���ED��iXᇦƸ��h��)�r�:��⤲�'M�7H��v�?4��F%/J<����,�P�d�� 
����݁�wf���D��G�iiD�nW��O�S���ꞻ�b��Ps2� � �&��$�3R��n�!��Ь��zh5y�َPL�GT�:	��8fi_�v\3�j�����j�9�2;c��]`
'�%�}w;��5�k�2���X>?7��_�����B��lv���c�\<rA�i������f$�����q� t���+������v2���򼠭�Oу7�#�E �.�QBK����S� <�p���d��1����3b�6ĒT�j�
Ea����.��3�<�ԃ 9��{�(������H�>�ZF>��
�KW�3����PnZy��ЗB��/f뼑}�V�O_�ɍ�Һ2�u���hNwxV�:���B�m��#'��$����MҜ����}g�׀��n��3
'U})?�ܩ��K�{���v��EW�,��"Tx,n���ܻI��N����� �&�=2T<8���+�4C�mԓ���{_ш�{M�u��)�Yv�� �c�����&��!y�ͽ��MkOǉӊ	��nW�I&�$!�3��<���D��jt�d��!�QI��3�7b�������H%/�BR�q�N�ا�/�^�/>���3;	h�u��@�����
���nau9��p�s��jP���/Rf�Ggbڱo�!o��+y��3�8�1�L���4l���?�P���0*E4�i@��z�oB]��[?le�H�&��OP}�jr��l7B�ϑXy��{������{�
��$�Q"ܛ�F2����r�2,�ƿci��������?��K
�ͥ�	?�	�����W�������٭�oa!�s�0	|��ɓ�O�a������T�[��ykZ��q$Ln��R&c��h�c�ϋ�)��� �|4�4:�g^�M�� �O�3�]TlTojK%t!K�V���T����������[T,Ԍa �\��l)�qe^�e5����+es-s+�O��j�,��q�#D�>��f	��|������UE�M{�|���R�G��@g�n�esn�6猝�����⴮�¹��'�1D&;�O��e�g �4�@|�¾sj��\�����N+hAt�;:^[>�L��ZL��RXƨ�������<���,yG$̳5���FhԎث�ʏ�@�*��^����B5D���pUFo�[�K1Dc��y��Us�菝'B�r�J�t��`&��:�Ye��\UD��������&���0��X�>ܙ_7{�懂M:��h��ב�SLi`{ =[�č�����PחbjU!<���U�uY�$p.��,�HU�%��f����B^5jI��ʽԅ�t����������Q35U�/e��i��x��K*�권��eN��m?5�L�ʿ�z*LB�%�^$,�a�=�ř�8���������FiȊ>J�%s�Q+���H	���12�U�г���ȭ�e�u�@V�)c2W����*y����]�"�i��= �:"�����8��m�ڇ�y��p��.�6sk�wȤ���[F�B��P����K�������-ٰ�j�5��Tb�+�f�Q����� ���vb/F�g�Bd�7B���M�P��q|ZjӒ��H�5hC�`�1 ��1Z_87Y��^�ye8٫�͑C���-i
P�$����ǽF�x���R�=G7 ;{9��tG���U0zd��E�;�v��9�����wMnD����\���Z�S葀���rv���&�,�בE��=��R�ΡV�x�[s(�v��E�(`�r		��Id}ٜ�Hj�đ�a�zlѱL���J�q�X�%++��j1���V��/6�~�5�1�d|�YVJ9=m�v��'ya�nmI%7�D���j)�`���D����J�3=Ƀ��X��gq�{�T��i�ZA��B�Z�����b�U<��Kz_T8���,�͂��sDo��^޼�[g����^{ڲ<�V� #n���
}��+:{��m�2�̽tϊ��F�O�y4�����E�D�-�A�5a���QZ��VB' D���]���s!��,6�A,�\ł����A�7@��)jS��[���aSiO:꩜5T*�
�lHgR��� �{ؙ-:z:\�nډ1�p��~.�0*���I���x]���;�_N��:Q;���5�|w�i&?���ԫ�N�}y�%��绒U��ј��焯r�epED��9q����!p���%3����,��Qd���(H����Ws9��O^���{x�9 �P��إ�gE��E��i���C��E�!�`�LݏXby� �M:N��3�A1�sG���'�n�#d)��q��=6X�����1LC�('A�R��5�0����R?5k�Y�JE�2�w���%W��NF��^e�w���ٔlA��,��&{KW	%�|f{6�a��uz��eGƢ\��6t,�����R�t[��;8*2	���G
��4�I�������70�yF�Ef��]�4� ]W���Ӥm��RN�`��ѝ���EAx�V�2�R�H�Ǖ:FA�dz`�?"�/.Aa�]װ��U���E����*t>�������>�	J\йᯎ#�ٖ�e�R��`W�>l/!n�eYi������N��(����O�Z�`���H�2�U/�@u|��uv^���|CAN�#zOR����.����.��y�.S�'v��$3%��.i�;��V�8��8b��bޤ[�3v�M3�2�U�����1�S*�O���dN�&��ad��䶵`�^0��>�+J�I����m�DX�?
O���S=`��R,-`��Jk(�����$p@�H>%��-�έ�e���b��˥�e��z\&���f?ŔR�/�	�5ko��*��O�:�W�⯅�⇬f�@Ж!i���,�4u
*o�7�	ŧ֔��!�KP�Sf?^�D	�7�*�w2� $0���@�h_��7WG�!�߿(���q���JN��a���m��.��݂���x���&\�P���T��|��	u� ���S-Y1�V��n4h��t���!��xe�RZ����Z���s���BB��m,�oc|�h��Vw]�����䀟R�� 8�]��.I1/M���(T�%X�t�\������0?�@�c4�{Z���i��\�L�u���a�tn*9�TQ��Q^g#+�G��a��M��:4g@h�ɔ\#)h%����e�ޣ�����Εmř����m�c��]���g�dݻF��E@&��eU�p׊�n�\P=�+_���L9���)���n��������ɴI��G1�>�,�?1�v庍"��ք)ިq/�?Z��6��Iq#�=�bR�HY�J�F=$m{�R<�� .�y� YWK�r.�<Y;�GD��xԇsķ&䠹�s�B�N�}u�[ηd������=���W2�wQ��.b���P�s�;���e�q�_w&��;f^�~�
��ٱ{Q/� #Y��-x�˱�pc�'��W�Hqt�Kv��I'�R�R����#�|u فtw	�����
�mCd"�\BI�9 �4T�0����<A���S��ѷ��H��|����������� ���k�e2��q16N��ZGW8Az`{��k9	`ʸh��J�0_sܫx�$y�x?�4��Ť�+�S�����	���#j�Y���/m0�r���S�oxUv4P�̵��D$f�k۽��(�x�0��}�2Z����֖]\_�_��V�����}��A���GD�N�fc�s�D��z-�¼�~瘃<Gj #D2�<f�[i����>�n�B��~�qժb۬O�@��	��`p��`�. L�%��H�VH[.�2Al��f-w��l���=2�1\R� E�xNjER�.������̐t���&��,ϰ/&�.��0gUlwA�X���}`��{�^as�9�*7�y�-�O�B�M<��T�9"Cs�Q�Ύ;�_�	.<D���S�Wi��ۉQ+���B7/J����z>����@W��E=��z�Z�FI��u��y����#����7���U����ÊM`yp.�Ȗ����'a�8������V���5�I����]�O�����Af�:׻���Y�r���ɍ9Lu��t����0L���g�����G��ߚ|4�����%]���b�[>0���Bi��h�<^�>}3h���3�x��=��t���b�2PI����4XU����Z�%�Y�=�s��%&NLiDk+�A�{��������Y1�j���#iY�SlU�t�C�K���@O/ʬ��F?���p�]f�bARC�5@N�eQ�g�����(�Ma���S��ߠA�d��,��M��v(���{Np�(�Wj r�8ώ~�#�K*)���Ds��ңC��6@�%��h���o��0x��AM/�j�Y�x�5}�
,ߧw,뎏>dz�n�'��ܝ:ꖐ�CYʜ���Į,��C��փo�����{�]+pJD�%�m�]쵺�^�u�L�~6�a;Dj��fF
H
����AP�� d�պ(Rk�����'��p3�"0)��Dˇ�l��X\�g�vu%�-L?n�spQ2b�sx���hYb�b=�0\��G��Uӣ��#:�����}�)p��U{����G)%��d^�`������#0t���o�����L!����FI�����*�k]�5���GB[��&�gV�ԝ�)�8Aj��.5�U���:�3K��y#7�+Wg)���vfT���e�g�.�?ḳ�1Ζ�T����}^�P���^?�Ad��H��zbj�@e����QRFGxV1�w]���C�1�=d�œ&�-öxk�����������P�H�'8��V}(]Ik��E%�����F���0O�@d:�:T;�B��c�{V?�Sw�^'�)e��t���("'U�Z��s���=�V�̟;��`D_O�Q"��9>PJ�jJ��*�	�\ʊ  נG�����l�zk��F�g���ݼ���.�}�e-���xZ�?3UE���xXG��>#�h`h����4��nٍo1�~ZXo�錋��YO�#,���>�?��ä�X斸���y�=}K~�ָ���0$��J�3��������Q~��ix{D�L���y�����c.tQQ�D\Wg�,߂��͟�j[��϶��a>�y�W_�Ȥr����Y��*�S;H{1��}CHmiU�ݒ� �>�;��SQG�B� �D��!���K|�ol��Lb6%��j��m2�ޱ?����7��(��|-�Ʃ��SI	lQO"�a�� ���mjYODEm�jz�ZP��N8��%���\���ƽkoY٦�g2kt�cO ��wW�Js���Ǉy����]�2�e,��I��:�I!*������U��ȯ�B	����u���A�Za�Ε� �|�����,^26�q5¼6�h�"�a{�SpC������I����7���"KۤQ��|]����`�o~��nW�L��ś�@`��r�xq��'�z⁠w�S���G{�q����(�3�kHP������v���+&&�qz���zv��8��o_�M Sǐ��;lf���i���
�&��1��S&�&z~`��$uĄ$��T���V�N�M�7�$���C�o,'{I�	p��$�٢6�,���y��-�{O,Ɩ��=�oe�i8^+��%��8�H�� %��Yr
<�^�&}$Y\A��!�5���O������
�C-7N���=�f�� l=!���l��d�m\�]���N}�9���>#6�W$Lo�V�r�T���ƒ��I���Љ�j�S\� �6�c���� u���a�s�7���ưB�"���t$�`D|�N��5?�'�v�?���0��°�-m�� �i�d���A$m�>�Z:�w��>��͑W�����v-������]����89�~�^���}�֝�s>֚�86_����~����O��[���tZH���'��J#�\����R��t`o�f^�����u�Y4�t;�����/���X�;��(g�Ot^N��4|�ӻD������gv��7_��lY�W�p�G_�GF�˿n�e�&(\x|�'3���;�K��X �w�m'X
����6�c��y��LI\kԿ��ؔ��T�!�Kt�z�ߩ�_�K��}	�	��+[�8�@�+��(+��By�$�]���2�bAQ��at_vo�ߑ����dpe���;������R�&l���.�U�+@_؂H HE����L�6����������h�g��&���r(��Z��o��I�b�\�E�G�m�t���S�P����F<֓Oܳ������}`�A�&L)�^$�4V���=씂L}sJl6��~��K�?��c�&�`���6z_��xdd��\_4�gT��*���Jv���?#�/]� i���y	�p�jF�N��=*%[󻜱����2Z�\&�h��⧏Y=�~�b�!��L��6�^�D��N��ᄗ��8�"ja��}���� b�k�Iz�=3�:;��b�G�e�a}��<�-6C�V����8-�مX��f�{F��� �b����`t6���5�̔lI6���=�Hn^7���)Ю^�հz���{j�M��qz�Cw��X#�R��H���l�����CF���3W��:��\F]jN�E��y)F>8E�=��K/zܸ@��l� +�c��nX��b;�hKK"�|���G%y!4��m��ɡ��@��e�I�����S�n2���T�g�t$��7�c�aN|󭷁y��u	k�76�S�⇰�9�Ѝ�S��G�QS IFv(�x��͹���v��A�&���L��� 8���.Kn�7�c�!�c�ݞ��hq�*L@�I��t��ؽ" Z���T�Q$;O���2b����Tm2g������4�<n]]P�h�)�>|�u|6j�B���R37Wm�>|hp��O�HS����^��p\����B��WkTJP�f/��rŐ{�JS#�HC�!���u���jd��K������?�a��i��,ܒd��Ѯ,��q� ҩ�S��@LPd��� �v/�.�p�>�J��c)	Ec�.��oX�:i��r]�`���}G�q�f���-&�nCifEA9�jې���ޏ�/k�m��.��6v�.-"���2���n�7���Mu�+�q��a��s�nS�|�si"������5��6I�6'}�� ���9�<�젡�"ٝIU���g��0UW���,�Ѷ~)�N�3�x���ρ���=�9cҠ0�v^��'��ҽc
;�x�������iPQ��e�K�ށ�[L^Dڽ˭7M� 'f�2��.�L3��ۂ_5����ݝ\�JQ女�?�Kw�]�ݤI�K���b�?����\��8D��ޖd�u|����.���{�H�M3/����N��`���6�i��R9��^w5��o�XԠ��9�2��ob_͝�=�觌y��ڄ��t%��V%\P�hpG�
=�*^�@�����	U�|5	�u.�p�/�4�Q-��,��BҰ��8�Pn�c/2c�������� YD�p5>|>_+�\��b���ƥp����`������7RI�N�V�me�<@M�Æ��m'�$ G���%\X��UC4�]��q����Pa|��r>[C�&L@_�������Ѩ�-ڢ��Pѵ]�[�̴��I�Wi0��q�i�o�^�rC���_®���gw.� ���VZèW/ȳ��Խ5����C��� <���u�:�81�(���S9�*&=p��kq��-m������0Ҩ��oͧ �� � ґD�]��H�A=��@r������Y�I�E��LpK�v
��������q��	�Ts�An��.Q&�+R7 �#�E8��;C��9������
���d@�V)S��:9���\0eVs��a\Bq>�Q����gB����I�J�)@J��	e�d�v+l��'s4���q�ԮjX\���J�@��b�[��S�u�;q~�}�*���OK#�T��I�ϔ|�p�=>�Rᦖ!w����o��M:�}}���~[�\�B�����$s�c�KEl�ѽ�e�X4P�M�Og؟I��t�K9��gU�S�I����,��?�3w������Z^7�P�p���{���֒��&DZ�&(_;����p�ȕY_R	u��қgP�\	�m���������s��D�*aƼ��P�sxOԋl�����X�\��
x���13�-C��6vR&����l��|i|5�84�1:]O��5�C�:JwΑ�ʹ�ɒ�M�P �8�/�6d��s_-�%R�{�U��}�]א��i�^�3��0Q��l%��!��GT�b��]I.[�c�5�?����`Nm3��S�����mK�=?贃��ָ��iCv��0���ŝ=YQ��i$
~�!/�V��;�Tca2#�P��y�ы���}B�m�C��^Ҋ�W��h2)�[�-/���?��Vj��(���,��~Ȝ����ݹ�~'A|j�"�#B{]��R�/¬-0P)E�O
�AajT���1=6lFR�#��!��8��A��Q%����=D���Mg�E	��XVy��9 �u�P' q6'���l�
��7�JI9o��.`R�����SE�1g�t_V@X�A�)pv�h޸���+a�U����?�\�T-K��;�+��l ��E��܆(��4 S{�������	b�=��������"��%>�i�F�q]b�FJ������pHw5�D�JU�_T@�[�<�����}Z_D7�vV@P���̱� 2�L�dJB�����e�|�NMi�M��%���ӗ��t�Q����s !���|d+ơ������-�Ŕ�wM�I�6T2Iw����'\��F��]��4���\C��~�F��ۑ���Ş���Nf�|���R���E�h�@8d"l�b�<[WA� C]�^#��2=4LG}9dlMn�s=��hk��')���11�I���orJ��2��f��	j�N���h�Vg	ٕ9��ij�Se�RP����R����ё��-O,�K�}�t�D�V�J�UO��
!�θe#\�6��+u�d�l�=���8<>m��C?w��ke�����h�L�:;��4���!�6}��r�|��o��g��~��J�W���	@�t�#�Rv��\nY��=�-f0"�׾�3w!�D�5�S���(��Ė�5���^_����(�*妥7�����*_���*��C�xx��G����dȤ�u�*>'=��q�c�D�$f/s���4&0�;�R�(�"��֋0b�v�΢4��Q	�uB	qj�(��G|��i��$[Ȟ��"��! �:����pҥ!_ �	���Qk68������{��;��"g�o6}���ȫ��d�;��=��s�Q����@�ndq��JǴ�i�"Z㫪�en��ǉ��J�)A���ߡ2N�|�Wv�eɾG��3U�[ë�B��w�[(f�=�������M'
��+ )��T"���E������P!m	�JF,��t���)zA�����A�����=/a��m���(w\���h�R�s��
��"Ç,�i.������1z�O��o�Li
萌�]�V$Jo�#7������=�-���@ϡ�?��tx�� �:����Ʀ�8���-P���/��G���'��y3��!�L�X���A��/�t�yA9��ixTp��D�Z9���$�?�p�k���$7P��D�ԥQP"\�&�Ҕn[w���@W7m�}zn��-��@xP�eP�����]�%[b��ͨ�o	���2C�?�W�?y�邕ժn�R��m����qf��뾡�A�t�����o��a>�Ԣ2]�e�%�y��� �լ��6`F�7)]'0Y$O���������֯��v���.ܰ�E9�����!�SQk~)*=��Fa�����S�p�h�����?���_5@ �C�jS�\�C�ː�k[11��l����7����<
l`�����a�y�Ě�Z��i��}ڰ��t�-b#��j��UFc���\!�sa$�uIM�ހ�JeD�=h;�r*X�	H�:���MiЙ���_�{N��H�����`�MZB�:�|I�FSXE�ן�L��W�ө��(D-fB���8��8q�5QiU��p]�Ϯ"\��ұ����	x��D���G�k��v(��ә��k@=>��7�& O�R��w�Xx�
��K*�	 ⠹�ӄ�m���P�����\���Q4�CDG	ߝ���Ǝ���{f��U^�c;��<d�۱�����7���?͖����D���?cǎ5��:f��n����4��Hg^���H�"?3���~Qp\��؟Y-�bM�r�5biq.���]�{�4�1O�#�.h�]�����0�V(ji��Jќ݉9��\�d�O��p�V��$�k�5{vXT�6s�#s�6ר�<�/qN��"<���]�c�ac�}�%��ލw�WO5.�+�#�����4&D�]2歱	%���;oϢ���f�DAw��U�9X5��ng57�	"���:
�hȧ%����}7����ky7�U3��N�(5�,��_��0׫�$o�ӓp�䉪ɐ�k����x]>���k�l��Zp���M��P���:�O[��ɣ�Щ8�tVq���c~f�y��@7�cč���L�2͒x�f���w��f�z�"�f�	c��r���[^/�9��ӝD;��6�}����j�|v�>��?�+�_�L�L�D�)'5�-y�,t�����]���(3q�(�b?�9n����eB��F��=(����1�T����V�9&c"����pax]w/_<K0U��/7M-.�x5�ᜲ�In;��yRW�}&qo��
�Ye�Y�|�`5]��i�����UW�.�Bv�<=����l��S �^�KncH2�q���f� Ϳ�&�rN�7�	�ڞ!���=itCawݏehII����֞ĥ�����D���g�h+�:�  �\D���!��קs���Ls�:�l� �=�A�C;�Gb�p��	Zk��?��/���Q���
k|�O�'�o��堾�+Nf�����8��E�������Ď�����[�qL4�Z4��ou��}~Y֤����@e��̞�x�wV�VXr9�YW�T\�8���Oe��˜H���֨��C�s��eՈ��gͯ���B�l?v#�1����B�ii�(�E?v���sȩ�P]|����y���V �2��Z��z��^E�p�M�a���?���wq��s��>7"��)���qǤD�og�.�Y�%��7��x3[����Ѥ^GH��֕"LfŅ��Ǽ��-�Jf��QCOj\G�`9��֞p0;���C=М��=��Ce��E�$^g��D_C��,��l�ِ?�e}-N DbHJL�u���T?�#it��]��s�9�dP�c^+$�ꊷP< �"�3ea�i�E�+�I}2�x_Y��RHl�8べfW�w�!1��|N���M�쇤�{i.	iZnD�P�W�տ
��-/�Pf9i�9M�Hi"���8�c���+4s�	�MW傉ڻ3!7����ǁ�<��э���nj������������h+��lw��1����Fl��7j}�i�?��@�L�	6z+)Oq��O���� {g�B�U����T���[JCX�I�F
+kA d��aڒU�qЄ�PI3@�i�'��|ǝ�2j���4�cK�_И�{��@A8�f�<8��L���.^ _�+t+�v�J{Я�#���]���[�v�Ҡ����wْM��xͥ��5�����L7��{����V�>WѤ,G�Hb�Vi�7[�-5�����p��b�<�{P_3���@7I�>Lc�Õ�=y�
�K���� � �uԋ$�U�'�)�E�l-���BG��9x65��2s������N�WQD�=C� �Z�BQ�n��ҊQ\��y�y�����%ä	d63���`���g�l����� ����_3�.��9��+�3\�p\��"�.�n\���
��BXn�03������Tf�FK�Z�ɶ+ӕ[����i��+�� 	S�����Dڲ.������DF"%�vW�a-� �c\�A�Zv��/��\��\�E���ʕ����_F���_g�����x6�4e-\i���_4�	:ŉ��y���ľ�:�a��%�|�h7��S AhSBK��%��̃���|��2Բ��}�&��Fl{�,�S�0����q�n��Uc��
� �z�3S�G �5��
�I�ܒAs�;e7+���쳅�<	�_xP�o��w�����/��*>�a�$��N�P(g7���q�BN��7��@�(}��K�廏�p��^�мC����U�<�M���K=�����FP<��w<��;Xop�Z'th�ɏ��"w�z�5&�<�[ul��m]"�4c�0��		�(����ga�Bk���+�@�B��.�� � z5 ���Z�1Ž����c�-�_��8��5�����%�9�w^$m�I���c}/�;1Z6�?�E�[�7,�'L/�k��;7+ӄ�|U��7v�:!�.��KL��O��[̑���Ѝ��3�\��x&��Q9	��]A]��gAjO�+*Һ��7	:%^�7������
�*�Z;�/�ʂ}წ��	����5������u���L��>F;>�a�����T��_2�	r��Chi�jhoA�n�E�[s��@~1@Qy�N�6�����d �M�c�3��IO lY��^0I��ጧ2T�J����w��2p�&Ƴ7D��A��X�h��Tv2��\��X��a
��%�C�04��5%?��e�
$`Y#T/��3F_�����:�vJ��2�����S�?��h�.	���sr��{��'��{,؍�����E�g�i����,7d3��t�x~9H�W;�M|�2'�Ծat`�r(�� <ys�ؑ���)��R�[��x�7S�,].?�o��{7��	�9\�ݻ��o�D>\��I��3qh��\���m!��b	��HC�ۢ �Mm���,&8��3 �-=�b}œi���}6�q5�R���0n��p��©~CY���Q7�o.��ێE�g�f���T~����Z��:ΨdN��X�
�Ob ͫ�@\@ӑ�%� z!�B48!V?��}�����'�H5S��,Z�o��jL/$Tp�������*�>�b�1�9yH�%�^�i 8�����
��*�rɠ]<~fp_}*�׶�Iv<�2�14F�Q��,{���l�E����ef��T��F��%�����΂�B�P�1��������RV}�]��V���~��
g!��J��~�>h!��e�A#�p�8��XO�ǡ}�E�~9GP�o/�
���?���Ŕ���| �t�5&��"q�ټ%�X�m�́V�_8�W���h��ی`~GJ^����ܟ�Lj�&�Z$at���5�kL{��}`C8(��E_״IX,W�'�*�����bbkBQ����I0�t_u��8iN�_��9nrx �A����07ӻT� +�����l"4u��=H�%v�)B�����YW�(�7Y4��������~R�e�XU]��;�{��Łx mg{��bBB�!~�Cd�a1hL3f/{��N�6Ws�ԡ����\5�&o 	t���5~P�D���1G�g�HV�oy;���|��#���V�<���M��e��{�$��w7aԅL=�>�<JM��ꄊ���sn˸���M�*�D�JH^�
S`Y��\��~z�Pi��1)�4�w2��R����LN��h��9Jk3ͳ5�VWc�<��礩�5�V���]���,��Y��ޚ `�c3+:������Rz���b�KhǾ��TD�K# %��$|jE���D_9���%D^m7���8+��%W~,V�܌&�N�k���h��dgx^�B!�e��-�~�k/�/QX���$a�ۙi&���@Ml�H�ҭᵻ'�{i<�34�P�sv�b�+[�9�4��o�4P�[4
��><q�@��b�Y%`������]�/uqej�<���/;�ڠT!-F������%n�sC��*����{�S)�;+O�R5���m��y�ߔ�ٟ��&����ą��)U!�S�����������:�S��:a���؈��'+��#<�{7�F_��r�|`��6HMrob�qG�U1�_��5����7�Z�����G#�!X�A(Z\�Z;u�(~��N�����u��������C�Vb޾i
uov���c��/	B��؏��#���L�j@!��D4fmɇ�	�����p��K�k����-��mT���B���/�X�ÛS��j❘��U��?��:��^43#��q�Q;�;�ZYcO���~ֱd�-m���cS�^T�/q;M�\ی�vs�fUg�x�/!�|c�6��G�h�Dj�T�
�����~���?#^l��F�5�۞��=�4�}�lQ��
8&���_$�{>�y)&lD�%`�V6H�a��{�b���L@�r�V��BM�qMZnP���N�x�'���kv[��n���&.-�8�w�Vff�0���v�>i��w-�ѣ<��g*�Y��쵎籃M���W���.�ś�ӷ�'�H��|>rW
	%�F*�
⯝q��[���P'��'W󋹼ߜ\�$�$hߔ2���}'ٲW����v5U��A�C�xka�m�������SP�@���P�� ���%G}���`�< !��fk�;� ��'"�'����1�)��k� �[<��&Em�Ǔ��R('v�s�C�a����%ֻ���1�x�$��;M�+� w�#�~�+\o)o���:�$�����&�vrxz���S'�[��̸���lP=
X*������0
�z�a��I�Hq�nH������rj$#����
:A�.:��PuUa�l�q����
@��ۖ'ݹ����]0S���Tq��^ �������h��8�΀����!c\��}t�#7'�/圬���"�4���p�Xo4���v\�f;��1���u�P��=��>w�c����k����c��L�lu^RRg|��v��b�n���{ll���uCSs����o2�%�z�]�R7v�9��:TS?�H�:F"Zk�7V���;(<ˆ]ˠ'��,�ƨp�Ji���>��uCZ�G_��/�4�F>Hj�4E�/_�b�(@�����0��	%�yµE��UL�l1�RoJ��V��yr��B�tnt=uoŊp� '"���F�?r[:��@�!�:٭������r�!��>�Ǟpd��6@v��o#N��9� ���;�m�<��bR��}n�Q�X_rٜ�Ӯ�)���$0��X��X*&�Ǟ�qYJ���0� ��!�q)⵭��,l	_��.�)�{���9�5��c }�$G��3����]E��f��~\a�U��-꣍2��r���~�h3�����V���{kX��b����`��<����C��<����cAY`]�5�u&z�M��-����e�'��[6�Q�kEbNzib�ת�\(ۀ�?�I�j�&-��} �5r�L�w5��8ͮ��g+�Õcݜ��.ezY��kf����51<\eh�2xYڇU�)��e[!�k�ٮr�1=8�(���=�Z;�xT�'�c�&2��d%�����Cũ������b2�%����D��0!{�(���pE2����d������Mw��פ|{�������g"@�M�@�C>h#3..�5��ƱS�7�x�Z�%�^R"f*N���,GJz�S{	�]��ږB�m
T��<3A�:}��Pu�R/ˮõ����xQ/���/�˸�l�TBz�|!/W��Yބ�֑��cT֭b�;���Pȩ�_��b`.���|e�P�S�6�7�ea��\�����v�����}��+b�JTܥAxB�V��%�r��Y g�T��͠�����u>f	XB����h�X�"[�q��ՌV�AϸK�A<X����EenaJ�ӓޜin:{�5�i��;U�h���Dm�Ng4����T�=EHʁǌ#�%���g��c]�}RⲀl��4?���E=�^U�It����<y�$53%R�P.�x�7O��:�C��ȸ��`�����N�z21�#������X���}���.�b]���󌦂D�̓Z��'�#�6��ҵW�YI<����
�5DR�5˦-
^5�o*g�]��D�)Z���Q�=A�A7��5f��QdsIY���ܚ��4
ͺvy��(��Kj�
L`݉�����yx�����9��!�6~K�x�I��-����iV�U��f�靭�j	��'��;�{��4+���C�b�����H�+91XXv*G~�?��5�u�(��c�0�򫁼sKr�2�����K,A���`G���s��|������Q�(�d{]�t�нp?W�n�|����ޅrj�-���|C�F�'a��\�V�Y9�$�-{�`xN�0�;�^�D��&ſq�̻9F��L �Ew2���);����J���&�+ޑ���_%%��=)F�5�6��ΆA���!ϭg5����q�,�ִ�Zb�
_��j�$œ�iHn�Y�	���"\'��%w�*A4L
��*lg�$Q2].�EVv�q�s,��90�T���{�0�aw4n:
6��,��w�X2�[��ʫ@x�!!��8o����y=��e �c-BI=A^:��И��2ǹX0�͚���D��J�F����ଇ�@Rt/o����j}V#�i8Soœ���2{#mq� ��5H�|�w_�0H��J���(�C}X�iɰ2����c���"��Cf�s���|��6��sw�N�M���]/F��Bh���p��ٟ ^���]����
sM�_�(�6<38��'l6��s�V�~Lദ_���Wҧ/��¶$xs-c�Q���v���<���Ea��1�7�hʏ��ᅣ�b���!n���h�iVHK�X�.ֆ���`鶲 �b��$)VᲲ��4H��Xu�ސpXA���c�_�a�H;�@I�L�B$���EkwCܵ��ql١@DVB�I��'��I����PAⷵ:�2��ɨ�h�.2["���=tE�{#�k�����3�9]�+�cn[�YCJ�n[���ԿX]���� @��U�X�DBG��5�@h��a��k7W�����\��in7����X�Q=C��0f��nMF��`^�yu���F��,,�f-N� �_����|�ƭ���J@���wF��m�.{>���J/V�
@>s2��0�ĩ�%��An���Y��K�8\5#M��P�,'o��>�\���tOc$����^s#����>;+���qY�?�*c�Vad��Kex!ݙf�Տ����;0On�`�i^��a��-���(��:��W2��ឌ�����\��R�����4����d���eS�`�x��@Zμ�y�ݤ����}�6Ao~����Cә�<�q��9�%pEOd�	��ԗ�b��l�~(�|XV2���{%�k8E_QeP(PWv�D���OQ٦v��ŋN{{�
)]8�<��p'ˠ^C�>\{r�S�z���w�~I�f�:��?D��l�����e4��wC�2nFFh�Բ����Kl����_(�Ҥ�v.��KM�@S�$|��,0?3��zjk57���/f̙��r����/Tws_3�� v��JD>)�fU�׷~��#sR���s�������щ��ߘ��j��\���3d���cܢY� Y=f��F&�S��?�hbPũ�Š����T�Ϗa8���jo����Xb��"��	� h
����ݍ%!���K�?&+�Evg��M��Z탆I(�#ci0Yp��́ߠ�X�^K�R�� ��êP�cDZ't�'x�@�U����Μd&m�E�Yu�m�+4G���}ji	�7�W\t�Лy����� ��tmZ�$���%i���
�8��][��v�ЃY��o�Zj5�� R�k,�4Y�y9)>_%1�9���R��Zj¬�F�.ߦf���*II�E��!y���X �� OZ:0�]��Z������5]{A"��s�_������#�*$kK���u�oojEC�ݚ���6'^U�8o�Es�S��L Zvd�j{1k&:S��y=����Rzvo�L�Ҍ4��b%Ux&)V <H˾�Z���9�[�W�(���O$j���tt�����1������(wNa�hD������Ր��J���<^^��%��]>�du��z8�N��k�S��1�
|��It���N���L��L&��4�'p8x2%|b��`����*����+mY�O�r$��	�wl�C65��O$!����	1T��A�x��@aVc��;`�6��Ȫ��Q���C��#$�Ҝ4ߥ�q��3ɏ����B��#�9a����x��e�c1�	Ñ����܋�{��A�v� n�T�A���7j �8�˞'>�R��8�aj�А�z1Knn:�[�ƥ1Z�mq�� ���-J�	GA�'�^�Vt��/�-n�N2w�u���x��5�RVl�Ѐ����~�xSX�e��hl=!����v�4���&wR@��X��r�HVJ�7M����΃,
n0���?rĘ��7G�MP��/6nk*�e��:�CP�2���qw�|�9^\<C�;� �Eݘ�"Qg�9 ��I=ɠ<��P-�uy��b�
}7˂��M�qQ:�d�y���_�� D~�W�ӏ&:����(l�D�!A�BѴ�XP�?bd���J!o�̘���O��Aҭ(�
��F|�M��5��ɉӶ� �}(�CkM'�G
�z�\��P��:Y�:��ʁ��p��!�����_����ʼ�<���C���c�5[�@������1�	��@����b���y
513��!�]�"�t��^
�~��UH��;�R���gh��*��o(k��ε��4�Da��n��V�6�[5��.;� �P[�c���>��?�j��QH��M��7:�Ȗ�Đ`r!�
�� ��u\o�^���q|#Q�C���-Ѿ�C�>#����5c*��$w��,���Iz#���`���َ�u#G&�����-��B�������hOȤ0Ù��,��G/6{�&��ȃ�)����X�6�A.=��oVQ������=�]G���u�$C��^�a���s�Mk�/5p�ɻ<���u��[���#H��^��u��9�r��A�XR��L��$Y�｜�S�O*Ԭ+f%1\���S>��)�&Q�<��c��r�M����tя���2�[Zx\˱I���p��
wȳ窴��E��h�=��r�A9���jcc�To���pp�6Q�+��O8lAK=��]�$�S�ɮ���ն��5[G�*0����r˝P��^;���3�6�Q5!��!8���;X�I������L����hV~���v� ];����Y1����3�ݪ�nK)�-�'�="�=��� ����6�|�%�rs�3�[���Nn��A-���6IxF� pt����4g�ԃ�Ey�&�E\%��Ǜ�I[��U�T苦CVll�:��W"�|Y6L��i3�}������o�e��:� `x됸��1��=�L��4��D�x����v� ����B��wΛ� ��w�̈O[!�dKc�YK�p������r0(����i��K�^@'�+�V�j�M�`�Ri�;�[f�)Dv�Z���-��NЇ#�K5n�RbL�8|Zӿ`�7N�[U ���d뤉�DQ&ŝ��FCZ���o`��H^ח]�+����ow�����j�͝�"�¯%?�����lL�q�MXuSl,>Xj��	�S���p�����k���V�{\�5J�Z�w�� J�Ha�j�.��T0>��v%p�Wƞ�ݒ⅀�<������Z���Hq�'�~�꣫{>~���>�	x��M��jN�"(�����*��w�4�H�P���oP�l�6��z��X�!�ԛJ8�e�a`gk��<g���.�D�~��S�5	����oF���ȿ�x�/]��1l�:��3���.��9����r���eZ}VJ��K�����}Ss����������I���8:)%{�'���h�8h�z��)���'}A��w�`�B�Uk8wB>ik�*^!c�U�q{��F��Kͧ����t��˲�on5l�K�����]�G�w�����L�)�+K)��$X{T���up�V販W7���Ey�9�L>��V~��ѧ3����/z��\�TZ���Z�), l�)�tK#���.�!xYz�h!��+<h�#TW(hA7�F� Å��| ����P���q,55��bq3���}EM=34�A�9�}=<�/�+J�| Բ�%�>�$-l-�����i���ʔ �nA�k!���?�)J��P�;�g蔇4�����	�v+2�홛�5�H�ќ��T��@�_<���co+ʈ���� 2g7.P�?ȝd�{Uh_��^c��Sz�!��g�D��,�<���42I)+|rsv�Z�M��3;L��m�o����r"���E.+���G��B��
hg���h�N�f�8����6��c�e�XKX��m�s"�&Y%K׹*II��
R��Wy�G��(��x�%&	�"�IL���[�r���`,����aK��E��p�y�i~��5���ԋq�J!��V��jں���+Bˎcbx�)��ǃ�{��͸��'4��pX��S��K�G�Z0 �9O�Iðu"i�<۴�O���&����[�51�W�����b���E<�4P��1��� ��ll��LPM'A�zǂ�O�d�~��MI�D,�͇c���J�u6��.�g$*aom�Q�>��+�`���E���,JA�Ӌ��*pc�́C׬��\�2�|NѪt{��S��e�0h!�v;S xb���T#���V��x*_%��eeR������M��ĩN�y�hx��l{z�K��H�q�*UN�=���Љڒ��|��h5���SN�rq;#�\��1�)�I����)���(~�� EF�d��y�9��l��c�P3��_<�VQ���C=���K����譶���&j��V�$��2�Vք���5�?��:��uE��.��o�#qQ\I;1�ޔ�!j(l���rm��o���پ2��Y��>�o�W�n�T�<����or����扨H�!Q1�J]�ȺR��$�1�� �Ia��!������5�iA�c�c���y�f�&���[󔧅c�01[��S�N���aۤ�-Y�b�>�VI;�������Y�R��Ÿ�]R�l��Y^F>��mV\y�U�k�ѳe.C]�q����Q����E�fFAD�&ŏ�#@������i%���^S��\�,D4��a��82�b+6HhIFe��� �+}�l&�q�̫��A��^r�ky4f��9�8__��*�ѝ�����Ɂ�V't����b}~ۉ�u���ߗ6ص	��[IeN}'��i�p`+��b��b	�l�4(��� ��U����T���^0�pv��e���L��>�8(I����Y�؇v(��T�K����ps�5�e�P�=3�!�����d�)��6y)��BM��LE�����W$b�� �R᳣b��!f�7n�����������n�F��>���.aD2K_!�P�cU��^��+�����\m �X������a�B�{����S���i�CPzT1���H�P�wf5�^��fÏ�IZte9g��U���FV^.7L���W���!y�	�]�{���U� Kh6������vP�}��1;�U��0hN|��qngX%���"	J�.�ҏ�7ei�'],���̎>�e�����=�=듧/�����h|	�>'�Yn�H^G|4�Wf�/v��J���6��j��e �L"�ԥ�7=�I��4��a��6�C��N�ȶTZc�3�W�Pp0�8�=�܃Ճ������WU,�a@E&[S��^��pz#!�w�s����O�[�{,ɛ�U���(UQٝ�n\��u�����!+n%#�����t��[>1j@�L剴+�Oc��@iE��7�Ł*��^qbȄL��*���0&��~hPv��:GLӐ&��h����P=�{���3܅Aޗ3G���_��0��٥��Oy��|�X��m���m?���RZqJ�1g©�7� �[��~@�u�È�8-�����y�0)މ���
�Y|�]��[F֯Wg�`Ms�������\�o$@� x���C��?��n�h��No6�XI��u�~;uD�E�2љ�AYv[iKte̿}z��dJ����^sI���椀<�.�����HM]�E��m�!�f"P@��@H�UU���]иb��'��7��(T�3PrYi۱�*Onz�Hd۸1��u*�:]�X1g��,/R�Du������N����Ɯ���~��R��7��(oa����h�5��Z� p���6�nt�Ւ5p7i�%�DiL� ����=���<5�r�0���g�]6��+'��Q,5��q��B�L_��N����b�ku�R���ͣ&p4̏{�
$�Lo�>A�S9;/��(��m2è�'��"$_��H�$��HR5�&s�A����9k�9���tP0夃N��f��_3��u;��a�$-\�����<`(�p��Qd�ap��.P�A���;���Ą�&�Ŀ��bCΗ��e�r�'χ�����?CV������%R��R^+	���[IoVhOJ-s�
�����1��7.p���. �xj�!�5�!i�j�}���0u�q핕�x ���K�g>D�[����X�	mkv�aO?oY ���n[�?�;�=8��l&� ��!�14�e��c����L��,Z����m�����Pkt��B)oS��Ue"�W�k\�Wme2���Z}�*����P�{V��k��>+��"D:��`�:v�إ���Z�c�J�8Fe�F
R�k�;
��H}*і|L��R!>/(`�aS�z�N��w�v3�҇�4��^?�s�$��u[��~����+NC·�gС�JΖ?}�)�'u�/�}6CCf�-W;�/����V�>[�UuO���a�K+L���h�U��o�^�5}��x� ��������=���%�ȷ|1��z�seR��+�=)��e��'b��5�������1 �Ǟ�!��&w^Xw}�5CZ�<��F��G�u���X���qX��q�FyVn�52��ܿ_��l�ĠFcC#��n6�����2�{r�l>�꼆�.U͏�I��� �xHT���K�*�!�������Aã�����"p���_	�{�{1�i������6�᥅C"�<�1г��"}ʝ+�aΦۀg�a��CY+�d|
�;�#T�9���W���*p��[dN�ӂt2��3K��mW^�vPa��9�,��|xg�w�n�E���c�X��c��ǁk�2S��uđ��(N�݉R�K�1gۄ��6�s�j�9��O��B-�-X磁K�� G�}&�ڢ��Y�g�{p�r����	r}��������}BW�/,��j���em#	K-a����X�i˺�T =��r���M�d�,�1�bR``�u�sk>H��7l�TR�An*�Ѫ���@hm�`���]�;1xB@���n^��my�	���ZX�Xg:�|A\Ő�	Ƣ����|��Le�o��rE�v��S:q��/
��lW�倝�cxz*J�y��<=)D�q�[,�p -����+�-�7A�g��Y�1;�t��x�S�{'L\w�WD����Ҥ��j���3y�ku|���A���t>��j�]�z�3�l��uŉ���SG��A�u��6}���r�Aû[ogZ�B
��I�2��v�cisnV���y��kAB�q� _I���"��zh� �Ϫc[�L�!Kc�X�^�f�G��m�@�j�cz�Z3zVK1�J����os�[�,O��2i;��s�mQ�]QV#��Lqf��Z���#tם��0as�%	d��a����G,����܈~�&������3ϧ���J�4����4:�o/8��!���_��>��t²�&�]]}��+N�OkR�3{��/c�Z �R�{�~�U7V���~��A:Dp���PsSƉ����}�mٸ���F0: ��2��kA�l�� }��l��ȪbO>�� �K���>�*�PƓY1F�b��É������J�rS9&���
_^�>]����;��ކ������~#S��qFSe��>�6oI9{t-pP6�։U�B�\������c-d���}K�)�^�[#6$��ʫ-x�F�����AM����u^f[�dGf�*�����Q�>��7�Q[��މ�ޥ�8�vW��\�-X��-'R|ke�b�N��_F�~d�ߕ^�MT�����2^3����m��3H��Be%~'��7�,Q��'�==V>��x�c]� �5��GB9��ch����Y(83�46t�8xx��埦-���`a*�g�"H.�Z�
{0�!v\�e�*X��m>�j������Y���B�����HP���(,�Eh�p�N/��#*�:�m���/r8�l
�z�m�0P�V�s�R�m�e[�_������Z�ܩ�o�)��vM���uٽvh��n4�*�{/�~5���i-�o��4���Rʰ�RŅ�J^�!��;^�H�G�*0w��a�zy����?�	�m��P^,���	��w� �O��ڒX��q�T)���t�H�nF����ά�n���A��eG��4�\�z�Y�k��A.Z�"
��䬂 �LC���Ý�N˟�eJ�)����a���`:*���1k<�{��n���wŮ�ZEn����|2Cj!�U_ k�vpzE5�(>D::Yg��g����"@f⏗50�N��<X'��	ڏD�&��"�\�ʎ�I��	l�\I�t�dW�q4���	/���ܖ��/�����n��ꕟ��