��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jåا{�\�u�?߷�dn@6�zf��r������;��1��B��dF��M1�ۿ����yE(P�|��MP}:�î����SМR�%���%,1�~��2"N0ڰ����f�Oz��,�
2���w�\�.J����.�(n}�-���~���N�]Ӱl�d�lh�L����{�f�*�c	�~�g�
(���r#9��ﮀ�!��e��e(�-5������B�C��gȸ�&.N�cB'%͠�ˋZ,Q�E��k�x6|���ƆM��85���Ȅ�������detx�L	���z�0}���=�$_91H6=}?i���7�f�4��&8_��0�oi�p�Q&bNx���-�;��5���ԆU ���3�G������"��&1x�(k��q�
3y7���C�_�r(<Ot�6*+�>��)�n)l�6��@�>�C�E;������z��j&�l|U�p�����w����	<
u-���^.rf����0��jE|+}.^��Y����Rhw��']��F��a�&�zu6A�+3�)�;%���'��֒i���i��C�9����'w�e�.1�&(':�נ��7�'t՘\
ǒ�U�2,�	��Q(g)�Ïrh-�M/d���s�������>�����n�u����UD�~&���R��0��	��sW��>�M{c�]}�i�7�'�-��䲆�U�F��PvZ�h���7o�VW���&�Ϸ1�X�g��	(�& �;:��<t8��x����L��1��6T8�>M=m�^��7@���:F4D{I��}FZ�Њ���e3����]��k��j�`[�\GS�V�����R#�mW��`�r��'�]8����m�	7�bY�˓Ms���z��.u���{?���xm��ݘ)-����P�R�#��l8�ECV��[kg��/�� �V����μ�v�g���eJ��̡���CH�=�n��2�M���3��v�h�X�Q�?ѫEl��ށ��*�@���_װ�O\{g�b*/�ޏ8���Ƹ$�;*��o��H.���j
��/�/�a�r|�3h䆂�G�1���ZtAR��Ѹ���"�?R�+��G�0� �^k�����ˁ�J�fljV�-�$������w������� �����I	�T���g���~m��(������L�o�x��	k
|�@�"]G��H��X�|�Ӥ	��6;�°D"pc����-��ar�רּ5�*ċ�j!�o߂C�E�կ�#v�MFKUH�40`[g��`�aنH�S��0_���)({[zԭګW�y�UF�oڦ[��[
v<�7���:�CEB�-Tk���3�km�2��~�kN�o^��ѵzg����q~xgh�z�"��l��)�>�[����zj��j���`)�$9���W�,��93�brH�d!�؊��ZS�u^ĬL��anJ�^���5�.[�Ǔ��@R'�6(͵"ʇ\'tn`��a������ԕqr�3��]o]�  ����Z6DG-���8I@ټ��1�}$nT:܊��|��mj�Ѕ8�P`4CnL�`&���E_|Φ2�RB�&�8�����Ww=��ငa�o�GUF)��O��Y�Qky=��qߜ7�04��狪��jo��S����K[��o8�����2Q3�����:���RW�8צ�HfS���{�`�ƣܚ�S��>�;��ݦc����дI'�l��q��O����7��JK<lX��tWP�*	P#��ފ�E�v��7nC>��]z��S�!�h��ݩԞ聤�J,��ZO3�5
��j�
L��"{��/�w�� ��~����B����:�(�d5��ոu� ن��oyi��&=��t+pQY���m�)��`N�^�#��)��6U�8�Hl*��_��qk"mڕB'�/~1��@|*����\9��+1T�����߀4�T��>����*w[Dd/���Vl��Qf�x��ߋ�����d�����P�n©Q(�w7�Ћ��xC�
*�V	�>%�(��a����Y��Sz�<38��:�+�{��p��m>Wh��n�{� ��5۹�5R8S��+(C1�*)F���#�B���Z8y�#�,�
|�C`�̋������;�q�u�p^1>�~u��\�=O0�MJ}�We�Z����џK���[��SY�����=ڕ��K���IP*^D��h�n���B0Q8�P���*S�k�I.�t���V:�`p̞��3� �a+�}$n��׈�3�z�҈���ց$�# p}'�Cq�7�S���4��f\_�H`�PHB�4�߮ew�skt#��`H��Ù�2�y�PU���]I��4-}8���~Ɏ:~��%lJ"��y��0;0�6g;!�4�C��G�mu+�Kq�Cg+�5�TfL��@�l������/q���+Y��5		��1��zCCˀI��Ĕ�T��M/��� �����fp��Y��i�&��ѵQj|=t1�m5����ʌ�Pm�s�\�Y[΁aȱ���X_��[�zB���&�7��s�Ҥ;�����{���.QO��`��z�_��s�S`�Ir�id���$)SK��3���}P�.�~e�+���_�y��ln�S���J��28wIFhˤ���$�ĂPܦ>ً�������E�8�vTk/}Ed�G�{p��-�ˠ>\vW�FY}�ET�0�p���bV����rgV����U��*8�xON������R���@|�⊹F��������>�f��?�fxD?A��h���&�U�����L-���,��z��%-vl�;u��5\��c[e��d�UvhX@�|:w�w�Q�����1�	���6�,� =T�e�C�]ϋ��	C�)X��V�����!�|�>�r�)�9�-�fWSC��\��>����S�!'N�qs��
�����w.����-�96u�Y�?E2�	nb�c9���K�Kb�@���IJ>���	��lu��| {u�r�RH����u�|���O�
��O��aA�Tо�Xu�X�͛��<�}�x/u����--�\kG����q:�)�J������g��
�L��D�;�Em���ֿ��Z%[3<_]ď|�K�%�~�7��0��!�Њ��GG��a�$=p]K���ncp�9��CoX'��U�S���Y���̛������o���8g3Ż| )��a`l���8]�JpM�:`��ج��u�6�k�>t+���Y~��Q���g�k��A>�5H4��i��������m���G�,Fl�\�R\̫�	�P��j
�$��J�����`V��M@ 0���C�A7�U�h�ǒ\�B�������W��meS�,����֩�y�:J�z����Z��8�ӈ�����d�5>R���(�آRy�?�ÈmVϐ�����g��� W�������� a�Eȳ���eJ��ƀ���u��Ɩ7�T+	�s\/�	� <-R��!ߺ�9A��[�R�a���t�f)�v�\���*Һ�7z`CW]�"+���O k"͊�Y�r�줳g�z}�az��3h�F�85�ItJ��k��7
\�{/R1��N�@3�C
�u����R03�* u-�N~�0C��݁�jB;E�l�n���v ���S_,鶭�1Sw�'T���)U�Y�:^,|�;m,��U��4`��^�e���@�e��k��rt�L�`ru���}�p��[44�j����k^�}���~濖�wn^� ��u�NsY|�)J�Ņ��#e�I�G5Γ.���*��Sk�#� ���F�f�2�ެُ6l��H$���|0���rjT�u_(�7���j���4�D�oB�u���}ǩO�=��ޒ��AQq1[=
oE��ܩ�ɚ���������m2>��B�W�A^�TT|4�D�V���RG1l���+�T5{9&�i�����u�]!zM��Y0��c�1�p� eW��ҥ�C�����pˏ�h
��ص��=��ƛ�z���hlҵ�eZIc2@=S_��eB���(Mx�P*��y���T�'KE�+�뢳n�p=�S���;��EW#����<w�a�Uxۇ�ФI������RC�ll)�'%{�������ADI�A��A�b�+�~Q�c3�ϩ
��D�8<|�`z%QG�S#����3҆��{�v�i.[K��5W5��=�U�*��]���"�j�V��X\�ű�=[�<":S@�[����COg*�#���8 �S?Bt+7K�)���N �p���$w_F�@n��j6i�p!OQ&]2#3�>�������"r�Z�J��8�M'׷��!���oɩ'��؄��J�K�S"���oұ���=�Q�MiH�5ru��$R�y�o^����7�W�"Cn�'��I)5��dٸ���w�t��H,c��C��w�n�QYƓiv�n�9��>�D�z�RT ����q�e�YZ�R������׹ۗt���*����tw���_�N����Ӭ����U� 	���EeS��N4_�R����E��(\G�L7���.\��{�|�R��Ra2�C�c���������E���J�g��T|���'�5\�`�4��x�*���P�XtfM��.�{7�H��b����0a�����^�XE�Sp.��!V?�y�7�Wc#������_�@fJ� u��U���y*W�\8�͔��Dè���Ewdd�/����E��aR�Ha�?���׽.�*Fa2��k��q�"ۑ�^��9��t8i}�|^
�a�̏O�fN�\���qd����G����^�T�$�Z
��^��J�PQ4��ԧ2r�WN�0�enc>^"i�)�k�ad������Oo'�)�J'@�Y�.ߞ�.АN�M[��3�� JGqA�4����*����{�h�y�03+\7��a��R9�R 7�Kd�i��j��� +§p�a������&ҝ�S2
�ާV���0c��v��~��Lv��F�{��r�T�:�F�6=$�ED�8�������?����1�����>U@�Grb�����Z� (���xo w��F��o<���h���Z�ܸ͸��'r�Ϭ�ّG��QN9�