��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e����d���f{��@����S��>���4{��ת�AO�Q{���$�O~��yL�̦�[�QF�����S@P�����L�x�D�&Ծ�SvD��lv���,���áC=8{�@&�+�-��/�F��])Z8	Ҡ���J�f�g�U�r����z�»_|p�ןYV�ן+z�D�z=���(�~���r�0k�����h�1B9�0��L���B "<�LV�IB�g�O"g��$�(9ZU�A����Ӏ&=!��<��Ѱ��u*��.�"�����6.J.��jN86L�*�8���m��0���h��p�Es��m�Ƃ�[d��^�r�e3�\��$��'�&��.HƆ�RX��^�6`F)�G����ZH.˻���/���#��c�F�� J� ���|_�V��(�4)��Љ\FE�u�����e9�M��>�/��M�Hh��&����w�9����z��(� �w�8�!�U��*=�lv+% �kF,�9�Q?iZ�ħ���I#�4��P���W�1?8˿�|۟;Y��7-�"�9�'�6��Z1���	��|���/l��a 5��t����`������;�#a
.x���R�EXF�Es�c�/=�)Yc��������(%k.�H"!ٲ%[��I��v��*� U���2Q�idtM@�U�0��"ZK��ER�m�(/�G~srOk-�m��(E��Q��S�Q4$�n�v�=T ����>��qn՝T��B؆��HD��`�*jQE��Qy���v3u۾#��n ՝93�HNY�x����@��m�	��p֐���Џ��Z��e��.�<Ъ��]C+#��4�� ��TB�mζ[��+�,��?I��4�i�}��EO���ی�L)ѥ��� �EQ[��v):z�f�&��s����l���~ug���1g������{�t/����=#��(�ۛ��H4�he�h5D)��I���/$V!������'�#������s�Ya��pU�D �����eBڬu�A��|��4������*�aȷ��cD{�L5"�fu�� ���DP�IW$m=a��N_)HA��)� Fr����x�O!���yi��Ak��/��,˖!�56��ꨔ�Ԍ�E	��#��'��[��:�x���4JB���=렁�����L����i��J �$������� J�N[�����YO[�z)U���&{m dXe���<�$�̫r�&d�Wh�O(w�2C�'��_�L
mV����m����d5���S�/ˎ"���?]wX����O�׼�S羜 �����d�ն�1�'<Y��yT/-:�D�4�AXE���D����`��^�O�ƍZ:n`����(�:^s#����L�D�o��Rc�:��y�=�P^J��4� ��g�6E���	�9ݥtӼ��R����v�xf$�7gM���b�����џ�6����ڛ��([<�މ~��İ��"ɻ�4��VOkw^���H<���G�c[0M�'�b�6ΆY`k�Z��|D�����#�ve��܂��H�L����`���V�c>�}�2�Rv��0�,1'�k<]����0�@?�s�M�Kl UR��?,���x�xN�6��p�sr��d߶rqir�ɩ,��r5{���XB�"m�4��N��PA�����,��8��0mZ�q����=�Y�ȕ�zG�m��A��٧��|�>�N��K���y�̈��]��Ҥ�6%BE�3��c�X��N�����q���`iʢ���s-7:�U�OQ)�m���>#� 角b�̇��K��?�}��R����W�Qk�1!3�A������9>�;�mj_�ZC�����D��R9�p��S�r�:~� �d���4�H���ML����]���μ=E�g���E"=�����E����ՠ��@��������B�Z��F��#�#��R3^�h>����Kë�>�W�3vVA��M�������:�C)x�'9��3�[�4X���0+I��N�N��(5��X��ͪ ��'t�\��'�#{:(��Ş��}e#$p�-�oKUތYxn��ƽ�� asr9�Om��l'��5X"�?x�`}F�?�/-,��,K�,�MTO�������kRf� �������)�'q�����M܌)��� ���E��"�{��[����QY�ұ���
i�*>H��aD�id-��"=�	Y�T��,�pmh3I)�Z�GW��(���EW��6*��x*r�u<_O,H��T�ޟٗ{�%� ����fM��S�0�١@�Gx�%W�F�����d�y��rv��a�Y��rk n5�k�H@ε.���mcßl�B}欀����7�������(�J��ޛ�]����2LjYq�����K"����+�2)�ZSH� a�dӧS�X��&��9�y?%G{��7�U�����Q&?Q
��,�®��$�%(aS��pP*n��ɚ�G Tԩ��	(��@�%��\��;��4�Wu�zP�G���䖋�"�?Si�t��f��:4��08-���A;���>�v� ��W�����R�n!�U9ź��V�|���U�2���-o��C{�uCJ��(�=�I���A���j�q�~��S�yHx;�@��
��ӛ�猻���b�/Y3ļ��#g/�����HU�%WXg��ut�7ά�Z*�F�' �� j ��ξ}u��B^�;�����z_傿윀I����34F"*���ת˱L�W�f
^6bՇ3��7,�K��
�u���٫�̆��]�k.�umɅ�ln[qܸ��A�������F�$C&�y+�b�TuA4S�Y�9��`�,}ߐ��|X[D~d����T��He�=�q�#A %��H����lD��'9�m�D�=�5��&��V6U��>�� ����M�¡�5�!���_����"�o�Jx�Ij��C�������dr���D��o���c�C������Uv0�iwr�*d&PH�LT6|��c0���u ��Ԧ�5�κg��W�p���{���w���,;7��1�J��ň�x�^���H��r�o���4�I0�E(�d�����B����z��u�i"��Wl�$��Z�G]9͆�����v�*�4�������e�Lr��>���d��L#�&����v
e#1&���B�7N��n��k�GO{���<N�uq� �m�Z�7V�U?�%!m|����h+��'�eM<����"��h�|�p	�n�7�;0�,h��'�Y�N�/cQ0�=�FSp���T3��)#@�A�a޺�گ��za�)��Wm���`��r�	K���&��si)�'����F�FY��sύM=);��s� |���2�l�����R�: 6�a;>�;ř1�g�yT��*�X���J��K��qT���.y�_h���U�e̽(�� %Y�JD���po�!��Yy
>O�.��F*�~���/	$���P|���;�@� n�}Kݷ�+rA[��y�ZLU�>z����]J�W5��-�� t�*�o7�^��*l��-�
l���b����v�I�J���Z�G;{݌�q��g�~����ẚ5z�l �'��J>s�@pcWN%,��%	��_!����"��m�z���=��M�a�EbwAY�uD:g?�I#_�
������5�ei������ ݗ�M?��{�6������G%���y�y>d�"�j9�vK��N�Hߠ�]}��c(�b�`t���Vvw��.�d�ʛ���р)S����/������2"�K�� �o��p�4L
p֦��6i�&U)��}���A��45��ސ��RXk�3�1�wv㳦�
�<�������"�%{���mB��X�b�	���n=
_/�$X�r���ȍ�2B1�<�I>%g��{����y���縊�62�uSok/M��{��5�	��$m��>�qV K��APo&ɞ7���O��O �2\��̙�e��hYw@�7}^�H�"eX�zk��3Wa=k<�����1e��Uू.��:�1\�?��}���G ��G���3ā��ԅ|�x[E����O�k��2��QV(���ka�E�R�ZH�q��?��r	(Y���W!*��0��R}}S4�K��B�^�Z�z_:�ʯ���������
�%=��Î���a㒡������ �RN9Yꏔר�K��9�1r�&^��*u��@i�����edO�R.�)�?�IANʸ2,��uW�B{SK.�ِ��\��~�����(�E$�w�ՋP�lH�L�����7c��\�������s�ai-L�b0)57ߔ���e.��=���1+�3َ���Q��Js�u:�qސs�A�J���ù���L1�\�奝Ip쉑��,`�_��T�4��e��v�cG�k�b8�3���:�cMh�m$� ��pb�2���Ŏu���~�|Щ�S�Q�4{����\�42�,c�&P�9�p�I��E~�^<��XZ�@��::�A}�,�c��G���s[������Qj���A�lKO��k�w�n����^� ���`���LVY��}�Ĕ�S�1�lߴmq���ah 9Ճ^��4T��x/~�˞,S��Wqy��*he�Kl�i/oDM�h]�:��-�>��U�.�m$����Q$?�ж�Z*��_��m;�/E����&\Ӝ,x�ih˸�6��������F;����)7p�c-�T�H��.�2����I�M��ZrG��v��z��o����݂m߆u��u�E�:�[mφ�F
��hsF�^?��o)ߧ���M�9"��o�
i��3&i���'����wC`Hf�7��j����d^��DU�����H6���9i��H�s���<< �;���%��n��X����$�2c��Z�%p8-(�^y	��o�yem_=Z��mO�=����:�\�`~�)�X��Xd��C����(3������*���ܠH�?�e��~��z�M1H���@��'HJG�P8�Yc��"V�h��ϟA�4��R&:ojQWZ�G"��3�������|�i扉N&���� �6�ܷ���i�L]�˱F���DP��T�1ih�����-ѐC�ryj��`����Y��v��<�[8��o�G7�(G��!.u!�^����`�I5��62�s9CǮp�����)c�­��=��>���6�#OB�v��G���$&��%�5�U1�s�_%Lp�[��B_�`h]7���ِnG�00��o�}\��y!5���� tO�r�}����3u!=%�.�oᆩƻ�rqn\���ݸ[��bi�A{���O���5��5��M�=��S��F�K��(1D1�緍ϔ�D��4�M|�ѽX[�ᷘ�
��u�[����3�3m����2Cj������H���Y�������;����.L&
�>�F`�5�E����<���d�K��rT賟�Q��}1C-O��qZy@���K�V�����C�[�	�Z����)!~h��+g�m�������툢U���k�	8����;:[�<*�pvG�k',�a隌4J�>9�^e��yC�=@/0�����S%�4��+��� W�2V\t%#(��w�����GJ�sa�p��:?�a��^}��$���>���ͨx�)�C6��#��F)U{��=�Ledb9@å�$"
��l��&`x/�W�G�B(KPo  ��`���a|�����|��mBjc%��څ�>�f<��w]��;�^����7
�3�H�0ꃘ��"�g@pb��My�|\ś�<s��1������G�vbr���U۶B��RX�&f���\��f{�#S���N��S��Y~LVJᲛ"e/;R��&�M_�:�Z�fd$;��U���`�%w���Vx6- G�.��7gc��������F�4�0��0I���2ms�x̘����Ku�cCE,��� ]'��>Ya�i=�H/d����׎����7ь��d��O��-��Ŭ��˭�Hr�o'�V�4���S- ��$�[�9-�5�ހ W�Z�Bt��6�Ym4��Y�����}�MŖ�Y���h���-L��-Z}�Q�^v� ���8�R"%48���yp�4�v���&��@�x�5�K9����@I��K<g �����Ժ����*�u/2 jh$�z�C�zR��g2Ud��Z�CWˣ�Mu�b\����&�oo�P�~�7���)MMx��m��$ϴ_y�t+���u��M�Wj��M'���Y�BeGPp��|��|eX.P���0z"�B��u/�3�c���>�K�Zh�/�3Ķ�uJ�J���݌��F��5Ӛ*Pw�@��B�h�J�*j�Y�Ȯ������-��E	Ҟ�˴���N� 9zL��Ǻ��8K}���A��$��a4T�"�}���o![��d.Ȃ?�K���F�f�Յ���0��er:ᰍIx �ҡ�j��(Oễ9KS�'�/���2C��w���F���\�q�տB������Ąc.$ɝ�*���Ѿ���>���*��=�J�J8�?�p����K��Q���E�.�fT���U��4L��� g��KEL۵a0��-.���w#���#�G�����vY��V�l� (�3ϋU%���XUb�H�Ҥ��@>��ކ���&͠�UC�<��k���踀�X���M�/�k|��=�8���֔���������z]��{hkM�V�{�#��V�[:�M[[�]޵��Ф��p;�tw�1�U�cT�s�c[�u��rj�!V�GŊ���Ju�!�Y��36nN��~��\�+*�e<2zu��:Cx�
��:���N��L�Y�]>�m��:�f�/�n��3�V��9Y�A�֪�FfK-a�O�m����j��+ 4��U�{�7Y�!��1����|��!&���+^�hN���l-��dfGo�2l۠2���� ^K<�P<�Ϛ�3��M|�mh0=k8Q���+��y���TQv��K�ԙF��è���B��+B{g8���*���43�Oc#U?�Z6Ϛ�\�q�2�ک~�5�ܙV�r���aa�"��)/���t�<խ7����>:j{ɳ�A̩F�߄�5b�����Aj���Q,W\]@y3˜;��,�������B��ߋ6n7�-΅n��yF�Ido�2_���2�Sn�J�Q�)մ^O��*[7������w�ެkv����h*�d滐H��I2���g�>Q�߻�!�S؜�r �ݞ*�Gv,fx�	�-�$���ՙ��
hrU}`�C5�v,1�F�p ;��oϕ�(en˙�p���K�T��/e�N���E��N�?��ez�>SND�;����������6UM���/�/\tuf`pg�T��Q4����MK��[U&w��޽��-/�)���l������W���>�{�u�~���u�9��G�`^	��՞#d<HG����H	�����	e��3��$�d)� �P�����RɼR֞׼߉��#�8���kU)��R�DR�b��G��;a$
�e6��{l!B��ȕ+wa�h wpx/Xg��3%������a�n=��M��<�yq���eh�gs'e�X��H�M�l��Wk�x�P]�C�6Wl����Zم��(�4��zV��Kp��S�1?�o+At��ʁ$��[��<�(�Id�!���n��B%m�k�3*K�4r#�f)�Y0��0|<���r`�d\�<�����FJ�]�N��`��B�C��{��I�ZWT|Z���?�8z��H��G�.���-��.]
P>�OM����8�.xQ���>1n��oo&sN��5���%MFj{�}@tz�ȹ�P�a�D����9 ��еu+ ��@1Tόp�MH)ߕ���s�9Y2�뉇	7�N/���S˳͚Ui�e��a��Qm�!#�oxa��I?�~#�_3���(ZnD��*�z��:M&X!����À�'�GGL���FD����K�#GMz��szz�Z�Y���+�P��Ɂ����R]1�E%�h�f���ؤ%�����{�������a!6x>[�A2!T9<	�#�ɗ���]�(�:R#K�����$���y�9�*��j�;��^�R��o���(�[�y��/w�@}kl�i���7ɕR6�3x�G���
�6�� 0� WM��o,RR���k�J��*"�ȩ�gx�,tuEla����|��s��E7��k'�H�Bo�#O�S���&�h]�A��'Gf�j���p�z��ƫ ��B�wV����g V(w~Y�^�y'@�Wѐ�.γ��;�Q��l@���"��?��Dn���&М�r|M	��w;q4�W��f�: ��+�`kM�)�7`�b]�]������.b�wNB	���~��#	H"�cAV��^�0y�
�Y���g��O�{�5|����	�0�|;h�@�k�
���m-�_Zȳ���6���Sř��!^��*y�~r�!�)(=C�����~ Ju��mj�ߐ%��=���=�7���r.��Ozo�F�^4>�ʋG�\���Mx��|⍱�P߉ށ�0�2�h<�D�nw�b��%>2h^���A�
��x3�'t`(���Gh3�UhT���i���X�}Ͽ��6~Bg]���(�i��K:_�naZ����uÉN�����6��d�2N��!��\'j��2ǩ0m�m����xj�x}	���o{�Hβ�+U'��+��iJ�)49� <�^�#$�m�%�־�_.O��ߠX����5֢�I�UV{y ʧ)	�@�Ws$�,w�a?����7��	4�l�]4��;pi���d$yђbm0�؄�z����#��� �2-Z(��V��'"ٔC�����0.9p�������]�$���zЮ	����@�.��@�S
7�g<O�WW���r����v箠Ճ��#z��g��]�J07ۚ�"?v�J�/^l��.��IlˮM�Ĕ��2��(��c%Kjy(h"P%�J���	�jmh��ئ+EF
Q���r�3�gf�L�kyY�c�&�
�y��Hv���^�8e����_����B=���$#���L�W*����k5���UO<�\���鎵�jx�bwuw�o(n�Av���ֻs2,�E�`d-oҔ�<�Qa�9i	꿺��N9l��0�c{s����S�S�J�TcO:gN��l*Ҳʶ�HB����]T�2٬.�>grlf���P�)r��!����hm��|����5}c��U��\�E�$�Ge��o�`��,�*"�aJ~~�:Ge�(���KJ�1gI��_�䂴�E���۬�q1]����a��R�M	0aq|8����Vha4����I<���Yh�C��)���Ίhr<o!�$܄�,XGh���%u�qS�ʰR��砆9�� ڕ��um�m+��q�7�t� �Ȁ83}�ĺ��U�!�B�JZML�H��V�[�`����N�	���j��.��W�����!��B_?9��s!]h�P$WKY��f��i��3-L͏`Hԏ^ַ���8 92)!��<~]3��#3�ս�H]!f�]��Klf���Z/��^!����~�v�}�"{�Y�#�U�J�'J3(G��"�%��9}>�K#|80�Ep@��Y��7��V�ܖF����EyР�	��X6��|�n湬@��\�a�a�yQٳV$���/V_��m��V+t �/D}JDr�,BA����H%�R7td51�{$�s���%x��}�^u�]_
���K�1�/�/�.]�+��Wq#�i�2������"B�ń��b��J���%<���*���f�����nf����(�E�IV�]�^<q��x|��XZl��#P!0 �A<��tF��i3��'�e��̘%9r )z��Gm^��6	�N.�&��Y��1�o��0	R�n�	�Z!��<K���w���%�5�j�̢)I���(α��/��e�r���7�WE.�	�~�s��:
PDK3;�Q@8�r��"k����ֹ�� q��5=�=H������(v�U-3ʱ��7|��tFs^fx�	,����_.��
����Q��I9��}:1mO$QĎvcP���~.�1H<i��!�$;NV������+u^��\^#� 
ϖ�X^R��q�Lf���"|@���o-=�i5nZ
8��/�km��Yx[��� ����+�^WJ�xl��tх*Lbӿ��$�Nc�Sw�Ap�~�k��bfa^���T���������.���LyA��DOH���LT�>�����ͱ�D��N�`�J7C���_��.��� ��)S���NC��o)5E��[��Iy���
'�'j�$&�x�a�l�qu�&�{D�~W{e�g:B��^��^R�����~�)1
0��!/�і��󼹒�⡰�����ᕕ*���XQ.�7/A���N������O���	�ۗe����Ǥ�����v/@6�p�'��0�r-�q����_��Z1��`���C���������ͮ:A��,X�E�k������eN1�P�^��0r�}��l��c�n�rO$a��r�u�_0u.�:���߄��D[VV �G���V��_��-��V�oe,�z��	��C�ݪ��ea�k���8��@�İ" 9�?b`�P)N����4u��r4(�Y��vعp	��i0{����@�¿a�O���OHK:�<dfQ�2D�����b����r���v���n|qt������r.#=�`�����*u���8�)��M�� \h�r�C��HC2� ��>#���k�S'JL�%���������$!���ô̚3,t����a��+�f	�����6C4;0�yi[ԑ�^}H)��/rZ �>H�[���(�n�֌��F�k�ɡ�ݎѨ}�|V�6��v��5�YR�-�sӿ�D��=S���d'FUt��,uNܮ�gt	��T��l��g��V3�U�2Ë�8*-���HEq,�=��X�0М�-a�s�ݼ��QP`��2(�ޚ�U:��k6(�gC��~Rr��1n�P˵��l%���b;m&������+À�+���� ���5R�/�
7�M`9�L n~���駩�\ ժwј:U�F-ip�I�4�]Yn���Ow|��֎)p()U�{�9�R�G�V�w0�!Ȭ��:^}H�M-H�l�vA49��O���A%ӛ-�J����َQ��	dv�W_��Es�*���S�B��R� u�����P0�j'�s�Z)�������g�j�)k�u�e��Ů�z�^My�A��;��2~R;1�I/�����2%�I���3,�e��Z)JV�0����r����I���$>w�����֋�*��~wd5j���lKS��Z!��3�F���=z��L�uM�󾷝��ˏ?(
�fz/����N�7c�u�Li�y��F5�����D٦߉L���g;�a�M��V�b#m��S؅���`O�Φ������l�� ����j0��+��_�A����t}�C)тGwoYL5��`�9Θt�(' �A��B���Kͬ%�`����k�i�y�5��t�̑$�,���e�i�B�8�Oܳ�yנI����+�sS�j��`e�R}K�Um��~�b�v��.U+��};D�z[]=��%�L�􃍙�՛¿��)� ����S��,����9#Ј���3�ga���G������w\*���?��#�8Iiv�OE('K�W$؎���d���g�0�5�BG��Vq]�2w왁d<�̼�o�'P=��Z�.P�!���f�R�JA��e�A�'�ظ���Y��
:c7A�O������KrC��F�)s�)�rȾ�h�\�+�t��Н0?�<b]UqQ�" ��S��ps�&��<�2�\n�`�lci�I��K3$�w>�@05%�m�-�2%Lۂp�#�ė�~SS�^��3�^'ze�e.��&d^p�"5����� ��}�"����|��2ݸFmiq!I���͍���?>��z�`:hW���𫨖��P�K���j>:�߷>�z��S�dؼ�Z>�NL��y-�Ԧ��!�US��i���tp�b>���q0������BWtHN�� �~�r�I�=Dt!�l��V"�@��ץ�8������>�HC���0��'�c���b��A�3'�N���1خ� �F�YU���9�/��:f��&�@v_�Q�x4�f�v��6��HM+�*���ourn(dP۪����*Y���v���`͡y�I^H�8#6��{ة�*[�<��^|h���T ��.�5$��F	<�,����7 *x�ب�30�Sl-�xJNv���?��
X�O	(8����7z6�OAב�j�����"���U��n#H�Q��*aoo�J#v�	�}�=_�np��3 S��|)(pGE�%���X���?��6jq�wJ���wm��>��'� Ű����=s|��ҳ��m9��͡~�:c6�b��/.غTM�;'��GV}O�ޏs�oV�]�|��==�ߣj9Ĩ����0��KʕE��B��N��&o]c~(ti�V�^�y��މ �H���s��k=<���	������{7zg�^���9�!���uPO�CΑ�?3����qFbFezãR�+���;�w�Ŗ7B��k>G���MD"�V���lBl�s�?����+2���0���r�;y[���B��nnחݹ���"w�Ӕ?