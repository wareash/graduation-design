��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|݅o�@
�nI�֛TU�PP.�����+���u�Jf]�ϫ(#��$�r�jO!�Q%y����m����T}�R4�?/䃭0����AU�(�ƾe��������f�7�m��v����of� 6�{�
|)t�]з;�Y7�^(Q�`QԤѥ$Us�fӓu�CQ��rƙ��t��uī3�m���j_Kn���&Yp"8��_�X���qS�������~x
o�{��0v1�N�^��uv�N�S���@:gW�����ם?��S Q� �8^�������?L3��j�+��ڎ����Y#�3��X��\.�#Y.DӪ��8�WkOo���?dJ+E|!�3z�E��t��z�s�ۛR��#O?�{DJ�l EJߐ-'���3����F{L��d�� �;[Hn��jy�"�E���si�嵙u�}M����G�㩠_o�߁�2�Ŝ�<v��e��A��K�'Xs�D�5+�����K��2���ͫL>_��N�D��Rzʛ���G@H_�Y�����"8.�R��-�L���]��)x\�`�(sp�L���(�G�;��
���DW��g/��+�=�͛�h����l��&�n�ܨ���ɠL���m�8<g�@A2v4����8�z$�}���@Y��n5a#�8���	����9k|>�~���TW�6k�4�����[�C8@jSy[R��|Vg�/��>�t5X�ūe5g�ֵ����U��Hķ+ð�Px� ~�3�.�/��I��-x����_����`�(���f�Ԋ�'���C�o���3�r#Q����8�������Q��sp+U�^ə�;5bNG���e�5����Y�9w�d���6����������8�S����R���fa���=��sP��i�?�?Oq��ոo�M��;�����u,!8+���Y<�*��m5��[���K��pҞ��g���C�q#��S�A5��eq���0X���MO�>��s[.���!� �BA݁�ғ^��*�	i�!u��5A�p3��ΗPX���A� �������8�yu�1�F����D��b���G.;�-�J`�M��l�1�>z�R �0����(���<�9�08���b�u
�Ց�φ��zpx��}���"2�1H�k_�:G�ͩ�>���4m�:���-U��8�%֐��$'	H����/�Z��C$�0�V���A��0^���k��OUﳅ���oD���Q�,�S�������{/Bu`��MR�'J��D��g`P��U�N��s
qy��<�OSOf�f��#̂�`M����UOC-��o`ZC+zS-����Q���ا�pCO��H�Ά>/?���'n�����~��~_���P~U
C�?V�I�t��a/I��b��A�!�؅�HpG�]@�@��d,N���*�<���L�̻y&���i��֮���ڒ�vbtvI[�XM�ǟ��}۹i���Z#�,2�q�}q���u5~�;�n��Y�u1,H��^M��z�*��5���$���;9���M
��4QO�/�V٦�g�����_ .h�q�������8��{9��n����?�'�p�*�܋�Y���97"#�b���<�r�H������z:�yek?��50��D��X��J �c��&/x��3���,l�~��1 J��n�4�L/��\�Ge��8�i��8u�Ź��ײ�}�v�u�`�{6QZ�a �����N��Ѹ͊��U��(�H��=�b>���-y0Oƌ��'�xZf2yfzx����R<ݶ<<(�����e�X5ҫ/�$A� H�����˲�N,���qك��\�H�Q�8��ߩ�?���Pu�w"�ɘ�XIU�'�u��l���	ּCĩ���>���o@�"����F:^cyV�8�\�U�YM��>OB��q�Y���SQ"G�c��)�PvΥ�C����:������y!ʁ�ʳ4Z#�3~to֪�6V�x%�s���숑6�ol���syK�k�!T.��Ý�*�.��t�)��~
^���2a�n��*O Y��&�B�[�[ٙ�z�_Ј:��~�ߜu�,��Y���&R|���7�Bg�����}���M��g�K=_A�HX�uQR6ۏ�x}�����x��!hj/��h=��H�^�'��=S\�t�KIK��*)����D��]��D��t��g;?ƭ.�ve�dD�Ou�k���U�J���Y*˨#�>�F���<
}0z�2��L��Rn�o3�&<m�?���e�vM�Z=򞐁�<��P��l��y������]
&2�M���oۮI�-���uaw$�	0��d�?<��mu���u�<G|��O�M��Y�[��`ͻ�c�g�O_�(ZS]T��v��cO�Wf���pZ�}�M�6\���}��ƚ��tN�[�A�.�rً3K����/��p
1a��_��YU�xP"|dW8:p�h���|^T~�Y@�WF+B�/������0ҽ!�\��h�����gߎ��o�����^3s����fҗ7p����� �F���8��F�^#�� ���A��x��Жl��vj����1� 2j*�35�](�L��W��b�-�ۖ���t�$kaMh&v���������옙���'V%9I�c�!@�ޤ1��W%O�D�e�ݳ�GJ��/=c,�w��F�KL=<�D���.j����̧�W�!�.9���9�����3� <(��Y�#�F6�{1%�cZ���m���ׯ�h���=�]�A<�D"[J迄ܯ����}кtP�=Y�1���&U�����Si��� �O�� +�%�w$�;�
�T4��so�,��)QYBLU��YD�����O��Q��Ƕ��MJ�s_.S�Jo�qj�\VP�'4�O�֢{5`��<�]<�m��dy�9���}) �rݩ� Qj���l�$g� ������un=s�u��4�*�~	CC%��쀱�����x1|���7�\y������IBoz]+p�$�n��xJ���D]�S8��H�V)�)˙�6��*:�]��D��'���t�I���[}������]sh]w���YRm3�2m�7ߚo�|���V2U͊Qw �;,c/�N�y���Ǎ��/���V�����O�Æ	5S��$e�>�f.���eK �!'�aU��gZ���������IpvS�P��%�bI�b�7���t=r`):ȅ�Q��� N�<lT@�ݍȡȥ�㋒N��9����2����M���/��n�R��#�9�׿B_�fV�q�5K�x0�8�Q�rw���e+T�Mp�F��Y4#�O���L�/�ް��z��`Q�� k_��>W��b�L5�I����hߞ�4�b������ �_L��{N��0����9�^?q%*_���z��{�w�ޚvgB|� ���]��^��/�b,�8l��!@�������P�̢�1�'��P�>:��R���>&�s�����:g�Ѯ>9t/��t�6!Owģ�B� �ʵ�w���hk��{����J�n��i�{pz~+�*[�`���dH����b��@��l�/ƣ���z�T��䀧?l	�P�/�]0*��&uP��#�ڛ��h
4��w��B�1E/��G�#I:R1�owlz��p(;���:�F�j�ƃ���B�J02W��_E���+ӣ�tW�f�5.oFA;�/c*�.��&C!�ϧ�z��N�b��>��'�gC�h샑�6E�����)g�sӂ�a�@�sJ�L��K�)6�z�^�sL����@�.gs˸n=�� %	|��5�@��]*� �o��ʍ��?�B�y��d�B�u9u/��?��z���<o���UjRK�Ĉ�gHR2U����
�{��m]��/V}^���rU�䶋���\cқp�M�gNFݒ��?�AۏTt��7$�dϪ���f
�t���>�rj�A��h�!L��|��"�����+V)v�����Vb�~��\�=�F*�%��b�C����E]�rpЪ�@ ��T7���v��[EU�6��d����E����ae�X5���k�ߑ��a��,�3�j���?M{د�d�:��nbπI��H��x#$Y Ks2���P��Gʷ�p����>��Ҕ_���ǽ?��+� �]=��#">��P��%G׉�����C���g����G���̷j�<|`�p/�4��e�"��_�9�x����h��-��V4*�5��®�r@�yHȠh���4��9D��sy�OR1�L�;�gJK'=e4:5�Q{\.��=U,�e�C
E�%�.���̼z�W� ��\�x>y���2蟖�)UgV<�O;�Iz���1��i��BK�qjQ���� �siۛ�j����1A:��m|���i��̚؞�E�|x(oU�Q��GKJ>ԫ=j�4H۵�q6�&�������z�	v�l��Aj5�.}X2E3M�|$@�ӑ�O��'~�H��L�o�؞V�m��������P�\KO+�1^p�+�N�*�p��x(�"��%A<��T����Xqա!��zL�7��C�ߑ��H���I��1`�Uo�D�����k^{���/&Ƈ� �]Hnk~����ٯ=��={�z̔�&	�W�Y��j���uߙ����6e�<o� ��;��Q��ǘ���Sk�C��_D��X\*�'��e����է>�PD�%o:/it����8U���o�_��S�`d݈$���R�R�G�};�R�[('XP�;�$]�o�1>F�{s)��9ؠ�3��'u��%;�9`�G,�_�9&�,8o�Y�l�>��G7�&��8��?ب����+���a�>a�����=�3l#7z.]P��Ľ����ɵ����G�Ό.�Bz*�ޥ����^�������H���p�ch�����R�(�t�U]�d��f���_bo��Ѽ|��>�N�y�#,�o�n��\1)�����q��k��vv��w�N �}V�~�G(���74)�_u�}s������,S�{�'��zD�����J��d'���ٰ������� �?}���%�����q!CM��`��N�dsx�y}j���8�]��Q���,I�e��o��&�$���ѻ�z�`U�2����!�T���}zx�YZ2��+��:��˶"�<�f'μ�����GM�x���f��7퇊�MZ��}���v��@6AZ��zN�9cl6��8#:�zE,9�@;�����l��>�}���M�q����f���{�m��6�Џ���ߌh���W�4r�Cl�1���z�<�~��h�ӌ��h��6�@�\��j�z����U�>꫘B�:{h=r��&�Nnj�cv�����myH�Ç�2d��3��6ۗ{_�0=�j����[p��k[�_$�q�u-j�>3s�J8�!�1�({%l�T�wU�/��-��(6��t��8�V�0W	��)����1���wJ���nW1<���;���{DnR�h�w8X��lْX�����K�
"mdi0���So�iJ�ˌ���
�A*'ϧ� ��y(���U	xqQt�~�u�}"��ǒ����h)�Y��� ��t�4l��5�1�n߃�٦y��9qMi[Yt��)F��iP�h��"3�ٔ�U���9���+�ʊM�0s�$2q�ء�5]~�DA�ZAd��Y岛F�24���l�J+)����I�C�g�m�9a��`hh��A�^Ď;��[����:HK!�x���iT����w��.Wh���9%!��H\����P��n����^C�b3��L���:��y:��]r�4�:-@���޳�3�c8W��X_��x&\#�k�x��MO5�@�4����4*����ҫ����{"�eud�\��0y�(����4籫���Tŋ-w�SvK2q)v��ך�d��?bĹ�9OP*�SY5�x����V� �8L,Z��\���`L��E�DJ`
�i�Ҥf����`��ђE<U�)�,2��fD�cT��<��"Ý����� ���j*�`Ql��7(��<3Hx�Hݛ��K�,L
�L������CZ�&�7�d�a��n�G-=7}
*�F(.q|1_(Vl�O�"}c��RYÇ��Nhz�J� �d0�i����T�
]`IF*���Ƃ�ؤ�#�&�'m�2�4E-������tW��<��,�e*,S>eSv+�E��c����7r��ET[�f�k��H��n��K�;+��6؃�-�y�����@�m�t�TN��=���Κz=y�B�*�vڳ�܂�j��̈��p H�3����L���K����$d7
�kl6gE'\�!ڌ2��.��C=��]��H�챔IZ  BH�I`�s��'w�k�N��|��5����n΀2?iMP�_Dշ��DQe*�JU�t4��fŖ/�j�N�y�-t���V�)k);}ny�����=\
��vZWU����e)g���g��8�����UK�O���3h�(���Sڿ�a����(��u���Mѹ���l��k�uk�6��I:E�E��6���;�%��zqkC���8�e�3?8�+���@X�; �w�Ӡo�ƾ���Y��z]W�7w���!����ŒS��0��ܲ��M��-����*��.uP���d�y��[��>!0F�k��s4�+���Q |��}ꚗO�l�u9.w�F��2�%��H��@^!�\X��Kɕ]�b�Zo#�?L^՛w)=������'�E�.��vib�8�y��%"݈A�d�pVP�cr ������R>*7	_���cڟ��}u�-�E�j6�r'�N��N�yTY�R�x�4�C��G�Mt�ޕ�*�����sݲ��	u�C��O]�Ğ7�2���7�H��{��W�?��������&�����&�A�
ŐcŅJ᭰Ix�e� ��"z�QCm�=|�Ϫe[=m���nfrH�{k'?�Hkͪ�^��u�G"���ct9���7�#��aǘ�L��y��F]#�M:�i�IQ��}ĸJ�Ld#{�V�[_1�x���l/!�$hbv�T��V�c����֝�x��1��_�7+��g1BW�Ss�/������w�Ȟ:8�-֯:�U߅���v����	r�d�i�_bKwR�\�@_[�H��I�[L�����4@�3�I��3�D��)b֊��#���#��G�3���
j�� $C���(�\�T%Ε�s�����������li)Wt[�B�Es�n�e���Rv�����n��ݿ0⊻�#0"��N�Ẽ��,H�����S�֐���ʋ��d�s��{�X��dV0MR+��ߔ�w��X���b���nʼnn����eXs��q~0y�8P�F���HI�t�Y�W/\-�C����X�B��;�LsDm��mP��.s��(����?Rǂ�����/���>\���Z��h�C��n�&f�b��x�ҟ�������"�s����p�Ֆ�ďpz9��7K��Y�7 %������y�OJ�`��	�!�9�ezT����eX�F�B&�D�6e�TK��z�g���6�	�,W��D����C�F��nU����pf�vx����L�R�m�:]�����(v�u��F#�Ji:e��?'M�/�}�w}0����A�@��Ыsj���$ib#<v{.�6,�x\�GQT���TYIX�sc����b۬�v�9��P�l�R���`g^:��nv��>��q��_�Sʜ�����Ç5\�ǁ�moB˵����HS�w	(jVoñ���>˄`��$<P�MS}��
m5��5 �zD�	`�t(���B�j���� ("c�.��!@�>E��AT� ���	JT���74.�p�$�B�n�I���v��ԋ���m��gD��
c�U#��$��xȏ���p��\�U7)���$��&�1e���^B����ӵ��kT�R)&���W����W'�rW�Eߛ�4>,�%�C�o�B�Z��\@^��l2��NFj��٢"�	E��͞�@�T�����ǅ	�����{gF�� �ߏ�U/{g Ǡ$+���B���?.�:��G�S�*�����.�GA��'.��bI����l??8�Ep�Q9�2��~@��ZH���!:�Fxr�g� ~���\𱇑�N�ξ�L�T��KT�l�zI���6.IG��_d�i�q�z\sO�6h�"��E*v���j-k�`8�]]��avYʊ�_
�s�g�&W~�!�ƿ�x�i���o0�D�Mo���E.��Z��bX�L(P{ۛ[ +���u�#^�Q&��n8�>�;�}�S �̢��R�:�p��m����#��4���ڟ#��n��B_�<����K��z��Cg��Q�;oa1���5��B�����t��MF����c:7�ЊҮɃ����";aC�2�W6I�IxG!�?r
���ek���R��+�[�N���R�������1��Qhbj��Pt�d�r9�;�d##}�n;�B�g`��8rP!�z��<�ۆlw�(K7��X.�!�!L��&�Byir�o+_պ���(S�4\����c��v7�7��8����ܖI��+�#U��g���� 1���Ƽwzv̐>��o����[ŃK=+Q��+����Q�!Q�Eo`�ok)oU������]~O�6�����ْ?�~�w�Օ�m����x/ܡ[� s�ش0�1�I�4���"D��D��3�i+����W2�ɽGS�� �o��{�GQp��r/C��o�^s)+�����RJ��{��{$6Q��yQ��M���i��U�:ޜ�O�y;���&�[�$����U�{�܋5�Oۉ=�c�ܺ�C���5
�.�Z�O0�㎿[�1w':�f8_NH���W�������%zlF����ǋ�	���b��zF���"�U5p��[�k��2I>^(J��ɲ�Z��q������^��"c�3�\��N�˧a���H�E�U��CG�-�����T;r#�6���#I�Vxk����ի���X�=������4�����)��r����N�L���8�����:c�.����ZE7�[�IA;hg�(0�RK��T��|>!�/%�К�'�{��<����#Q+�b���W{�E�춂I���+Q�F|=�,r���a��ϫaj&���7_ �*�|m(ϫr��������K4dwQ�*~Y�e��~aw%нFI}{<#ȏ�<!�Id��/#ܪ5��d���<�oY����GP;� TS�?�Ҹݕ�žֹ�rAF��d�����Q!��V����s�1Y����u~�BeFA���~�|R�׮�e~�$�a����A��`�x}b@�x���fq	Usn�����M�!�ooe��*2(��ɜ����}�2����5�b�5����o��8���y��,��UD�Af�E��_r��8���n\��x�H��G���
sQ�����ٍ���&��|�^8��]qg��C���g�b�6/Z0C�ܸ�4�����f|ș;+7=��jԇ ��tل�D1���ZFh���L���r�q�&�[�b��E�:>��C��(�<�YYY����u[�����
 �-L�z�z�����C���
�ݡ%'�c ��G$����ڬ�_�)%�EK>���5lʎ0��Nm��������d;�x=�2\.*�9�8��|-��]ɡ�òc<�HQ�~e� թF?�H����;F#��wJ��a&����e� rEl+&@jQ'�kr�����N�ZE�1��̀c�Y�ʐu�.q�']3��2.u\q��}ᵙ����P�L����-'���?��;ߜ�NƐ4��n��k�٘�>AA���bį�\������ �Hu�c���Z̔�2FK��3�h�+���Mɿ�ޔ8H��6ȼ�s���-��Y�v���3�C�q��|J�����J}����[������,!�?N�7;�<���t���K�p�����R�J�������
�1�.B�w@���Q���	�կo���S�⬣�o�~k&�bI�-q&���:�g*M�����#%x4,徸c�K��\z�w�2��3�cu�������0u��_��8^�l��;+j�CVjJW`Wٛ;���+e�S�
 ����GuܚQ|e+�(@�S��ڦhxW��U� pW���gLl�+���:�JW���7eF���M?���B�����o�/Y�8���0)ST�;���^�N�f�b�K��d�KH"���XB��ƌ+�r��|�>�#�P@ď���P�j�����9 t��A
��S񁩝@������A��FCӉ��9b+�,�"��ʞc��-��J��2�|$#�V�6+��-����Al-��~����N�Ʉ韏(�d�Z�NN��C�H;�w�������� ere���B�$*Տ#��d��ѓ�ǞI�j�����[HlXY�\�y� ��z��Fv'����V���=���mS4�\�o�ZO��W���W�J�d�t4Ӭ���F�PX����.x�C�8�8�:�R�^�d��>�96�4����u5����j�<2x:�LdO�@�m3߈�Z��$��{������2����j�p��d�QO(d���%H����^f���*e�>-��$��@�����m�����ǚ���q1QF�ۭW���j4Z$J���ٳC�V�2d��/#��0��냂h���	�/��g')���J��Sy 2pĀ7(y��͂uX-�+0�Q�vƶ`��U��d�s��S,�6jqM� ]��jQ
�e�"�������Fm~�p����~u�]G�ʣCy������歌	��卡�\�}�'Z�~	�)����`},�>�iT'I�����煏�����0��UPk�g��aXT��SD��g�Y��!X�.�J�Un����uu�[!��y1(�$كZ�9&���a���UԒ�݇҉a-�=P��b=�?W�{��c0/����aڂ�Ҙ� OA8�������%W5�`��l��|;T���D\;!0����V���{�#˿�W�a��=����T���<��;����*��B�-��j��2�����$:$�5
2E��"�w����Ȇ Oif�w�-֬ƕ�6�aO�6�T�Z�m�\y7��Bs�	mgڣ���
�%?���G���c�E�u�Sb��{S�S�F]��k�m|u	.�KJz7��>�����	��[�q}0���¶�<�?�X�vA�Y^��i��tgf�0W��� h�	���q�?<ߕ���F��p��LAL��@���i	<��QW���v7�C3�'������UE�DI���9ʈ1p̴�_�&�9��p -���&�:����DWa�tX�l]x�a�)��o��!h���ڵ�{��Tlt�c�]\�����ީÜ������3�D�ɑ�*�x㞙�"���[��OT��3���Շ��iwsj�N��4Mnu�{iz�촼Pǟd^�5SwD���pg�BL�I[����w�N��
�J�`>�ӛP+ o|�v��b�^��Q箻�ƍ�q\~Un(��	;z0U+��sw�Q���H�m�ui ��uz�?뺽����R�:�K#��0���#ē�X��8�}��G�����⏘�l�Ҟ�ag�y%��7X��7�W@�J��u����r�^�|�,u��dd:���r.c��#r?5����4��R��}�b�(dW�ɟW��F���x�Ja#�_�r������(���Mb��ߔ$��sA�q-�L�~��R�}>�R�ϐ]	τ~�M��.\2��=}&��@��x\0>-�3�#��q��cNC�kj&�lb�5�4M��3ʄ������sI�D{T�V�כ��j�W��C	X�M�m��D���B�Q������y;�l��6W3ȼ��r����`���^_ܭ���}HD�v���7�:���su�Y���������<�f	L&�a��{$Y�(��X�� ��:�=4�Ǟq�{t�cY�#�2YoI�O���uN�$3���aZ�2k����>6��41����9h�/��T2R��ޱp-V�\��i<�
z^�R��!��r��B+��H����"z�d�u���/�z���(^4 �"�;S��ς0lW�����C'�s��FM��ڷ����PH΍�n�E)ʕ��G�6"�*��)U�fՒl�?�$5�
hI�br�{5���r^y �ÿxS��m}c���z 8�A�s���sTDa��襁C] �8!pҞ��F�]���
�+�3��Y���W��[�&�CG�]�(�Gy1���NGh�w�E��0�S�^��9���C�H���9��p\�r�Iw���`$�}[M�29�ע�6+r�"[3�J9//��<U�����OD���./�`�is�S��zc��j�V���A�b�1&3�S߉� �h�����'E����<ڑu��:�M�E����!�?��5�O$���%wh�9ɇ��c�g�R��ua���/s&�p8ˏ���`7��l�V>�$���e�2�v
;F��H#�$I�(,���pi�o�lp�"���K��!@hβ��4
g19���O�ө� �g���!�X^�	��1=�͛)�e���?\�-�s��.u���a�a	�Z�k�	\�UU�,l�ٱ3&���%��^��_汹G��Y?Z��Gq5���:��$�)5�{���7��n��D+||O����7�s�>G5�v˟�^��{U��B�4��Sa�S�8d�7O.���p�!9ST�Kt|��yQ���D���},�h�<m��?�,&ln�"D��Y�gl �<���S�+����tڠ:�.��@&E	��2������/(�3f�<�tR���%¶^��N�o���!�8հ[@��et�=P�9Gc'�8\��j��b7~f�3F:����l���@7����ؗ� �bT��J:��E��(�~��{�CcL��l�Ó����~<l�~��DKt}����?��A�7���`�?$�� �1�e���D�Cֈ� y�+�/0"\�A	�[S�[5D�滅dR'�ȦQ�ch���?��:)��(��z��Z_W�����7�;wj����_b�-�HI��a %sLy��?��m�@B�A��J�5��x��=[Y�s~頲YM��c?2E�����uh{:Eb�����cp �ʲ/՝d*}~��k��,-}��f",�j)(_(�#U���[�(� ��YN�@�/H��3Ls��tF���!.���k�1�A���6��W@�dq��~{	;L���M4�Q�@:�F)��u�)ӛ�ןO��K����f�u=�zȈ��BK�K��?5��9+���=i3�(����f��|!�[m� �8?#����{��	ի�o �m����h:A��Hg���W��<H�qB��ա�My���^��9�b�x�a�u��r�2�:�5���1�R��ϯ��c���<��U����ľ�<m�h���z�7�Q��� ��ݮ������<�CS�\ ����%������_���Q����p'4��Ix���U&�������+��%�8T^|k;-HY䪩�"��j�����	�oo4M6@����g�P[}W�@�f	4)y�Y�U�7&�!����zh��.o��k��� Б
��V���xǀ�i�����ѠJ��S��ϐ��O&���s穻�z�+oǖ���E��)"S,��'��^jd����Ư�P|�;x��XJK��?�d+�%l��aA�Z�ќ\�txT��ZQ?�B�#� ��v�w���
�[�Vvl��]����o�H�����A� ����!�j���LBԦ+)!,��C$�\��X�(@p�g�f�Ǚ�Ƈ:I����曡'��c�r��К�x�F6�P6웉&��A��[����h1I���X5
�h�"�լ������lY��������9w�8�e�����m�WU!������-����t�S�9ߛ���
��"�������tY>��'�����Ic:�ج�`kx��;�\�inl����y���A�תo��G�C'n�)S���	��~oP+v�pG媙�)Bkwu���h�1P)$cG�������������S�9.���w4��:ڻK�E>4�j�3j�L���?��ܘ5����'���:��%�h�Қ�A"5�}�� ��v���ȏ.�H�@��$jDI���J����7m���d͇8����l�'��_���7X�Z� ��Q;2ecy��,h��4��x �͚���S[��?�����P�@�����+u,X}�@eMM�a�~R����h7P�+�/@�Od�� ���Ms�6t	O���94�Үo��~��q���S��|��g����U�U�����m@��Ο�h��\�r��R�	�õ$9�zP9͇����;v7f�z� ����h���tUv�~/�����j�ؑ������>1�,`��'�T��A�_hn꫊�1��/H5ʫ0ׁ]6�Ǐ�W=��bLs�K������{j�KF[����W�~���nބ,~wA��@ZN��Պ�/L�R�r<PME�N/�E�o���#H�{����������䜷	.�g�;)����r�};���&�Q���]5%)�8���#)�MK9�/GeΈ/�~��������2E�D��oS�t�s���iɀ�*-noM`�lRCO���D�޵<6:(�r�,Y� ��C/�����gHk,GWVq�r %	Kvl4M�6�!���h1/C�\ݿ�[	����D�g����DKV�V���"_�N"%�\����6�F�W��%!�b���_Έ!�����\�B��3�e@�	� �v�ʹ��(x3�g�ڋb��譑Ke�;d�z�韐�ۄ�5��W���4�nO"�&�O�Du)}ą����_f��	��׃�-�OL� ��y�3��7�i�(Fwv.�\��2G�s���=��\~�J�:!�X+��.�xOkv���=j8�� �Z��A6_[OuR~����Zע� ���I#��ܠ#>��#�ϭF�J4����^�+~$��#'<rj!�W��	���H��٨���O����i$ɲ�>aN$ZqѕP�-�(�e^���	#juF?��928���ɾb���b��w=ofU�sU�b�j*̇�(�=�h���O��٤��}~M���f��>���ҮH`?\��t�g���o�O�\�k��
�������`BH���9����]q����8�"��NQ�vyZ�=9i�s����u�-�k����vw�Nr���� �����J���MD���$8�qF��v�$��*��\#zY�71&*�cۥQ0��oES�G��l�ҍ&��\ڳ�\����U��RW�j�)y��F��&��2.�'��K~��jo�`OS�e<��iiV��ŗ��zٓ����ʝ�53y1\FS�FH��%[;�)*�K�7^O���Z�G��D�f����'`<#h2��-T�#�dY�B�B�
�;4;�=sx��?���px+�0���4��Ʈ?���\1�\�X<����J��7ѐ���	I��@����԰��u�^�}%	Ԟ8}[A��w��(��X�+k�Uܬf*#q�}d	WG�Jq�b���\�!�� �L�F���.��Ǉ��y�EmFy��ԉ����<����ހ����-0@�z"ek�Rk	� `Q�D��-e�-�\��NFG��Bs�[��gj l��T!'��� ��?�[ﺂ0�G�ܛ
� ���x�`(8�y�������5�JZ��M�"ⱸ*��� ��9KG6�;���`�&2�l+������r�,�Y=������_zӭ��n����r��O_yYK�t���/@�{1����cZ���)Ub�B��<�zႾ[���#ӋO����e���������H�����y��h�B>�'�%���E++���'�r�bOH�=v5$�T^��M>���ø��ߎ�X�.�bG<����{տ�WV�R���ήetK��]i��_�E�ŜO��k���hw���
c��bɳN[�M�q�����TVh>��xu��^�xu�h�i�*5��}x���L�]쏊8�%�a���Р{�����=�O�y���A�g�]%��'nɰأ�D�a��mi������N~�9w���ٖ��71Cf�vho+L��z
��D�5��=�?$BH�}iWF�
��ٿ�v�.(Wr,���0�ah}�~��_F�n�����f4o�_4�'��Vs�#FO��hq�Y�c�Y͇M;պ��6"t�E����
�9�$���Ti�-}s�<����S�_�wD�𯬨ssQs�/��8Ϟ���ڒ��XW��t´-����!�I�}�E^�<�i�%���&��f���J����[)k�g��փ70����G�{���Ӌ�ϰȓ7_����q�xS��T0�/�j����'�L�� H5��f5e�X�0av0�:.�|<�=��H�O,+i*�c�}��,[j���*V�ЄH:���dX�{�%Q����is*&�/ѧ��`���a�����HC�bgpW$���a"�ׄ�{��r.��K�8���E���>�nK����+��!��~�gH%��]����,���ͭ�@��O-f��+@l�S�a�^�fJ&�u-�tp��
)�E�!9�Y����I�5�bIeBgeQ��U՛���m��[/���9�q�y1K���Dz�%�+1)�!�럯�F�����E�Ԙ4���ۇ���7�<m����9z�rY�'����@ѿ֜˾�"$��/T�6��1�u�D�_oH��
:����>KS͐1�.�Y���zqo㹬���g��� ��_�1�g4�dq]6�E���3���ǭ'�X�g��dL|S�X�D�wE�5�n�E��6Ѳc� ��_I� ��?wu,= ��>������E�f�ʡk�L'r��EB��D�4�H�ڝڱ����u��dA��%����u6��Ѩ^Gjk��U�k~�ri�Y��T��(V:��\��(P����L7��ʷEhIl��FƑ�!՞��@r�[qɽy=.1�`���T�	��0Z74+���#�;=eea׀�ݼ�nxhk�|������s���!]F8��b���>�3�Rf,U�:���{��2�`�/�G�y\���v�uӜ�˅�v�de��Ad��I�
�zM��
�P!Ԙgb�wa�P�[���'�R�L����ԕ;�B�& A��D�6R@���Qx=������6�d?����b�J�4��l�j��0���q'K�sUU�6t� Xi�V�Q�f����ɲj�D���/�
�J��[�~��x��{Ęm�w߷+~��;ߗ�w�ݦ��c�겷j���𞈵��YU�FJϕ)���p�rĦWYڶZכ�!*!��K%-�
e�͵I����2�+v�E)��e���l@�J+O�2=FQgƊ�VK���/���'�� ��!h���I u��Z?%�F$OWy�c�FK��:��2�Ծ�Kτ��i.r��{n}�-�gR��կ��wK��G�@g���-h ��*����h���� ��.�� �7�1����e!����wu���S�Mv�25�b����P�Uy0а	0(��m����E�S����r��ƪ8J
�ʴXƀ��4S4�I�� g�Qv�KD!��_y s����ҍ��'���ħ�l<�"�pĸi�P�-�!u%�txD|�a�e�%:�Bo�I�O�Zp��5<���"��E�����MQK%1ʈ/��@)�~y�x��an��_��^��i�Ӊ�Ȫ��W�E6�5�6g�
 �?E|料��7W�'���zn	�D}��/�K讑X%�:�/��a5?�S�4�v��)��!uA��� n+��Ƃ��kzXc\.���N�D��O��P���\�Z�;{$N��XiYP\in.6��Z���c�GP�U����m�
�x~���w�U��g˹��+P�Q�`	�i	hӑ_cmt]���0ϏD�q���'�p'`���*�)!�������p�����2�q�8
�%s�f���i:��u����j_�a[E-�1r+ �a��"�ۃ�Cgj�\��*̒wn�߉��8�,�������OG_k�'<o׽�ZcȮ�˛�+����Vu&S����ڸ��>���">�:G�Vۑ�ξKH�u��|�*��h�5�����8�E?�Ud#�D<FN-T�Cr�����I�ϖ�-��)a3s�3ɝ�Τ��?A1 ����Q��t���_�����P����%�q��>A�jsҽ �/&]pr8ƽ�l���ފ��r/�#	?:�-��M0��%>{��D�,����pP,�c��i��K#�$:�0�!�5i��e�=�N�
$�5����=�V��ג�됈Q,or��pj��RL��~�PNɨ�%�K�7�!��9([yQK��x��b�F7��p�&�o`>tg�w��Gԅι����q���~�����{�8���m�m��4Q�C�sM�wFn��Z	0�	
�F{��^q�]A��8�㌱][L���f����XS�l�O���-�X�;Qq��w���UEjy`�Z�/��:Go�W�^����q�=X6]>!����ȩ5�]��67.8:5�fdV��E�`mb�u����0�s���:D� ɑS���(�ψ����BtD��dM(m�z��-
g�&�|B�#�$	Z�ͦ?����4�4]�ޢ��uJA�-�1�B��:���1^�5:��4����ņ`>*}�Y��T� ��a=Ǒ�4��t���{Ds�D��b4R�v4� s	$�~`3���득�~Y�K�]�a�7����y�}5=28��e�E�?m�Kq ��3`�4y�4��Y�FZ�ҝj"͗3++�m�э���;�-�n,�c���s�:~�5�v=j�*p�^~.�\x:l=�3�F�d)O4��7�[��"Ƣ�	~V��� 7��x��w�Dk����d-��e5�ix����b`��o�]^�� '���~dJU�
��-�� ��m�ŹZv$�-��v��lD|h�����G�:,�([߆��N�� ����YP����,ۏ2�@(���nsikO�����ȋ]C�K�@V�p�ye���0���ک3��.���XY�S%`��=I7�̱�> ��8]�b�����/�я�v�H�m�EcOyP?w���	���q��^�A�㫷i����ӊ�7��($�a�C�����잔Y��m����H�kV��?^h��/��zg��d/���f���iF����p���qH��!y:JP8�d���0�l2x[ߴ�'�I�9^,n���K���=�< ��R
���A���5�颢�h������,Ya�iS�F�*6Z@NKY��� /���l���F�~��wX`!YP����C��Gyv]6�<i���|]��!~Ӌ������h��h\�b��A�m�*+a6�kj���e����ק�5fD&X1r1���;��q��;�	K�(�M�o�t�u�B��WM����� ᖘer��n�נ�%�@��h߹?�PE�AP���N\�}�܅�FA���Q����fU/�����+��j-3�����P��03G�^�$�=zGh�`jP��]kְ� �����N�t�����R��+.��A@9/vڢ��u�|ϓ��7v��]���	��NwS�yq�y�Hu���S�h2�-��Vi5+Y͝~H�Jb�*�@���O%�@as_X��9p��� ��qTA�����9��s�"�@�W+��C6n-�ճ�r����i�"㋕��i��ͷ`O�������MgA��vdY�Gɜ���5�	��V&�2��n���땗Ǔi
}@���c������sKr���v!�nO����?ko&=a\�
tLz�e|��/n;���W��c\r��pg�\�	�����5���|�l�"�>se��4�a���X$���B���Ucm���s�a�����U��O�x�B3��iF�A��ѧ~�P� -���w�{K�nVb#+�!�L���g��|�8�S�8��b��0�������˯x�_=#���'(��������W�1�/��`�u��^�ܜd�h�V-���Բ�?+ 6%��w�D�,�Qz�`%70%�_����%�Jh�]�|1	'�&�D��xj�ܳT����d�o��V��%����=7x&�z{����K�g�� ���v�3L�q䱒���+
��[<������Ã�B6�*��-C�iOܫ@�;ݠ�+d�ٞ�A�5ɖĜ��'�7j3|.��˦.���B(���Ϭ|L8uQ�4�DPe� �Al���So�UD[��Hl�v�
EFG&�O{>��������Q�1,໥5�NO~pA�KZ
�߻����\�&y$����>�Y��8-)9� D�Kp"Q�q�X)��<�|�d�?яX��b5>+���p��å �Z�5V�W'�L�z�O�A]���'
���9�4���<Ϙ�1m8������o
�Z5��U�r�I/b�fԯ{EM��|��T�tcs��o�����������WH^��ā,>�����N�sWwE���������j��h�wY-��t6$7�$t�	�ƍj\�*�X��`�#��"��b*kG���%��g�`󩰝�^(�^����uq���/*�k{ld�b�'Z� ��	p�mr�^����9=�U/�����r���������ݐv"���V��~N����t
>����`$���*�{jA}9-gb�K��Oɚ�w�:��)��;$+������,��WM@�%Y�r^S�l�$Ym66���)n�RX��t^ �&ަ/_<#T���iA�#O�4�b~�_�Wܠ!�Q��AJN��