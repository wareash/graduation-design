��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf�&���>b��z�P��!Y�������p*s>�+'��g���� ��1��yaY���X��&/Y��l��{B*Ն�����I��W���9����������˟ ˮ�9��~�s�M�?"VYZGЊ� ]�}�D+���yniW�o��No���󖿍߾�c�/��W��"�2�˿��i��W��w���f�Mݚ��39��w�B�%��C�s��u�3����ށ��fn?S��D��>�Z�ۨ6P�td����fJ���w��s�#�����OσR�e�]��"�p��k�c�U�uj���*����#Z��Q��N �Sm��՚OO�!�O�Ӎ,��Y�~�Ò�"�O�(L{Ӭw�w��ܞ��L��{��Y��vn��,4�+߃]'�uY�&���VW^�7Қl�mw01f�P���8тN�:��,X>����ؠM���K�T��`�FҤy��Bj���-O��Bmkɵ0���Z 	N!쵀*�o�����|�B���n�㯳HR�S�V�A'�Db8 ՗�x�:'�������hm%�K>qa���Y�wM&>�&_s̴��w	�L~���gRLk��Z?��+n��"
��[3)qٸ{���}�i�<�7i���"܎��k���fah�v`����͢q�?z�K�5�F=�I�ͦ�>^S;�t��^H��hh��(�qL�$_��J��?�~���A��]V)��&�=��������%(�oTbR�X.��	@Q�Y0�@~�6x@��F0�ivZ�*�/���Z�,���4����052�a�?�fȗ�w��%,�Yhߪb������8Z����,�U��[���=>��!q����M�q9`P�
��7]\Ϯ��3�#���0��9��Q2$�VDQ=�Ã]ە����b-g�
"����� �eC�bUx�D�	0]�Z\s꿷�i��Q��{�<rqH�)O�>�@� A�;�o�Nɲ��gfY���G�J��, �#��4��/uƦ2q�޿�͎Ԩ�k���"l�vt������?����T�hqh@LM/"�=�@x���ud�|^��AT����s+0W���4�M�H;ĵ�H^=i�F�!��D�������K[·f�|��۬F3v�b9���Z�OP���9`�I4�z��V�z�z��B�� 0Kف�MQ�W��*A��T��Di���n���@����)�eϓ�3���7�����:��l��<bEIJ��9%�ʥѽ�d[{��v��B�,�g0G�t�#Z��q�3T�w����t&��^�Je'�<�݉O��H�I�M	�,�d\��
�?K�S4�� i�q��<�8(U�ɵ��� �rY��q�`�~zÊ~;���y�Z�����ݸ��F3�z���]���o�2T��1�ٿ�o@W�\ʕ��"MJ57~��.UlT�Z����"��^���w�N�򤰅f~�TN�[Z�Ȧ�.@�r�p[SdR<����Pt�qv���z��u�F�ћّ�Gh��5�`L��rF=b�䛅F�V^�Ol&���Jv��.�Rۗxy4��� @حH�O�'��PV���"z�3źT&q= D{-���ߥ�˕�4����P�?��9�k�2�d�J�L#sx���.��5p5������ F���R��Du����=j5���i��;s"`�/����x��r���D^�Z(0@Ɣ��,<�7$��Hbނ)���"5��a�`�!~A����c�$��f=_<��'9��{��+�c4��;g.s70� ��龬ӏ�9##o�{���>%P��Y�eh�t�E�P�zn5����L��y�X#�9~��醴����N�:�E��������~å��L�:�7��М��w�DU�2s= �,`���Q�U֎�-E�ZA�`���T}��t>���d��#�I��)�Iʢ]���_[Y&�F�.1g�kL_@�-����5F2ߵ��ھf�M¾�������4���5? �����p��W�q,��lȉO�z��=߫k���V�d�t�xB����>�l�t�&���!����bW(P��2D�6��N�ͨ/�P�'�	�8x��(��Yo ���%2ʐd�!����z
�B��m��ԁ���
��]u�V(���E��B6�㮴<�tY\ma(y ��p���9+�!�gG�0<'*E�v�Dj�B7�u�E
���ip#!#T��\i�X%�9�W�n*M5{D��L��
s;yTz��%��&�
Uޔ�HZ��?�C\�|4xƅ�ʻ(%�(m��-�}`�)�G��IW�!NFd���ZPԕ�N����5�]�d���'���_�N��ڡU�p�ϋza'�2�[�#�MXk,/k�4�Y&�ߔ�]	���
}�Cd&�t�(ԅ��	nQ��@aX��[��W!�!�PG�j�6xݧL�6Z߸�_z��T������:�:U
����P�Q
�&�,��zp�.�n-v3�hBRu��Q�/�O�PST��'��*A������iM,u��R�\?�����W�� !X���E�rg��g��� ���[jA��Z���H4}A��}ǔ+���͖��FC(9��G�h3�_�;�L�Q�*��؁]a�C=ͩ��C� �i��k7�]l���0�G|�I=?M�e��ֿ��Z��q���P�����
 �D�5s��ѷ�*���G�1]jp��]Ԇ�B{�y$��#��,�}NqF���Z�I�^`�r�[�<�Vӄ���ݔ+�w�8�q���6�U0u��V�F+�T����q��S~��Ѿҍ�CV�X�,�z2�s�p�(�N����(Y<-���c�c��fzU���Pu���C��=�LT�.u߭��ջ�/��|y�s�;�����*�HO?���~�[���?5���6Tc�s1Tgb
Ϋ�����S������УfU|jV���:��Vn�m=II<b�r� cp�w�;P쮈��~|o*���fBw/1��T���Z+���kfo;[18��˼nW��Hr�͈��,n[���J�n�+��,6�|���c�'�W�Ӄ���(#zi�5{�zH���8��z�'��J�⯳ �n=��kX�� ���$��4�Lݛӊ��O+���cA�l�I�:�7��Bu�`�ۇ�<i�?�;}J��kr�i�}
[N�e;�� �|�~�+�6�Š,C�/|Cm<d�%�_'�̲�`ć��i��Ba���6 rBT��eɪz��*HuD [�6�#��M�S..}��7xJ�W��<��d�Z��A;�\���ʖ~95%
3��O��go��ӕ����Q��t�[?R;a^��j�K;`^�iX }�e�S!4
V��H-��ͰL,�Y�ݳ�*���CX��.;��")�G,T�g10Rįj�� '���Ќ]S����9Iz��&?	�rˋ�}���׼	��3�o*k2��zimk�(�\�C����-Μ8����B��ig*�NE�d�~����r�_�`�Uj�c��`�[���>�N��l�v��S�v[s�be5����X�jFG�Ci���Ȁ��%^	�]������.#'T��Č9Z������}Ӏ#��āA/�;�@w��k�r�G3_��Ne�5��uhj�

�+�����~$k��4�W�b/��T���ګpRhrq)]G^垶�d'���y�U�LT@���h��?ᐭ�S�.�ID3='�:��&�霳�ƻ�����,C���5�1�;@�ư�y��~{�z���Eg��=�/���}����22fCSR��+b�3]�M����^{0D�fUG(󬄾�̀�"�U�����*T<&7�އ�g`"�'ך�\J��(\=!{C�e�+/}���μ�I����4w,�_���)EW�S~�W��<�e�P�99�T�Zi�3x�+���ɖ�+��ÔS��U��3�wxU�}�����[ۡ�8$�=�&��8�U�@Ԡ��B��uC|��p�V D��W�Kc�V�g]ؙgXeHcr���6}8�*�bz�i9���
whc>��y:{�V���J��UrG�2�z;)P]�3�0�nh �!���7����ʟ�J�� �y�B.�'�>����4�$�,4@TO���L,�*��gGn?_ݠCaȂ�~lWn����{��'f��]�?���d��c�J�{� ��P ����΂�c��X9w�z�C����@z��H�Nio*�L%Ĳ��|�}ߴ�.K6�_ȯ��IY��B;�:=��21��"���y(GYo�՞�=�{�<���۳�d��ڒ�4�֗�FɊ?[ A �])r�#��O��4a�g%T��懸�z3!�z!^:9��ѹ����3
�4�i�h��ʇ���AF�Z��2aF�\;n��㺊m�f<>��4��O�J[>��b�yH��8���y!/
*<ug�4�縘}���k�j�]�T���pF��*8�����)���.��Uws� �*9���I~��y
���_nG��.$��¼�G0!��}��2�p�;��u��V7;��z\ׁ&E��e�Z��¾y��y{DȣZ�o�������r�<�"��FD�?��Gҫ�Ϧ�C�)*�L}�+��"i���g�U$`Ib>p�beg}{Aq	΋?C��C0N����x�>R����"͠��IEJ����kt�)�8��*w�Is�z�_+���s[x*B��iK�˔$^߯���5�mk!&&�����?QÂa�?��ӡ5�	�5��^J�3@�
HB}����Zx��BI��m�)�h_���oz����nK�@:z��<M�҄$�~'}���`�`3��#6V��N@|	/�&L�*7zx%Ev[i�@D�*��$��t�ы��P�Ts	���οR����X}�Tt�:P����_n��u<]#���m�.B���׋t����{�}5�?�S+�m^�(6c��&(=;ұ�ʜ.S��g���?���4-7�-:�(���ս�ś��l=a7=�C��/@<����޲y�(�w�C����)��2�K���&;qp�?��_[�qq�/l1'�b�B�ޞ�,5>�Ƚ�ƝY��g���"W�g�YOi�����x�a��%���q|�޻�S�è�Y�x��m��������ªF_c�q	�k[-6l~Ɨ�ͫ�{���#V=o�,�ф,�XT�@?5��n��N ���B����$��0���u��z^����w�5��KH�{��gKR���LAͦ�y+���xᔱ�Bz��S�H	y��!W}+,5��Ŏ�6a����Ψ�  ��;��0����? GF%�
?�oF��C��ԛ�A
'��#����[��مW�l˘������?���`�"*��h\�Bt�KXl22d�xm�C���-�g@[I�E]˷��D��Ә9���!�Ȭ<�jK�ڟ5a����"�$�!�c��`�ExN�c!o��e6-��EF���AU�����d$ud����@�I��S�9XSK9��j����ǈ&�4{��2r ��W�Ք&��<�WԀ�
p�o�}p�AߺH�f�k�z�u���	�y»J!�#�F�z�ށ6I����Y���}4��C=.��eR��޶��19��y�e�h��e�k.[�D�Brc��*��mV�i��+�kFN�o��H��e�vl"����9x�.�̋>=�O|�����=j)Ħ���כ�G�$𮨅1J;�p�4��/߂h�F����v`]� �K�uެ2��Y��2;,3��e��=Z�cz6�1x%N���/�V3��]-�u�&��֖�2��恔Ņ�h���Yf�����Q�,`ZCϰSfz �3s��E{�j�]V'p���#κFYc�	�����y�αh��K��;��*="�2�;���՜|�q�-�oJ)	�}|�Ϻk�|Ƣi@���}ؼ1\���Ss��ةG��E` uv�I�hz�Gr�Dr~� H�f	�s;,��ʆ��D6q��i�+���	��v�lL�IW�7[>zP��M{���v�[j��.%�}�&�PB.-+8��YZ�>��2�^uUev�k娽�#b�X�qD͝i�G�|�n1�0a<���0徙t�V,�+S�HN�T��lg�x�g�HE-�Ԍ��t�~WAi}pʳ'؊����i��9�GePP��3���xq
���`�7,oM �X B�T�u��8����c���S���[�V&�Mҕ%�D�꿏�_��y����ٹ!�Z���K(��m�u(|�<#Z�n��H��4��G��[����,`n��+Qڰz�f�5gd2A^�p6�;��S��)TH;:K�j$��#�G��a$���)p"a���X�/�"�-�b���C���`�a0�ј���+��|>�&�������4�a������2<s�k.�Y��'v,V��(-J���&��