��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>%��}w�K�
y>F�GϋUX=��޲z Xs���rf�-*f�ŉ
���<���Ci;W疭_#CW��RX��:�g��^��큙���W�o��G��?>g��+��,^t��ϯ�FI�a�,����Ƥ���023�ٗ��=+E �����j�t\R��(��l�&���I\�߾�x,���7�Q�� �sz��%�d0<�M�AK|I��!�`_6i��5H�]+a��y�|h�%�~\�������y�Ov��������+5ӹ��i����B��smb�2��=�������8��_��ZHBs�k�T:f5C+B� �a�Ɯ�1�A��}W��C�o�����Xc�:�?a����q�^9pU��Z[+>�5�y��m��-�(+sΐ�P�t�a�-�A��*uxpe��VB��gF_�bx;��^��S�������}_��P����V��*�Dw-�a00_�6h(�iw4%�_@����p�G�ےpQ|;����n��t�źO���C_�	Z���:D��"���a�q����=M���w&��k����GҭV�$��]�V�*o82���ҴpZ	?�r�r�(+*�G1�"+�������4��e�>��y����i�궟@�<:�r��}j���9�:)�;�	�~��4��p��������u���ӭY����+���:"�����;Eړ���[�ZV�Q.
/�2|�\Qx�2��`̞�l�V�c:��M!�E`�-�f��M� '�* A�t_g{�����$r�>��6�d&A����z��9�FqP�[`.�P��=�%z���T�fի�0�a����9��'%J>B���կ���/�g��i�Ũ���~M�"��$����[� ��1�v��D�D����/!(5��a��֦�;J$'×+x���f�ڡ�'PQ�8�t�+.ivз+�JCj�ۅ ���DO�wS5a
�_?�*��#wYA�H=(��_f���rm@���2j0��V.CM&�E���My��?n��h*>o��8����3/?�Ǟ�	���3�h�C������wBhe:����i�(��ʆ�!���*�[1�n�1~���7.f�I�kn������m��V%q��s���w�Y��ĕH�Iv���=Z�:�׀�\��WLX�C���)�1��)tA�#�5oJO���^�!�1���bS�Ԓ�� fQ)����k+�H��dk^˭up�T��։��8�G��_R��eЀ�@�|B�A0DWJ���l��y������إ5B�Z(���Ծ���?����%�ռ
�k���f�W	ئ!�'����9��w��2aF�Q�ʨk�����fLsu~�)�KaC��g)�3B�u��t����ႎQ�jv�\�a.\��ۿR0|[گ��s�* Dt�ؐ���٨����EU,�1�je�]���<t�'�fSҟ�� �gY�xH�(Q&?򒼪�>��W��$�� y�ׅ4I��Y$���pod�^�3��x�f ������{�&W3QF�֡Qفx�s�.��i�����4Y�D���f�D�1�63F������I�T*�䏗(���/-͵���H.+�tHC�we���8=V��L�w4�秐02�P�h"^���X�����u�:�����c\��ȥSB�
[Dl���S��:�~V�%R�n�8�۴g�cV_*��g��pc�/n_��"���h��>��� �Pʳ�N�Ll������ſN�	���+�<�RU��O���'A�8�ϧ�jD�r����.����P^�wg���x���w�9�G�͖�DJN$�˂Z1�4�|�&�(Q��B�l���4��~5�S(ltI�']m��rA �B�8�*�C��j�A�f�\����X�aJt �<��M�E
[J=�K�XPF@m��i�K��ps�V�q4��-��~������W"U�P��xx��2�/�V���Y#���W`G!�O�@3h՞�c�ό��u<Ƣߡ�굞/�q+���n�iB\2���kJF@ǁ�����fi�����m_$;�>�z"�ΰ����vx��0��*�i�F^����,����t�S\U�,
��q�w ���#����i��#+���x��i���<N�d3�^����X�WX1�2���$�p��  Wn���N��,PQ��J9ֵ����i�੧��̀Y�Z��T�{�=��v�IҫDL���-Ffҝ�+/�����x>7d�f�P8D�� ��է��Ŗ��3��2�ͷ����-���d�������EM�Β��Ō�=��Ê�XJ���7@T,�H�%:��)MH�Cu���������;΀��*VqH��!^QQ6����8��;U�IL<h�S=���B���a�p*�)�U|u=��
�v}����+��?R#/���0n�.���:�J5�Xll0ֽR,��4��r���X|�]�u��Be@�p|�s�q��	�\w�����'\ӝO�@�8z��OF��̾��F�J���Ġ�g{��y��G	��"BEYu�hذz�. ���-�����\>�u�A̷݃m��Ӱ �����K"}8e�Q��;�q�F��,'R��mk.�_�]��:o3�{�'��Dp�}@Z&e$���AO�n�=C�laF���u��&�����t{��A��B){w�+#y�\3�,}�nQi?5�t.ܫ���rՌf>���踣Ǹ�]d��[�p��[��[��|E�&�]o҈҃НkZI+��$$�5�`������*�G��D;\�~�����8�	<I $F������,`�7��T[���3O����qYU���g�#�Б�A������@>	�xbhS��<�êey���i�K}��!�n6�"���/�,�"��Q�ϑY��3��ط����� in��D�ѽWټ��Ӣ �u�gCjU��}VyN ���v{��!�A1�8Dn3&�� �	�Sɴ))%R�XL�D1K�O�_Ni���U�xu�S ��_�u������g#a8_�9��p��O�V��*�v�cl�V���=�9==C���3��jk��rWh-�2��������q	��ӒJ�<�Y�}aX����0��E4��aq�¶A)I�Q3�7~l����\ ��6�������G^�Լ����S�I{'��o�,��N|(��b�-�U��̨�9��;)�I1��J
��i��0k�hk)h+(D���F�X5��_�F3����/��gy{.{P���Z$QU|���K�0��nXū��=�8�U�۷pt%��C�T��
�?��7(c�������'��E�-x�,��3���X�d~c�4Q�����l��0R�%
v��ю0�>�:���*[����Z2Px���C�A�,���g/C���YSK��CaC��=�&�t��i%�~p��WK )�o<�����O-�lk�'�?��cv��*�ɇCљ�/EYƁ�Ԩs�i b���r/�X{��8���\o��H�
\��+H�i�{�51Kmb[0�'? ���#��K�&r+�,{�x=A�;�!���N�Q����=��j)e0���J#:�jQ��y�J�7c<"�II���8�kR�k��{J�XCH>���%�׬�U�t����k�=x�� �,~�����‎�}���T�'4ҽ��%�k@��C9���>���j��ֶ5bd�[�նE�1�n6��~��+ܞv�d_�Pr����Dm������k'k/ʱ©�\@���iQ1��PDVkxe^	�.0Hi��,�N���9�[p�@_zT�8J�����Hx�$Y�Ix-�ĕ���
&��Eֹ2_�z�5�-�+h՚�#A��-��^�>ES���U!��_(_�n��L�LZ-y������g��zJ� ;ߠ5��e���ɪ)��r�[�x���O�;Dl��*�;$�>�] �PY�nr^�1㍼��$���^.Zzk��`��JO��Z^��em���rQY+s��9�Q��gLU�>�TU~	�̫,�>��M��y���FN��-�'��a���XG�ӏ)��%#��Bm�dY��~-�*-%�Y���\���(F�g�c��
u ��(�p"U�>Q��G-���>- �Q��ى�t�X��B�^�tT>�|zL�n�@��:�o�_�؇)�]ck�?�����6����4�3U|�e�o���n\�/�ua��;�S@"���Dj�(��W]��4�(xi[�̉:�q�b�~)�5g�e��&����=��
�r5�ڡ�SU��T���/ἥ�3�!���V^   ��K3��V-�Z�d-�p��@���S���r��|7`y���5���*Շҿ�P�a�������Ͼ�{�u�g�C���!�9�_�N�:��xf9T�{'LT�ђ�E�h����sS�Wk��ּ���ឥ"j��ҮW|��`���<�X����EsN\gƖ�rk
���Y��M=?.�DeJVy�}L4����rh��ZUu�Ll��~�F�Tϣ��LS��Fݯ�<wF_,����bs��O���� 	+�V�l��=�
��m��w�GR��Y�j|�L���N�[.3lI,X��M����}6�".a	�k}�+�z}/Ay%��ubI-Hg�1��i?FJ���/`)��p�4Q?!�@=RቛH,YJ�ok���ʽOb�D���OE=���f"��a�&ֽG�u�a��h(�w^Q�S<^S��Q3+\Q�YO��Tj���� $X8�H��m?R��_������;#7;�Q����Yex�L����5�G�с(�|�m ����/�Ʒ���%��DԌ��n��j~���`��GYBԽ�����'��Ux\t<�6�n�Hbط�!o�D^�OX��fG�.�| WR��O�Z�h�u�x/���i�>��1Ȥ��)�{ϐ��a�Z����ɲO��q��sT����>X�S��cv�(\`��2 ��Gy�R1<��g3��#J� �_J�K'�R��G!�I)Q}�c�@��J�B�P�@������SDy�Z��0����`_�e���f5'�S�@�:��;��K����|�����x��Xs���'�xf?����� ��4jغGT��@k�YI����K��řO;��EeN��?Z]�/�⹅l�V}$ߞ�X��W��YۯC���[��X+�H^�unn������*tb��ٗL�f��b>$��^D!$��Wt�~,�i< �O�1�!��.�E{5�I��r/��EB!'C�>-���C/6��Q=C�_��M�෤G~D������'�d<N<��tж����u^�W<!��<#]�6R�X�3�D4.�[��l>�8���B�d*��{���+�0@�Y��!�o��!'3��G�N|�Pd^)�����@k�Md���B�ygZ-{zWЖ���b�*F	\�)J�fw�1�}�n�f�;���L�UJ�KY3F�|�����bȹY[؃�(�&����G�F8�H��p���vd� �^��Ir�Pi�u��o��AZ�I�Ba��9@��Y����X� �_IO���v��5��%g����ޜ��Ⓠ��A���h �ۆ{��� �L�H�7����/�!O�L9�J{�wE>h[�_lث]��"MA���Q;`��R��"o,��N��_�=s�>�/�5�_ZumH�ײ)w.��p���ë˹aOW��[n=@=�ɭ6Lx�uõ�5�7 P�r2�"�`�(��w�̼XyD}m�e*�ɬ��.ν�H�G�Xҏ�j�	��H˔�_m��Z��U���+w�,x������a:�3#�q����G�*|���QW���+9��R��H�)�'�
Oyj�?
&IxrJD�j�b���70~���=+�3��x ,�o��4MP葵5���Jt�l�%!��i=�)��K��,�N*��F�Z��S:��a�5��6�1�6#?a���Q^Y�N����Η���h����� 7�D�l�;��c�[^v�)�?-��u�`��c3�������F�}���\&`G�RЪrh����~R��<ۨ��נ�d�s4Q]Њ���q�'Ъ/��o�)�P���K��\���� �2�����o �e>�|<Cqs~���C�H�Io��z�����Zj�.�3$����v�w�A��?Q����cP.;�#�|����lW:�E����	�s}|�4>r,
�s��)��R*�6�npE)���2���l'��VI���N�+�7}��WЉ� �3�>0Ƶ��7�虇[ҟ}�� ���3t���w,�lc*z��C%P`��Pg�J�1�e��_���M�p�OüӉ٢�����u�w� `�-��S�����^W��)���1�{Zض�D;��K�Y������?g�o��=�!^%#��AFGt�T ��k��E�ms��I��í#��{z� "����V¶����v�ᦑ]V��
0ɬ�-4��� r��/�A�R�����n������L"e̓���+��2=wIJ�!�`ba��Hy|`�#��=Ac�u�΂9 .dU�R� ��H�k�Si�`. :uG�*�e6�	*"�ruȂ�O�--y)I����8L`�H�H?����p#�:v�u��e��r���Jȓ��Vŋ7�8mn�
a�z��HDD�0�W~�aol��_ě^P�J��ښ@*��������7�~��쫮heB����:<�ҡ.bu�0��,��' �,u
����f�5��N��w�q�G�����]Li]��u�^xt*חǹq�LSq��T]כ,��ω𠢿���Y���CU7���5�����IG+�B&u�E�gKBe��V�W1���M�F�^���<׃��2QV^h���x�����%Z+b�\Vs$�5��i�g�w��Tl�_�j� 
��i(G�O��Q�r02�H�m�a
x^���ll�:���nt&s�=�.�-���r+��r�������g
�Mz�Yg�&m��j:`L���Ϩ��o�B���L��u��(�2���X��֎H�5,r�_���+��"��b�!%��͑i��3��v�i��l�������bCk;C�_����_��(��\�-R�2AϹm���3tB���cC硒��b���?���)����]I�Wv�x>ƺ�G`[3c��h���v�=m�w��2���3�A�g\~^z�����'oc�K���t��HH�"gH^�:�W�F��#7�[����%��)g��� ��6�E��3�YT�v�	Y��h.���mw�m�I���DX���|��Mh�|ݓ�N��S�4�<���hq�C�[���2_���әߦ}���`R|!�t%��A�س�����N���LÞz�(��G���+A1Qi���=,��+�ȃVǾb9��c{Yn�\�ii���b���Y�M��lX/V�U���m�ꯑW{\B�3s�O	�h@W�u����Ffl�>��g�N���h���]WTP�c��y`1sR�L���6Z�O���j^��[8�b����^x�b�f���Z�w�O�R;�=�FE�n^\��n��F�X����B�m.��{/ �/>��Ѥ�C~���-&&x7�cK�l8�a���E�;�L@�emfZ0v�B���S�#���*�'�	�K�t�%�	wK�,#0�c9�}�jj�*�L὆�G���ŀ�������/>�Z�Z%�����9�s0��w���(Y����췼��o��+�>kE;��]�� (s۵ܚ�ѡz� x
L��	�G��_P}����na#��F� Z� �'@�~�z�5��A��e�̩:�h��K���-���`�ܢ`����x�o��A�Ǿ��7�h���ڐ��*zZ�̜��6��Z�S*{d�n\�y��x1=���ɡ���C�����N}h��n���KWt��p浾�`)wOM;��w}n-M>.��C�bC�:��t�^a���{}�σ"��)�t_��S�5��4���ׁ�*�����K�������]w��W���y=�E�+qu~�"
k��C{�K	�{�=M{�Ĭ�Xᗙ���[a����`�2�3��l���v�>���(68�d��@����0P��t��|7H#��~^�#�D
�]tG���3��oÞt}����:��c���H�`�u�銿"o�ti��8��7�v�Aag�����Pb�l��׃�.a�j°�B�Z@�9�,��	}����P:�z(���M�[�J^l����N��d��Y!;��}�k�`�po�|5C5D	���gw��K?�D��D"}�02�� �
 �_��!�3�K.��r!�"�4� �/,�O���8�P���As���$A`�}ٗ��p�C�<᣽�	���{x''�����YC�~�����Y��*4 P韻���w�YA�V������}�u�.�w��B��g}�TWz?=t��ſk>M�@5�,L�RƩ��6��F:�s��r�<�Z�W�v�DbHǿN���$��W�k�h�-��$�^���o�����ڽ�&����oOI��P�	ƨ"8K��pLn���ט0���3<�{�[�W��[|,�����
�N>33���� W,��H�+V��c�kDj�jʈ�zB�q(��r��Ԝ�>�?���O> 
��S�G�:���\*M�Ea�;�2g@ܧ:��G�Z���&�gIn�"i�����[�?$ۉ��̅�0�����C�
5Pk��4�0�A+Uakl�_U#M�������iTU��|�M�3�0<[&�Wߊ ߳���Us���<c����܏�Vc�޶�w�JBfkL��9=�Ye�~bҚH8������Wi�m��<|x��[����6�R�3����}@T�1Lv�SYo�-X��@_`�vN E=h�͛u~��χ���[o���ĝ�ps+���*p�V��l�ݏQ|��6�֓ᥤ�\������`���d��{ϓ�Y���|z�r�|�����y�LJʲZb���s���+<���>�u�j���u
�-ۣ��ݜI�s_�=��\���kn��l���6�ض�'m�<����eX���I�#�̋��z����� 3C5DeJ��B*�K���,��C����+�,��Ù�5�yͪ�O��)#�V�7m��q`B�ͪr������5%��	Wnw�~8 -�ꠌ��d]�W���q*e;�H���2��-eMh��N�#�3ayL��;8����}R��4Ȣtw�y'R����*��` Dg2����?⣬�>�LM��F�����w}>p�� �)��Z}R�Lw����LU���7�h$�<l�s��n!���nq[�9�ݱ*�X98 �?�e7�je̹�N�GS>�Ӌ`*��
�3A��i����#��9Ѕ�!Ð��y��@��F�\��� ���LY��pbٯ7�� �&���."gX�f_��P���X#wl�e��g��$��vQcZ����$��Q�n@@G�r֑	�D�Xn���Rc�PO�2��O��#�9�q������M���؂&?�(q���j���R�S�·���IFIY�?�N����A��pW*����Bw�'��;զ�y�ZW�q��h��P(N��~Us#]ʸm���h�y����Ɏ
�p*���K��i�#ۺ�>����wjYWv�����"4QY�����|�V_?��t��V,(�ӳp�j1�;��g/i��p�n8 �˭3�LfA֚uwཆP]9l��G��L� Xx��q�=����������p�Y,��q�;%q^׿���~�^�x༈ߝ�=���$�OZ���h�&�s��5�|~�A�Q���������8�ǵ�pe�Hp~Ζ�#��sJ�m0Fp�G�1�����Bz2[h��"�`�5�A�Z�a�~LR;�r�I�%��	���)�����V�8�w`���i�'�>���ͭWê�0k�E�����o�a�����X@0�/�~2�\��2 3������F�G>9�0]Ƀ1���躳�k�UH�q�Bw��!NlaH��}ϛ/J�V�yA��5Z��>Ɉ��
���Ä�Ԃ��B�i}<�
bi7�rY�W'�Y+܏�蟝�;]3�Y
a@��
O���G7�`�k���wC>cE�]sSZ+}6�}\�����j���7�ˬz�Q���%��(��Q�� "5�#��
N���x�	��i�-�'��,�R�+>g���W�5/���-��r��&��`X���1IG*d����i�K�*���]�O����Zl�J>��RS�[u�'�����O���*����q=uU�_�ϸ~\����r�����j��[��I�����d��x�
�i.����<E�[�T~pU�ƪSH�ޮ���ܠ�έ�)���ZN9R��wTBŏ"�����Ÿ���3�\G}v��;�Ӱo�ة#՛���zUFΦ�o�Ar��)pt �
���(c�5�grE�~��H�Y�����:3r�e�1�&����&&ՓΧSՇ�� 4�K�u��w3���@�5.��#?�}�*:��@/#�˥�bMM��;�)�/AJ֔�SL��{�f��m�_i0&�Q��Nn�6��V��q0Q�0k�	�y�h�%�,'��$I'Q�ӣ*D8c<�i8��-�y��隄R�/�ӵ����O�G��7y�$-��$��I�>Z�k��I�fj6v=Kd�Jf�=.@����Ng؄Ցm���bHN��^x����?�L`����������^ȑ�+<���"����N����-����*VG�mO_��gt�‽0	��t"S�u��M]�D�s��S��o�~���~�H�g��]�3������o8��l����Vx����Y��P\CN������f]m��7��'�Uk@{�(��E�2e$)���	Q���r/ ���y�W�&����EIVR�����}���Ŀek_�~aΉh+늾i⬺�A����$irZ��u[���YS�DyV���}��eK�T����"�+�i=A�F�)�"�=y�QEu��h�����?Q��F��yl�"PqS��Y�-T����:n^t"����S��h2^3./$�r?��h��}�? ��T���q�q��+�e��Dn�%A�UG�vc0Z�	��a�Gy.��㿾  E�gPdU}��;O�x}��~��������ra�Ğ��J��6����&PQ'����7��c���iֶ6m+�X`4(�Wj���J��҈�%�X'ΣR����~kyr 8���p�N9�n���pˁJ�}���C�Z)��S�>+�;}�t�U/����j[{G�O��$
��N�"�~