��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e����d���f{��@����S��>���4{��ת�AO�Q{���X��F}|6�$�|��fH�}c#��'��8FY�U=<�+�y��)|b�x��}�f-]���f}����F��l�����������e��.C��GX��8��,7\($�[�R 46��X�Q��ó;�N����:��Ff�	'�ghތ��0�����Il&��f��/)/M��Nem��lqc�GC��*���`?7�uӓ{�N���{��1O������]Q���bZ��ܳCU�|pVX��!3�������h���[����GQxY��fC� I��h��j<��o�BKm��!�K~�֎r`Y��˿�Y��c�N��A
5���	��{Ȟj�P��ި��"�q|Y��=v� ����`/U���DC��ve�r�i��UgDc4��Fа���r�H�c�_$�p��uC��	3��K�����V��1~@Y��h��QQ�Aż�K�y�)W�Ϥ�p�K�vIvm�L�;��1Y'�朏���$�ʱM�NR����D�lR�o��!��}F>�P!������2��� �(B�k����8�_������Ȕ.B��ۻKξ9|���WF�~{��
�4�Ʃ�^i$89��f�a�(,�U������,�Kx�b
:���-R|B��v��T�S�<��d>OC��o.��7�(���Iܵ#�����N�S��)a�r�T_����B��@3x�f��2�=��m1`EaQ[��&�G[�s��#N���wc�-��@�����o�9���F��~ �7�u�^��7���0�m]���������!��C�ķ�{j�U���s �P�9�d�yU_:��޴��b'�S�fm�>��(I�fj[�V�:�� ��wي:�����عT�7DE�;-ٍ�q�^e�'�{}<���P��Y��s|���
K���H�)��}�г������wd6VG�c��YC�yjY�^K�O�
�07���Q�~^iF2�;��]*���V�-�k�߾��٣�N���D�|,XH&�}s8!����'K��k����Oᭀ�G�uJ�8���ܞnq���eGH.�KSwj~弿A5��H{
b�Y��/��K�6,N���+Lo*���!�.��46f@s�E�ol��b�R�H�˱ ��B��o��R)w�g��SYt]]{�k��*�ӧQ���Q�6/�^hG�:�(��v]����~Yw��NX/%��.����~���������~�X�'�4�	�ZKE�<�б�����H�Ǯ*xI�G��G>��̗z|��|�Sȍ�s��8bu\�f��>��Ҳeo�ۛ�f�c
9Y�J��R�A`F��
f~�(^.�zU9U(:>�܃����\2GA�?�j��'�s�NB��p�,�R��.�cr�������@�1 ]qN#D����-�iJ�z��CYd{�;�����lhY��>c*�e	�����o��q[�3.�"��օ2!l�Ɓ?�6 
�d��!�V��Μ?{�5PQV�ò��6���]��27ީ��8��c���'CF6��w ����]��qd{.K�l���fs��|�`�M�լ뀝YLǆ�0���u�Z�%�m�����C�n��pL8Wl���K7���YK$X�����������}%�e���)�2!��3�h������P%!<q���|�V�rs��
�:���>�p��+�%�X���	Gqa�?�#\�-c��(���[Z�r��%<	@�s]i<|Lf�����Ý
����Nt����1�Ǘ�9	,��,�l|���H21U�M���_�If�!�!��	�f�Q:�Ġ�%Y�VbY]V��bP	�oA��赂~��t��yế4��!̨H�Ӱ���K�k���_%�H��:abwYh�U�qvR�/*���g]?80w:�h(�p)�^�o�-�1u^>�͛�DTwҍ����Bi�f/�Y��=�kB9B���8&dH{�o93්�1D8����:ufA�'�&����]%|��s�H�`�4�_i�f0����Nf��vd8�3�|�-.�2`�����lX���o�j�=z+q�Dӈ�A ��5�,5JXQC���>W9fpU�����J����[19>Bʂ���V	���r���6�S{�K6{���Ʋz�@!��ԣkd��MZ�)M�.P{}�>dp��@��{#���|]��U@��+�������޺Ier+��[!,�WɺԘ.y��7C����k�㟧�W{���5)���POBN�yW��**u?�X#��mHXyC�υ,���E���8� ���p{��}�p��Ѱ�蔫�2�?2��*΅����1U`�G�����S�k@���l�LиCsz�L;.!�F�v�o3�nV�_��g@�Ш���;�uW+�6�7#]�!\����������M��H	w�S�N�nvo7� ��k3��%ߕ���i���r��p�3����/������٘���r��-�1O/�e���P��?o*���%uy��A�nG�`��.������ɲ�e�R�*^$~��������T��{M���jV�ێH+�A�x��P����N�jQٲ��(��T�����tX>�䅤�*zq&=_�>�1�2٦C<fs��%`�y�C<��VB��I'�k��p(�tf�f>_+�[�D[/�7�@�<3fG�L.���j�1L�����s��)&��QUP�{9h�T&Gn����:֤@��4e��� Z�֢�Zj3�61�8i}Xj���-j�_��u[��3`��^�es����{�"e���bQ�������� �g(�y#44.�S��'��r'G�~��ҕ!��`Y��E��5�,�B�m�4�[�b�KL����$�O%�p����_r�*�͍���X�d������B�jm���5Ľ�4TD��1~9'�3��_�/�q7�@7�L�Tp86mPy���.r@�����s�8��;Ӿ�6�)O�D:��_/R!�	!���jc�Y���WMS�S�	�9������-�T:x����4��-�Uf����r�����E��L��w��lM�~��f
��M!K�f5l���B��2��L�ZU�A�t�?o�]�,�%�r�����7�~{G�o��{�+�st~�1��ɽ|�T����J�R��M%���7���x3�~�zY�l���u�����{F���>����7���Lj�G
�.�S	�`�["�w��Nu���4�FG��4��"�'�!�4��/�s��ҋ�_!�@G:g�-�i��.�/^��u��j�\bp{�"����N?C>�"@��Ң�WUy���0�I?tjidW,�`�����Z�0�d��5�s�(���\�-l�L�qd��/a���b�+��&	��+�$���'��~0���� �`�#��
Oɾ-�+�����"Rlj��0s9�>�'��x4X�`�^����1�@R"G޷3D[N�˼��,��(0�[���|N�[�v�k�]�n����6�m�W�@�܇��hsÝ�b�?�YQ�a'��d�8?{�``�����!u���=�S�o{�E�p��U�'Մ���`��CU��z4���:����n���I�oY��-4���bjR�Ы��(�xT�^�24S�ؿ��?aI4�������-8�X}@�T�Ȭ�:\�[�X�%I�@t���ϣ���H�ǖ��Hg���k0N�!-8(���c�zH�7�k�A绲~�����Ih	��T^�b���V�j���Uɼ��1Q}���2��?Y;��xAϞu��צ{�gpPm�2�q�h׋��B��k���s6��/�(XL��^۪D_�Tx��<�Y�p������r#�JuK�l�D�s�+'�.�<Y��L&_I7�q��%���-L�~�V3����J{�!����c`MZ�עg�A�Ï\�yY���<��/{�&��vN9b4���b����T_�H�7�=�ú�:�V"!������"���\TC2Ф_���H�J[�԰' �x?�|�	Np,2կۻ�%�>\����!��͚MX��'H��,@�����j�Dl����,\������ ~�֝�����L��L����u�i��碤�m+��$:%c�ҹ�E3=��3��� <Tܣ��v�6͇�����0Yb��S����*��Iٴ3�O
�I�r���h�|�o�@Ne5|50���b\d�BX@pj_� �#z��fm-���(t��>�t(U�!>WW ��jڬ5r�C���1�b�f�j��jZp����� ��Ob�"$Sg�����f`xp�����ªj*J���Q���%oZV�����y��Cޥ�}����/�QWz�t�Za v��|��"�IY^��Ry�0��w��n���ё�t�p㮥�o|J�����k����/`�OAE���.ȭ�Lߙs�y]�C~p��W����k�eH|� ;�#�O;�l_p9Ɲ�Uk7�n��#�R1�������#�)؜���U1��[ػ�˽��G���mw>ƚ��Ғ쭍��Vue��p�'�����ʫ��pLMc�����{@�����b9#��\��0-�������R�x8�k����+���piYZ,a�xy�Ѻ�]H�#F�����lj�w�̱�7��0�*�:���� )���0�=<̞Օ��}�
�Zs�l�A��'F�����x�I%a�9��d�wB+�A��m��$���`?~��v�
�IkH;�A��l����I�z�H���|/���("~��e#�>�ct�#�÷	a3�mr1z<��&������Y���H�R��l�oo�!%-,�k��`�M�Q�O.q�N`B��'M2�z�)��!`���U�aN�(n�$�y���#`�]pD��b'S��k(��ou�������G"3�J0��m��a�` e.�9�G��(i��b?Tdq���Ns�h؉��Wc����[�U���KA�
�K��V�WϑL��Zc��(�H�M�@i�y�k��1�`�`K�J���5�;�,v�Xw�ΐ�ŒNL��o��9�<":a^%*�z�3r@�gl�$äb�$�����5�ъ���l�C�-W
��MB��$@<��]�Fnk.�t���=d�ǃ������Ѳ���@����������� ����M��֩i����&�W���cy� 1�<�P4װGb�q+�j������i��I���d,O�k���L�D����'����"�@��+[vF���N�)|d �-�6�m}a�o}�~hz��r�;B�&'�)ҿ���н�|����dϴ��c���J���[��\W��u'�d
�R;10���;0F\���Ո�]�`p��Ψ�/?��U�W�x��NAg���Q3@�q�ʂ��7w�ݸ���+���Χ,q�&�Z���Й�l�~���E���I�5O�T)^�)�X��c��	&��:y��Lm`1�!b#�x�hBw���(�#�%�<���_(n+&����u��=�Kq��]�a� V�j��\��h������b���Ĝ���D��T�����P��Ƙ�P<�������*{VHHR�Fw0ݩ)��$v�|�e(ƇZ3��dA�H�	Ȁz�]@��شRU��9��g�G,A(T�����{+�셊&�@�f;��uq(��e�P���+�rN�K+�=�>j��sO�~&��e+0�nΕ�B��3ρ1%* jrW�1>6WˢĢ�k���2�O�Se�?謌-k��M�\p��"Ԯv�h�@F��eh#��V^ �i���ȴ�Rx�L�VN�oX̾sHˈ��)�{N���{Ѭ�g�؇����v��8��3�M%��� �(���#V��1�3����yX�^��F��k��f��Y�IϾl���m�T9��_<��e����Iܔ#ނ(ѽ��J�F�@\�����l�9��/��GB�eT���f��<1����`��2<Wi��ZE��f�i�`�Ơ̊g�'(�~���QX����0��ܫ�c�`k_�'�<Ċ����M�T���$����M�t�gj+�l3t�]M>�#�qO��f�S��[�1o����4���h��l�[¾��o�+uq���xԙBÔ�U��h��]C�n~�#M�YϟCeGz�Oǁ�*�ήU�;����������8���8^5�7�&�rfvbr�ߝ�+뛼�E��t#�Z�x��ߏw�Q�~h�ri�K����;Jؤ��J����.t� ԧ�b��Y@�fTq,�r~���Kqd%�5�Lv�;.3g������ͫ_�s>���A�u���w�L;,�@<��,���?۞�@��Xi��W��C�)�#��	��"��\nO����pB\�ʏE��;�AD޲�_�Z��^<�.Z�Q4����9�ͅݞ���K��ʗ�r���$@Ӵ"?��0y��w�,�1:ww�rt
���aU�ԅs��t����x�\�cL�u?�IƎM��j��Vf������b���9S�T"y����Ϻnr���+q�W���݀��ms-3��(�(��9��>]�e]�*���2������?�/����L�c��};��y����web$5nID,f�s�&�w�����:[��bnĵ���w� `�A�v�=��2e�0)82��и�k�gKo{���m?��aC��q8&�'n!)�,	���y��W�=���d�Ҏɞv�hR;���XΖK�F1��@�a���g�V�;@=�
��a���)f����q��q<7G��)� m �n��Ic*��m�[�NH* �����U�sR�'Um�|,ŢA
�^�jK�"L�(�;�����'��.ђyH��l
&n}��5���\}��,���x�SЏ�-g���iA.]�fC�-�Ʋ%�A�ȡ�с�r԰��������x�})`���^��B����	�ȷi��3z;g�=x���
LDo����Jv�Wk��
����X�� gk~tx,Gi~t�������=���J�A�sxl���i\�g�o�*�
l	�o�s�n��5�����q�<�\68E�ر�����f��^QX?�FnU1�Ԡy[A0��<�����J���1�4�}e�<�J}_���,�['���R.|嫻��HC �0��i���0����w��f^��#!�Mm5hK��5Q��79e�u�ϳ�"8���a��^��eb���ɽtᎼu��a���֬���