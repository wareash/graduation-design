��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�k�۸�m�i(b[�{�㇌�]�i�5'�`;Etg
<������H�W޵α���N-�`��6����ݾ�FF��eF4��_}<�ےA�[,�|{�?r+-��]n?���A��#��Hb�а~�g����o�+5FL�cu�ȗ$��ƃdY=�7��1��2~��%K+U�rI��5��j�d/���ޗ`KZ8�M�07�H�4��n��@��n��P��u����������i�5��6���v$`֦�Q+b�g@�D�N�N]�܃��|Q�?�AW��	��b��.�Z*\���W��%8�yB5���xo���Q_���8���5jz���v�]���˩,	��T�.���B��N�l���%�OAh0��E;����08����}R_Y�����|?�I���rX5��1#�σQ�5w� CY�>����^zIbf6_�/�n�j�}^Wgf���jH�z�b��;�j����q�)�8�M���)��p���2���uA*#˾Zil���\���ȉ�eIzK�u��y*LmU�`��߭��A��\�%�Mˉ�(��N����A����%�����K����g�������..�o�D?t��Ͳ%L�ZP���ͬ�ȹ-mJ��}}7�t�����)E�s���o�����(�h�Íڳ�ݝ��P�`�>���T��ɮ�s�qT>$ΚY��N�˷�.)~y����4$S�Hi��,�Q�~|{���;��#[��6��a��w�H��nɮT_Œ�����0_�y�'ʊ�E�$jD��sT�rgx4v:�`k��<NͥΧb<��F�4��'�[Ωî��]���p�ֆT��9{~u�;�'��-A(��Ȇ8Vɮ�a�M
���Y 2K�{���w)T�^p:���DS�F���=�1�J�"�S�%`4ڙ~@��{�q���N.�ũmG#���q�;��u2�	<��f�E��i�?D�57C��uϫ��i���3&t/���^t\W-�{ ��S�#�+B"�諺��R@a�↻Gs�8��	�������I��&��,#� �)�&Q��$.GC����Z��5�wT;&�7�X����#��.]3C$ݣr��Ɉ7���]{*k�4�� ���C�O:�n���c�I�Lo�L޳]I�\X��x�F�CU��G�BH�����#��v(����u����'�Ļ��CGr
x�DG��Y�mJe3�?)�j-�K������Â� �Y��#�x��p�
�GJ��L�.��I�E�o^̃Fzޑ����g�3�/�t�FچL p�-�P��D'�鏇��V���:+&#+�����8��UVl}F2\�0Y�-��2��LdE��Ry$ �-"�_��i���	�ImA{C�F3L�4�`���<�2��@��#%k��̨���$�\͸`^��*���gMx>a䒍$M�2o��Eq+�@6�j���jk3H��9\�{��.4�ϫ�X�}������Y	2}���Z̀G0c� �\�WtR��E���h=r��l�&i�1�%��Bҕy��+��f���w�JJ.�>�c�n�=VR���@��.��=R� |����&��fI�}!���/Jt��;}�l�u.�m��~U+>���>����΅���
uJ�q1�]P$%��Ct`��%�v���h>��㽴�;n�҆�Y�T��^�����[��i�����G��������s�Y=pL._mS�G��5Ӆ�\5���
"�ʡ&�՛��x�/u@��38@}�
���{�>T�p�s���yN�TDR�V�=�\|'�i�o`։��u�V�Wy��X��W���N�Xs�I�
.7f�2�Jd	!,@���\ʨCt��@�M�>���L�N���=^��6��xAH�_#+{d{�;Rޛ��HꬷV�!v��{�����>�����XA%XO�E4��  ��d�� �%A�z7���]yO����jXd%���s�
��p�J	uL�޽(Y��
�AAPI�ևО��&��;&��mQE�B;�n����4M�f�,H��A)�dS���U�����&S7�F�A�6�����H9�8x�ly���Ku׬'�3����$:���CP�$l�䆿���g]6�)%K�%秡�������� �I=�a��I��;�A	5w���(��������ʔ:�s�2�8����e�� Z]��Sm��4\���i��hi(.�>��?�K [�g%�^es�6Sn�ۺ�!�M�Uu�ICZ ��F��1�f�MIƪ�*����xE�7x�����e}���.�	`�8�w9.ci��6"���Ȗyo�@	XXz�b'7a�	H�@<$]5�����)	P��;��	U�J3�����Vl����Ku�#mW@�Ty����|߉�C��$0N:t�K�|[�}��$w��|�����E�;m��ݸ��h"�1H�:+NÂ��F�y�ۿ��*U�qQʩ�|�3﯍.��-�}\aVN�8Ԙ"`�W�3��a�@l䟇����KN�r#}ܤ�X��`ζ,�J]��=�}W���<0�0/��R��j C�ٵ�o3B����� 8t��yk��e�����)�r~Z�P>���*��_+h�m��E�FC��Ɓ]�	(�O�TW��֞���ZT��I��ZsO��U�Vݯp[�x�q�>h�$����월
��qt~6%(rv�8)&�Z�n)ũ	,�.���U^����\�eB9��hxm���;�R�F {�@%_k�#c�=��̉�j���-d�^3�Q��fބ.<1�CD9j��`c%�w)�ʮ���Ŝ�s#�D�k{�����1e�#9<�w���,����v�r��B�'��U�u{W{��q���E�VA};P��x-�䕀x���o�a�W=�`O��dδ'E��f���\����;�)�]�`�~�[F/�#/�&�ibV)�.d�0���R�h��	�F���d��#]����,����.�C$S�8\ڔ4Qٹ��>U�I�|V�]_/ƄD�y�°�,
�x��7X�^� �T\��$�w,t�Y*y�ޟ�pyE>�R��'���q�r�E��]��PϞ��ѕ��3F+�3�$7�߆�&'h��b4t٘��b��}z���s��
�G�ڟ��������7���.�_RIc�
R{�i�5ZBZ���8��%x�e����[��2�>��ܕ��ӑ��T����A!� �9
x�FX�?S��ZaԦGKM0KI���Z���t��/�� �ZNW�V�y�lH�c�K����,&|���Z��Kޔ[�./Хbf}�&约���_�m[{/7ڍ�;m��N=#1?m)YB%��;c�sE
{�&v�٪t�pډ�>H���r;�D �̓OD�qW��>�;�%p�8�����y%"�ެ7�r�'���hQU� p���I@O ^��΃_������sHƮ]Z��q�lL�fc�@Zӽ1�R�5&+�ΚpA�]~�Թ��gd��|�g����[k/긴��ORv�\��ؼ@�crN)W鎚��\K#ƣeQ/�tu�,����Un��u]t��m����˴q�+��=��i����}�Was��uqAV$g��e�"n(�O�O�`��X�}o��p�6��d����2˫@V���N���1��{�Y���ꢶX�b�)�CQ�7|�k� 5��}�a�@D�s�����iߝ�[䑐��7HW	��-o	RюP\�#{�b���]�&MI@`��KU����A�pow�Gl���t�ܧG�Y��#P���� �2>f�@@ߵ�{;$'�=#ب�>�HJ�n�.���8�3	��
�lN�D���k]so���c|W!3�$s��2�+iҨS 	P�7����u�'03A��k\L����;W��q;Aj�Rp�RC7��: t��\��]�`+8:� �����*wF��|����4�"I�=���ݡ�Y��fz��:/�_�DD�F@���a6>��i�դC`hOܖ�S����VƔ�	�
�����T�]����i@��jNd
�s�g_���[O�M��A*�8���tH����}�D�ҋ��%:��9��e�0�`*�P���ؔP���zq�������pAtщ�9��]՗�yl��Od	c������G[�z��JՀ��~�_��o�B��`5�B�bC_��׼c&��zӷR!_ړ~��[}�=��"�����������c%"��J�ް�'�JO��,w�	m�)���G˘>Rͷ	��OE�]��&�7��%xW�Ŧ4�.�z08��o��O���Ҿk%Q�i01�q�;�!k�>�zwo/�mP���잾��G:����Sn��/�$�,�1�i�O9�v �\�6�b��5Q\�SS�ț|�䭸�J�X�O�9k^-|�����ʡ/��c|A�i����w�<�-��G����b�;�ˎU�!D<K��_B������c���<��ǟnWֺG�;�a�?{f<�i��p/��>�MUKܩ9�`'_�@�H'��D��h�|������Dw�1()��9�11��Fw�E����+k��Iqm|�nٌ��K�=3�.X��xC���%{��z��2ې"���}���_�Ko7�ؖ7�c'�WCݚ�f2�m��	 u��$e���^�!-(uM����X��&��<�.?5ƨgh��د�E捅<�a-����nB�^k�Oz��5/�4�bs�A���_y��0�Hs�$���f��`� ��=r��J1D4��#6He"BRUI-��TI=�hS��|��-z���) )?Hݽ/z5S��<