��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jåا{�\�u�?߷�dn@6�zf��r������;���:B�� �*�7�0�=�t�������޼_F��X�6߸�+��Ǟ.�u�b[dޖ l���\�.+��)��`���i��'�	�=��@�0Ƕ*C����2�/|��U�W��Z����>;;�������P�V4~I��Zj�9���4ư��3�o�
]�B|s�n�?�E���˛d�0�t՛�pz��̝U�ψ���uׅA��a�+�~ ����9��P��
=��O�$9�Ed&S�=9��|o���eu8�����(p�Y���dzJ8�2�䜛]�q&��{W�x<c�VN�;�$�x�HO ݝE�����MOHl�� �,b�4�g�m_x�*��ͼ�c��(q��i,�Q����242���O��R���Q�Ǝ��RpRQS�ah��Ukrl�Ң(ܳ_�F�B|yϳ���?��v��OWM���b�1��Nl�����a#Yt�O�U6��Woʉ�/~ŧg�a��w���H��6�X�e2;<�����	L�z i�/:�-��v���+.����b���R��^��̚�{YgV����	��0���'2���z�#��CM�Yw������ĵ�}O�(�nU]�,Z�3 �A�K���[qr�>
�����(a��'�T �$t��]����#������A�
�.^�?gns�r2N`�j7��sߓɖ�84s ��� �S����[��&�a�Oio��s΍�9��L�ۇ@�0��8T��&�z��uC�~#G�)1��5Q��a=�߲m�i��׌?"�W�ie{��]��ſ4��aբ���j�l��B�fEM{Rs���2r&�A���c�Py[cZ4�޸���Ĉ>*��扥�ٛ�YX������ϰ�#����@!F1�/��F{��\P�y%� �TVzN����{h9�(��,���+]ZGu~3&�m|ɟ�P�1=�lCw��3���h���]e`hs�N��t���?��e�U��$�=jE�3���`�qGw�A�Z�A%�c��0y�E�	����̀�X o�0�cq�_%�&���PV���"��
�_w���/,��Y��Xř.�lt��X*YY$d)e2Fpp�&%'u��7�B����+OI% ��,�]���lO����y'�_/����t>�m���ʣ��3�9�F�zo+2�����rԀhn��,&��#|l��*,�����ҙ_Û������R� ,$�� x7OWƎ")q�f(���~�«2���p���� !�$�(T�;{��V�x�8�!�GRfF�
:E�i�Ƚ�떻�̝**����m�Fg��|��g:����$Q�ӭ9�g�7h���X��=c��Qy��~}�ygJn�8�`TK�R���Df�h�Z� �?m�F��+�<}�#4�Y�bl�ԺŅ��Wa�Lz��nB ���w�]����$6�6qo��=V���M%9�}ˑ��Z���w��p��˄K<��L�-	^X`q�Y^r�X2N$)�h���2,�B�5��;�1�C��I\ x1��.�]'�uΣ̖MC��e2�E�l�B13����5���9�B�h�I�=hy�J�2�Xkd����vG�[�ĘnN���������h<e�:Lc��c���,D��-�hB��He�@ɌO�Bz�ɴ�>��H*�$�bx� X�6?�m���(�P*��ѳ|�]Tqe9;�]o�u���ԭA�v0�򿹢�*�X�@�'�6z�6HĊ�ڑ07~8R�	V!g�[��	4����ޜ�9�JUC2V1��M�i!i��{�!���h�+N�1�S2B����z�J~W�UVW=��x��< ���jv��?TI2�C ~�wV�2l�7(g�,jf���R/�
�y}��ڄ�D?�gz%��x�Jb���%�y��ي��9�a*n��v�2�ۿӪ=���{�`�_B�S����~z�i�"٤vk8�r�� 	�u�hъ�5�0/�׸��ؿ`n�9�����ӱ�W���6v��8�N@��JeNX���z�N���&��pF`��m�,���G�%^�.����GbJ̐�6Q��Q����(*V׶8-�L	�\��L�p�K��pd���ٓs�щ]���`Į�e?�Q'��V�fΏ�T�4�U���f����q�iD�<�	T�wQ&�iIibGw0�4$������ȭ�d��|8�fŭ�h�:�9�����3�!��BZ�ca����@v����.|�J��X��3���ZI������욆�!{ =��G�;�N:z�(h�=���
��XN��yS%�%6D�A�������O���m?���h���ŬC��c>T�вs�P����pק�8�V�,ū�$ƕB%p�߂��g���DZ����`�Fw��qm��
C��0 DKV�L��N3�Տ��I��4Dfv������/�Y�����\�`y WYg�Rr�����uf�$H�R���y<�]�X����$u �M������vBS!ò��q���B3�ُ�o�4h��-���g����(m=-8&����P����N6-����z&h/930)ֲú{��͔`���(d�e*���ϰ��ܫP�P�$��}�~�D�����_��&�vtU��K�&�2ˋ��|���Ub���c��l�Ý���.م��<��VKB�©>��>X�&a�y"�!T@X6�mCd��'o=$'��ͺ�"/1��s�)6�gI�?Up{��"`w�g����	Ϡ�� 
�LM�'�,�"o���nRF�^B��2�t_Y�] �H��_4^�gυ^�a�Q/��EM`�IO�V��څc�����L��ʕ���>���h�C&m�u��N��y�M�[�A��/Ӳ_��[p��-6),tS��Z͹W�3��$\���Pi7l�I�S~)�a�6s�[:��U�H�6uu(�F�Yo��1f�iN>Ck�P]Uŉ�x8<a��QKF�XH:�2<�������6]]T�$�+=R4Z��BZ���./��r6�Kv�&�0k�r<)�6$i�ݍVKQ/鶥8�{Cl͵����z{^�3LRA��4x�Z�z ��;	��po��5�'�Co���/ߋ�����D�M�
�jZ���,�͡N��v�Bӕo����l���ybp0�X����ъ��Jl|!`�Icv�K}���%?�Ì��4
��: "��O(V�@8֚�y:��� �[z�!4�H�x��+s�H��T+��|7Z�Ez��v]���c��%�]pV�\v̧{n0�M]e�^������ѯ��+N�J5��u���o�V����&3����jRfMI�ʑ�Z�e��R��dl�!z��1��%=�U3��ϑ���إ��/W��ia����
��-��v*��'��;J�������Du�r�)�e
P%{:4 �VsՖ�·�%�������h:�;�� ���zj�?�\sz%�)���#�G�%�LfͩҿG-f���>��j��C>������C��]B�Y���Ç�֩Ȁ��rB3iNހvd��p�/*d���;1%�#3r��'��TKP����c�Q��K$s�󜃆MǫTg:�ڋ�v;�4�9��2s����a~��MIYCw��_����̥.�P�JݲI��(��7�K�Y�U���R�F�D�#4h�BW�4�a�R���N>�����<Dla�b�wM�>��<-P<��OU�[E��I;C̨����硭�3P���:��/��'Z�.!��6F��o7�5'���l:+����t�鉢��/>W�:�D���)�k&���#W6��#�AX�#2���m����Wqp��u�gM8��h�9�(x�ţq���ͭ �4Q��s�fd�%��t�'zMoR7sK?[���I��?�!����Ȟ�Vٴ���dC�|��R����ܑ��=
�]O�
(Y����;2��1.�#
!9K�9�V�D	P4�=޹a�s�9�����l�{�..�\�;�s�Y'�U�~�����H��?]�tys�(ͼb	(�4��1�1u	��:�·��S6�6�O�>��S�gj哯a
�LDtT�Tk�oU��PHs�9m��N�k�n��S��/�ٶ~�ib�i���Fe�ej/m�x�X���h��n���DR�竒eNW7c/��c�%���h���n��Um�>A[6�0[�1J��Gg��Y+@��<��(5�H���� �)�d����$j���w>#Tx���Xa\*�>�<���jvT,uM�`���;b-�Vv
N�X-p��_�{��B�� }p�HNP?F��v	�^��r���#��?�co���"f�O���I�"��hU�1�6����KU� �Pxn��T���+<��w/ �-�h�ŁG��H�/lx|��?$�R^�����ǒ7|��+߉��2N7]����@�>g�\� ��k���X�by^��C����.E[��{��ȩ�*���Ľ�<�m�}�7qRY��c[37��F����4\�������n� ��<,�@5GA��q�0�i�#7���W3�J$�OJ��iB#+����KygC	R��}�њ��b�*�AZ�=�M,�ĩ�-tD���a�ֲܪ(����Lft .4��͑G�Q�	������ڂ�F�V��ڞܣ%ٞ�_��y�]���{����$
��eǣŅgD�J�Sg"<cXڨC��  дтJ�9���0��G��Ⱃ8MZ�J𰅏��˪RisnKh�<��[�$ʊeH�7X���A	��������>S���Cy]g�uUU��E>@�y�iS�8W p�����;�����m<���5}���܉ӽ�	j5����t !	�����ٟ���]ձ������yI*;fe4:�������HǩB4x(P}������1c!-l�7�`�7i7��bb��J�]UϘ\9�L�A�U�)~��%m�s&���#wv�m����Kv����OX��=�������2+�T~I~��
�w�?�':��7���.r��ů9���V��x#�hM5dD`(��-Fdu��CYfB��MTaM����������&E��+<��F)i��zo$Q`@���u���YV��qYM�ն&'��zi㤥s���ҍ�us���Ӎ`��~3^���X��۝���yI�h굒��s]1��eޑ���r.���4���l��o���I��$�U�Őf[�f`���O�D��&���� �S��2y�%�f�Hը��{���13�R�@��0����c�p���Og'�[%#�7��D^K�	x&r"��lS���D�َ]�����)��.�y�f�Z�ja� D?�!S�J�	bu櫭�XP"�\�>ǋk0��#��(��\VC��*�!�����W�0�fg��Pn�t��"�q6�K�0q���Z���}�Ժ��y�kz5����R��U�Ӳx|�qM�����w��ey;Y��}-��۴����k\�����Lmġ��C�����g�1 | )�<X8JOv~}俈�G.z0�i]r�Q�vȫ��yst��阾� ���g���!�U�oEe�9�{b��.���N�y�'��� �э�R\�.G\�n5 �R��8k%;Ո��|?̧��9�R4}���e���G��Wl;|W@U���=x�w�=x�=�Z�L&�~�-(.J�Z,bd��>mf�|g�c��qmM��4��AS ;��o��|A�ںEu��Fq������ط��ɔXf.ܛ�0�ئ^���\{>w��?��N,7����[�Ń��oͳ
��fЏ��O��J�iA���"/C�Q��=OcF��c_ng�Q��+&
��,Xe|%Z��� �3x�������I6����d�`�O����O���p�:��s����c�d~�Ӽ3��l�`Ĺ�qi���dC$�mv�;ٻdrDB�����.��d���n[D~m�bu��J�bo�n7z��tl��c1
|I�}��ۺi�&�z��@fԪ���1Z��O%rVE��#)�#����zE�W'}J�����=~�U[�0�U�j[C`HA���l�rxp=(ZYԳ����_��+O���GD2ў��2܌O��&P=�c@7 �S��<��6��)F�W���K�;��� ,�4��Q�6m��%B#�ѥZh٥ky���"�"h�E�/sO��j�w��Q=�s����6�~�Xfsz��U,nR�ڒ���U�f��wP���VS(���՟�u$��ܬ�&ltW'�dA���h>�`�\�HO�t �Xi?VTzd�w���sb�s{�����B��v���?�~�c԰���`�%�M���� �Q��qr���;3�76��a}�E�̉=.�Յsa�:�Zh J �YI�!n�?�%XU�W�D�!��L�Y���-TʊQpXZ�,�e5��i(w0s�páS�F��	p�.Y�B�xR����#�\���5�{��8���ҧ�b"�1��ʌÁEL���/�j�ϰ+���jC{j��;؏�Dnc��P�R��:��z�F#��:��h�_C*�@��r�vS���G��+�fG��T��Z�>ê��%-mh 6�^�����H��;Qȯ�x��_s�׫��2ciѪw�ϥZG��g�� ś96�bo�(��#����/}����w��:ǚ%��K���l!�04��w��bYa29�Tn)��@�v���S}�NO�O�"��Ԃ}�Ψ�i�;Z�;�l���|��R&k��'�s�g��-�$UC�i�Ԍ�eړB&�P��.8�_VC��1�c���?1Pw�*����{M��u�O������S�j���g�^����%G��dmCI/M����V�vogM��,Ir^�ڃڨ�ņ���B3m'ώ�����P��PC %<�(������y�4
�yp8x�]��ZQ��t
�	q,�d��kgOWk~�L����Kd'sV�:�)���m.������X�́�3��OXe�1.e���v����ٕ��ÿ�y����%�	���#�i@��@���w[G��'��d�R����\u��bx���-8�l�o�3W����v��{`��m���6�����]��PüM2}�;~���*�$���n���5�;[ŧ��K@C�����	z`�?���Εp�̭�6|�_�@
i��|�nT��پ�ȑ{)�J0(R���c=��c`R�2k�Qn���t q�o	r��Y�-p;��v˰�S�8qO���_�biϱf�x��-8t�=�%Yc6p��5���+�nN���EC	y����Ne�o���_,x-��Tv�ze�v^J�U+��5B����
b��áL/=�c�|$�P*�o,�������ٙ,���)�G����Ҡ�{0�z�g!�9���e��d���c����єXDM�k}��Q0�� a�g�l/V>�2��k�ZV��8(=�Ӥ(��M�}�D���} ���u��r����ݞx���&:2�=f����B�UH�"�7���hz����N�b`Т9Yq�>-ʮ�I�����1��ےO|��P�/��]iw�沫ڏF�E��'����@��`��~�\/�����=#�{�f"��(�Vv��.?-
�᳊�}B������%���9��9��3�)_�� �3���_�/��
O�Zf�_BlNx��O�y��'�$��5�qwp� �2t��8�s��jed���3�Noa�C^�,cP�}���Fg�H����3�}�kn���%%�(WT�ܾ{�O�?����"y���R��fƑ��P���֬u����,b(�Fuɝj ���q�QxO68	�׉&{kU�& ����T=(�_u96'b�[fDПl�{��1�.����&�q��� �G��,Nd�rS^��X��_�i�Lg,L��}�5y�h�4&vZz�Y�R�@�^�!���[��U�^A��p�ś�\���kʉ;V^<k��}��q�nO4�m�l��Bʰ�ֻv.��ˊ lbޑ���&*�n\%�����A��&�Rٰ�R���9,�X|��: s�C�b�2�-��ԅ�I3|h�8������b��IC�����n�-���3��r���V��5%���������Ґht ��.��B7p������C�Z�g`'�I?����FP7���~T�����3~w���W��8D��8Y/w,�;(��-S�|䳻�tV�b�;@^�`����K�����;WC%*��w$��*R��bCe�􁢠QH�N��l��B"�bԇ� q_�]�~� G�*!?���������4)���"��j�5�y���k��O_+�Ʃ�����������K..�c�;����=R����Щ��-��f�Z$�?��_�:L�  �&ς�!@�����7�S��iw�} ��x�z����G�[X=��jNz�c��ZcT�uw^'*f�ť_�J�Eu-a��,N�RQ���?jɊ��\�
�fw�ʻ�}J�;