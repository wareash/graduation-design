��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��/��Q�w���a5P��B�~�/�'̙���S{���^�qѝz��'�hřD~dVr�F�!5�=��[�\�bYzy��d�(5���*���D#����=�6�c�p�GCE�N��+�xh�Eaa�Ƭ�z�5>��>s(�oƤx]C��F�i�TϚo�2���E���W�۠N	Rw��#fa�E����ǁ'�iM�$r����?�W���aݒ�3��L��'�ފ�q��p��FU����vJ�k�~���l���wFpe [�29��Zq���)Rq�� �CPu�)�;��/�V�2��'cu�*�Q��펊(�Ľ��N��������PDEL��DK�/9pD�P!;��V�P?t�;�B�D(�E ����
	lH/i�M���rV�gzyK��N�	wX�k��2?Z]"�
����	Cd2��K�Ʋ�o�o_H���zm�����)�I��i��z�d`l�� $�r;.�6�o��M�S�>K?����W���X�؎�ID� �K�*�<b����/]�Y]Ka�����Kg��Bj寮b�:^��]sn��|7Wʙ$V�u�qb��[��%���RM��.�!j�Έ����v{@�Sa~� �=;�	CoX�'���h�x�f00��2�����ȧ3�|&�w/QSLC�l�J���mt��Y9��E�9�9�]%$@�}�vpw��[��!H��K������%o��L�p��_'W��'�����tB�����XĠr&��)���	��aF0��[p7(���Ēĺ�/a�9���SHܮQ!@���PW���THm&:�Ru�y$]� �n��<�A����/���o������{<fv�I�\;`��Cڴ;�@�s�#<B�3Q�K1�ݾhH��/�gx ��*���]-���y,M�N�1�bȟ^�oɭ=F��}GAs�	�~&�lre8��	s?kA�aZ��FaY�53o��
\.O3@B-��?�&D�jw`�)����'�g#6��}ae$�c�?��9��b	{AY-�8c�m��0�n�i�3�`x�_�/�j�h��ŕ~�%
2���	��l,Ak�R�Z��)���վK뻬8���Y���-@��@���!����u~�0I��?��C%�h
����"���k�6��k������0�E>b�|�o��M��O$���7OqK� f)i��2'=X�htOXe�glY��t���׶<��N��>`H5u*<�+ǵ.��,�1��� s�>m�L\�_���EJUi�{�gE�2���d�WQ�b.O�nZ)[#��5�O�h]�L����ԧ�8��2c.� �p�}�y�q|b����@���F=H�o�f9�<���� z��u��o1���)�LF�w�P��f�֦/F���q���M�� {:v��k��ˊ�2h�i��'�k�ٞ���J����Nt?�y��\?Ֆ�c�d=���ꊂsw[H;x��203NV�u���i�A�tP��wˢ$�[ѰV�(}N顫�=�Qanh�ܞ��7�E-L�i`������C�,ى����2 ��7�lav3o�;�_�����OL+M�B�~,�����R-\O�N>�|{�Ư�)b^�@0"#�̢;H%��'�PS�h]�+�cQ`�"h��L�x�X�C�L���e;Ssٓ�/�@P�ҩu���b㙪|����M����,aP^��ʬ%�W�N�����,�X�ӳ�1 _Z�F)��n
xYՃ���~���
iԃ�^�u�X<�l';��>hQ�𿆣ݜ��vb��/�"�1�T�Q�JC����%N
�����'�!��9�-=we�/Ri@�j�I9T-IIԇ��=�\Ǹ��T�q���o�rQi�jq"��|`�u$���)��ֲ��5�!�.��ye��pVx����Q��mU�{[:r�t5Ѥ������q�vQ�`F�*))���:
F�M&:�Qhi��ơ��,y���@�yA�\���%AƁ���W���P�sL���\�?X�l�@s>s�O��[��'D`�����p:�rNq�����Q��������P���^m���( ��Vx�l�1I�����g2@��E[#0�ޅ��4M�d����,o�Lr����T�J����� .�C�,��&�&?���l�4Ģ�C���>��*�	����3�V����I=n���.�ƧQ��I%�Fߒ�ȳ.%,ǁ�`&<	�r�Er�_A�X��К���̌���M��V��E������'B7yˡ�6�B:���!GQ���va���/Ǩ�������9�!Ug%�js�c��>��s|˪��k�p2;k�|��Y-2i���S���� "��a���8�|
�ǙiU�I�X~1~�=ڶ���i�����4��P(����Rig��P�����Ɯ,R��i����&�U9���wΝ�M,������4ḘV���;9��L)�E����$M�lg�n돓�:���so�O�7sr9/ ^l_t���p�����!U�\{s�Đ#��*�,��~;9f�I�U����4)@�L�g��FfMwh�#�ϭN!Q+6�
���/���4N��t�p�ƤP�so��=�������ƬǢ�/JQ�`��d�D�?�nTI�v��2�M}�����:�Ѿ���I2_k�W�=��4�w�*
L��cI�>{�+�j�rhV�;@��UYG��u��Z�mil�3�)h�w`e�}��
bWo�yu�hQ��
��^ɨ/�!��R�t��X�n�	� �Z�0�khBa�ϔE�Z/��D��;�����!�5t��PN1 �^��l=��P��h���l����4#��riJZ�`��91�b�����%�5 ��k�ؖ/|�A4"g#.��(ʰF�vj�F�dcy+~C���U��Ek�4LM�C=Dp��`hl��\�����T!�g�� d�f�T�,�v+�$L`]��/�|��+�`�ԯ@���0��p�w쓚X��S::��cJ�fg���{�Mb��m���lۅnH;z&Ɛc��[��	����Y���󬙷�/��X� =�VKGVr�@���@z��B��^!\��k��9��������f2U ��/�!���2j���ߜ���u]���~6�g�c���&���	sW�Zl�+xk�jv$ ���1q9���������q��#yS�nF'E��5
y�T������Øm)��=�ܴhȾW�Ҥ��q6�ա�ې�'�CTR�>�S����Mtq�mɞ4}��;����$܂oڡ~�F��	�;sk��'A	\{����3Y~H���2#Z�L��`�@�`̖���,��ci�21�]U�P��1	��W8mx�=Oэ�m��-7Z7Y�* r�F�{?��P��_r��aV.*,�y�?E?�<�8�̻4����l���7�dx���z�z����[��Q��b�@ ��!�V��k����]���.�a�ml��c/�Z6;z�Rd�J�o�?~���_��DD`r��+�!Q����U��Z���Nh�'�=��Oe<���"$��㷃۹�)(2�eԩ�5����t�=�/ �[�6��n{��#�~�)�+�	�/:��	�Xi�d��D�1 �_��S�4��#�U�+��@�������R�ب'&�����0�T���������_�z�e��2(��4a�$�U���ܢ�ٵI��D�X)r�P�nu�U�w[��m_lQ�.�2�[��Σ֒@j���v��׌#RV�I��g�c�v2�
]$ǹ]4'��׽O?_URy3)�����^��f~k-˫z�-B�������~��sS��1ٽ�$�f��BȂ��f�(�D�ST�:E��V�X��OF*�,����*�#Y�����z�u~%���u���*Q��L���d�p� e����Ğ�mW>߅r�v[5qi]|��ƋeOժ�݃,/��|a������'I7�0U�s�P�
}���b�/ H�A�'�h�[�8,<L�2~�N�/�+#���,ǸK������ ��e���򣋺��"A�sdY�3WʇTT~��(Ϯ)��#���/a���Q.]�T�'3����~g+�I���t�P��Mխ�B��i�v3F�˻K}5��
lg}�G�|�^�<-M(:}�Dv�F|
ç�W6lS-`k7��1�1��+4����GbL�w׌fr<��x�m��:c�tKN�T��*	��H=��q��5�u��_�ص����]P�l�a:����~a��x����,+� ���,RH~��_Dt�&"	P�&�bQ߸*��QuF�W�F�˽�^f&���n�熏-���1�z/p^�ɞW�s���>e��M4���9��1+���q�/�OQ�_�c�	0T��qtUʞ/���-\��hɜx��aF;vV��|7��K<\��:���ί:����)��e�I�o$NZ_`�8�0k��������@����Uj��<��k&�,�ۺ��; !�g� x�g��N*��NޟO��̘�0tW&��4Y?(@��(*g~�+��o�� ����H������q*;#�1h�ݺ��ķj�T���0j�,y\!��^q�Le"}~�Ӹ,�u���/TRģ� ��4w�?Lm_"//�P��R���.1��3��q�����V���~)1"O��FWb���6j���X��L��^)`LJ�6��V��(i�[�%��^-��c�y�͵8��Vn����ڶV|�'�p�4�&,8	�N��&�`絼Pu,�J�g���IN+p V����k����{�L�����P吾�K����T�>�ĥi|�t��dZ8�:8^s�,��S_w�g��D���嚾�B��4���,�M����X��'ɕ���i}�IO�
B�.5���Jw�ȯ�q���;>6x�>�R����V���Î:��O��b�K9L)��<���>�G�Ab1FZ��w�	��$ A%�xY����I,vrtX]�d<OY[Na<Hz��8K$�yy��kh���հ��&�rV�1�D�O�*�ky���E@#FL�\�)�>7����B#bIw���A�ܹie��d�	��:_�WY���N0)���- !}Z_ �q�:	y2��^[ײ�{~I�x cq���A9@6̋n�1w>Q�w��
���`��b�	ܕǬ��>0,���2��Y�/�?̬�iG9�`EV��1�l=�YO�'�6�-D-����B�MN��Y�!?=&+d�[/X���sv`���4��n2i��]g�{4���QH�U�����8ƭ�{��D�51n�x��ڇ���Ȑ���=��dU%�����X�;rR��x���r��<RG�S�����mD�K�R�D�u���0���و�fc�B1(��Ǳz&C��\Fr�sf�MW�c�#�}���X��Z�c`@6 �$��»���K�o�CR�M��w��]���a8�D����f�&�gZ���C�hl �Yw>�Pb'�5�+��Dڣ���1&b��~|�����!��V͛�a���Ĕ^`�����˭{�S�#�bN0s�fT��<�#X^LC�&W3�	���	��0���r��W6H���6#����]���Өmjٿe��3��c'�ar=bBg��� ��6�~7oT�,��˅n���G�<�
�w(���Q%��Ėu���aN/�iC��Nb���7#���./�`�y�s�U�<���m��f����Ϣb��zO�ݮ��i;EX�������e�p�8���n!�®/��$Χ���Te���%�q�y���c�~�&��S��@�G��
�X��<f�;�j�����S6��4jg�~�Xu�&?�Sx�iDkʑ�bX&>�9J�a�����`c�^�Q��Y����va}o��������Y �����4���b�nN��Ä��$��<nJ��YIX�^z��Sf�OP%O]r�V�E�,1�!���_��k��T9Aj��N���DN����ݦ�vx�'٭U}���.��c��6q�9�C���c7�3��뜓Ftٍ��_!�֎9�Lf�I2I��x��J�UVV����aF��jТ�:�Q�9(~��'��@�$ ���֚���Y`r&c�#�]� Wh�:���j�j��e i�ڇA�6nt6y��fM�+�А�-���A�������"&�`c3)/k��M������KN �v?֖3�O͘�%�����������PU6��>�j>�,���ԃ�ǆ����BC�u��]<܇d[
��&�O���*a�;}Z.�����WZ݉Ե�Ԧ#��w�D/�t}�l�A�l�$_�w��u0��Xꇸ]��
���YO�Qi�:a4�)��8��H{����Tgu�B��F)���/8��춁�x�͔�������Mkަ�05F	��F2v>�e���?-..��r���@�����"	q(30�g�Aw�?"�e��;�/������mC3��h�E��!���XD���L0�i��o� 0�͋O���������օ���:�V��������"x�]�aKT����Niӣ�Ex����_DN�Z+ ;�sTg�{��v�1,,��G�iM�<��[��B�զ_}��8~�']����^߁�)`?�R�����/�"J��d��a@c�/���&�vE���$�4�h�!?��ҒӴ��΄M
�+#�8��m�[&��m���f��**�����$� R�ߤcl�6�z����&��qFq����O������eH��yB�k���V8H���@�e���E��c�%��Z�).x�Fr���b�#L���f��	IJ^���q'�-��\�Ŭ��]6�w����m�����>M�b[FZiB�AX�BΏg]kQ;0!G�_[&:m7���a�o(ɻ�
s�%+�:c�	��|�"�zсE�`P�����I3>Kr4V�~�	O��2rE+\4�����:�;�*�$y4ġ��2�k���]���^h��|��Q��9�J7���bq���v$ZCPӗ�Ss�ƫ'��D��M��Q������Ͳm����I���)I���殱~WN"r
9��'����p��HxJ�.����0.m~H�>GiԾ:�������Cln�J�"�G8�l���V��Z�H�-�'�j��f>Q<��t��2��h��\2 ��B��$M
����C= �S�M}J�JKep�lң��Jx@�MF�W: �5k2�ґ�P3��:�֤����w�D'_5�`ױ��-ߵ���vI
p�KƢ�rn�M����R�������Қ("rD������:��@F�wuR/���u�}xH�5�ģ� �帍�N2M�6���ٺ��������1|�$|H3��4,/���j�Q]��'�Ҵ&3wٓv�4.*��v��^�а9<;��(��`6���t��R>�K�;{�ێ����Mz-��!�L�g�1��C ����5���5,�O�8E��ö�����S���3�%�eū�OBڷ��c4���\������4 ���[�z���]�2@l��E��.�����3T������Q��ZM�hE�)D
�.�h;`�Mw��F^7ыa��J��|��Ʒ<bşI�p5�V�ێy��
��ӟ��,�G�Zw���-� ��S�9�hٵ\����J�~z�:'ɤ���l�ᬢ�[��:�x5��r�G,
A������2
v������5M]��G�%,�׺[�g���ȗ�VT���q�ꍍ�y~ԩb�:��4�f��ݡ�	熜��6қ�`����F^ o�T_fel��^�4���eՔ�]ѵX!���oH��`coj{�YŧDN ��x�f<�
����(2��SS{��Z��4�0p���#ڧ$]?"k���QG���T�
��bi�o�:x�]:���� r��cp�1��R� ��H��kY�[�>A�X��A"�4����-���������E���3%�w��H9O �3��J	��C�g͚ԛq�/��Z&��0Ae
��� GW���7�E��|(T��������C��>��;��bv2��jSH�/�-W�\�Z��D�p삀�6�r s���\�����G�y����k�q�� ��)h����鳣Yؑ�C�/&����O�x
��N�w�%q���:�,�hg1"�������O5���d�駚�&�OI����a���C���{59e	��g?�X�K��vY���:��J����w/#�����q���(���������p#R�CG�d��x�&Q�ȞBPV���;u|���hhC�w�$�x<�l8�������;!0Nw9�N$��(�Z&S�0�LTs<Fo�P�H��%�χH��=������ټ%s�35��Q���E;l�^�=��4i]�<�Q�=�G�v����&�ۭ̿L�t�1�HgF��ʏ�'�2���-Mw�cB�I{������u��w��(�E��������B*Y��8�e7���q�z�"���t�4����X�
g���F�-H��amu�:�hU
�顚���2�L+ِ$p��>2'q�bU���������-*<��-Փ-�k���\��Ix�N�aݑ)�3=H3�{��~k���I���N������g����mb!���B�4�bS�"��2�8&��&������U�fLl!�/��_(�	��H��a٥_hA9_�xQ��c(Ҭ��4BY�u�����ܨ���id��K�^�i/$��d�
�<t_����rǫ�h�Z]�9$���%`gK�W��+n>!0���N@��bNg�*"��9��R7��7&�k������g��)C :S�󠡼TMy���w�Cm�#�=B�B�&��o��4p���f��6�>�Y���Z�'JHR�6dȕ��kB'���LZ6��t߻F��/�6�I1=������!���9����:�3R<p�&����J��r6��3�X���a8rj���YRD��v��z&U����iI�xa4h]45҅���䠍��Id��bC�H�˴�*&���ؔ_�,I�o��L����<iFx\�Ӟq@3?������)�����?~��>/-p��$����d�P6�Ԍ�V�IhI��!�ȟf���ָ����d����KY]6侍p�຀��՜�?�Z8bk��&Ie�vq�Ņ1�r�D����uD'�hQ۳S��1��.�� ���	���Q�	x^��ᶷ*��b+kY�i���޷�7�ԭF��T�7h�'��K���\k9�p�.��s-ظ}~�����찬�k��u�c��Ajt�箳����g<ͫE]����G��i�r�F��@W�GΥ��c��iH�i�i����K���Rzb��{t%x�ZQ�)��ٮ�d0ǐ/�r�|�l6+#�#-�
���\�++.�����Q9�KMe�Id��7�˦�����Nތ���S�Bq�d~9��s�R�-�����u�c4 �G���� E�Da2\�D��<�Iω�V���l�I��dk�Cĺ��_��6�-��cr�T�24�?�uS�X=\�&�y��Q�5+z���H����%B�v7����Jof���_T)�2�JX��4��eF�ğM
�!��5e���*K%4��o_�A����j�#�0�z�L�}�R�2���yF����'K�z��C�{��z$�O��g��ˮs��F�I�C���������B�����;�A$6�]�Nk��(Զ�b^��<ɶH$N��^�~�z����I\�r	@���=�	��x�������5�I�:��gIT����#V�1[�Rg/X�ͩ_3���m�g
�S��.^�훙���㙙(ә��1K<Ҿ���2l��8-��R5���i��Au?q�����߼���!Q�k���Z��u���ݓ�1�Ȅ���v,�W�4�Q�e�Ɉ͍ �q��6\'X����~Q�><�eHï���$LV"���gZ>y�ı�2|��rc��e �>I@����G);}�㤦�	a��%�M�=i���9�O�)�Sצ�?:�J��\%�<ѿ���0D��z�dj��d�g��M��W�B�?�X��	����D�t���Rj�봄얢�#��1�(`��q�pÝ{UDM���寓��<�?�/����o�g��ű��K7���G�]�BB�a�rI!�X-zt5R�,�&O�8r�U�|b"|���Q���e�B������e�}����۪�&��Gu����u·&�yE.�y�s�^~���d�_>��R����M��xxdN]v_�̞�cP���S*����Uh���A�:`��s��'������Z�#��n�k]����B�y LY,v�k6��O#s��ѕt�<�V-�$������v�Ó�ζ��ǎ����e�t���rO��E�|���;�i����{'Nn�\������u7�[Vg窶��{�&���kE/Q�02kL^5A�=��(��Q˿|���0������|���S�x���y�T1.NGG��ς���sj`�q�{%���P3�K*�1⺟-8~�����H6y��Ks��.��έs�[�e�Z/z���Pq����w�y�����{�j��׫y�Q��B��h��n��b�S�l[	�W��2O������k)lf}Ÿ��������f�o����of�^b
��o�D�C�O�0�\���W�H��˃��DT%;!��˵Ǚ^�e���������׊Cs���)�
��/�l�ĂM�[KvV��_r�h�6���C��ٕ�D~���*�_��	���'����@<:� �WOĿz�	k� n�)�+[ߣ(i �n�g3����͟S�B��&�b5p�\
��`W����;�bQ;��L�$�����crw����1�g��L;��m{�+��	=��__mq��q��ǳ�1���"��a+>��/^��5R��6;a�t�"X8L��i��aGn��4��uە.R�`D*����s� ��"�E���p�k�	f��U����SI�/��4�v�T�*w>yۃ�+:{l��͋�ߧ��^��Y�t�Ҟ&~+�J3���Ԓ��U%��/m�3@�>s�����|)���k�m��`�m������U�o���8�h��rϼf�V�u�bJV)�`��B˒�b��A�</��0�GM�SL�i���Ubi�gإ@�e�2e�am�;}P"�&>�~	�����G��I�8=��U�u&��n]�&���)S��c�!�10=_YI|B��>(4�I���j'���-�s�˵)��U��Yp�5��6�.�/v3Ʊ���05�8��2�v!�K�H!=������
E���M��ϾR]��L�������C 
��z�����M�<��,OeVR���7������x7���\�����z6��2����u�d8W�v&'�X��f�^��>�J9��_l�>�%ɯ���@������E�䴻��Q�����ӯ����(q	�C��Ӊ�<!�̅ۇ _�єx�|g�焬P��_�3���+�ݗ���gӱ]���ٰ��<�㶕(��WiŊ�=��&��ꤔ��f���12��!�~bY܉�3�­�2����@\>���x�v6c��
k��X~e�OT�ׄ+�2��V�H�b�Un ����D���p��L�^>�7�a*6Z�H3����"f�wT!���b����� /�[�#rh����;*``|F1/��
�Z��o;�b�qy�C#���5�6����,~O�>"^�AiDc�B��%�pB�-eI���W��A�Z{���| �3�Pl$���o��4�`����$'�A���-��gGQ`�=9��b������m�Y�����Frx1O	w'}��8�rP�������2&{)��JD���sp��W�gɭ}�n��#eQD�dF�l�vڄd�2�Hꞥ�\�X��a���G��$��N�H̠
$$ҿ�0���I��Zzb��sYطK>+�z!����a�[h�O�L��������[,E�U�\r2�G:����ͭ���V��L̬?-ZK{>Y8R\L��)�!"��4�������R�..'�0a��^[��ρ������C�m�X�	34<�e�}�݋�nސ=$S�5���D��s~5��� [AY��c*�	RF��GojKW	d�{�����F#�ŋjJ�f?�\N*��[;z �͕�R8n�/��ٲ���A��3v��@��^p�8X���y��_HM#[�{ �+wb�#�*X_���4����V��ߟ:G{�E��/Z=7�:�1A� �r��o܀V�`�VP}w�W�Y�� �p�DSz��d�@��>�v����&�
7°�C-��xq�ۤ��j���\�� ��-l�k�VR�oA�q�Ê��m0
6 ί͞���q�@�[Ø��b�U�=�ل3���ĺ;�w���n���@T�ܘr5�Y�
���k#zV�5-����{#M7�-J��@P{�$���,G��$���ɥ㬧U
X6� $KzV�(�n�L֖���!l��Q���'���G͘���Ef�n����f�.����5%c���td$�d����}>���n'Wpiv�*��C��:���3�2��U��ZcK�#�ު���W\m?Θ� B"��A������Tאj[S����3�qC�P���o��}@FOp�8FB�X�H�X��h6����䏐�4���>%;$A�H? �N:=XK��mV��1yv�e�Zع�ܻ�Z䋈[�R���(����`�ш�xD���08TF��mk�?��}=��"�5S4�̽vdD6p�N��[���nR�v��[I�\���O������
�[ӓ��@�+����N4��,dD?�t�Ob�a��tf���~2�I�Q���bqr� H�D)TuV[�V�ή<�&��I�F���ΰ�����63^R�lE�7~>�J�����@�"��<�f��Ln�i����ˡ�ź�YAɁC���JG����Aur}B�����r�F|��E*q��^Sx�;��S��%�s*��O��2�x.��jvYO�B
���A��u�O�G��گ�%�L�0j�$l�^�۪H�u�s��q�a��@4	C8�}�L��9´��3}�q`�	f��ShjI:���v��6���F:�W�i�B
57q��U�	*_�Sں��)5Ɵ;�;_XN(��|�QA�l��g��K�n���h
�?럶�  �
Z�K��˵���ux�d�1����(V�M���@R_�e��њ��B�������/l��P��_/��s�gy�*(��ӈ1��J��L���δ�!�x�V��Ὓ��T n@B��6��U|�a���w���+bY���_;g�fsԔp�.�Mݾ߫��៿&/�R�<o�iR��J�I碼R=�T�Q����4����-�9�,�F<s���"�2G��Xi	x��5��� _Odu�/�S�?ސ�h�1_t/2[|a�{����@ӛ֡�X�����
��B�Q	[P�լ]��j����I�`g�A��"6��!�8!�����*vj��3:�1x��/�_5�|��k�V��E�1�6�>n^'�N�>$h�;��ƍ���i��q�&;�f���̫���&�G�]��c��i��H%��s7%r��>�K��9���}�k׭+	�(a��4�ӵ����<�!`h5v=������)���Qb+���=�����+�s\D.@fI�Vzy�bG�H�����0y G��J���\zt;����F �2�]�Fr�[���:�Xb_��=���pIq*�i]�ڤ�J9��N6�Nf�����K�fh���Kk4�H�~C�˪����َ�/�Lz���)���J�W�h�������Ϙ/p�ѝ���7�eFR�E����v���1�0����������L�#�������ׁ(���X}/1�窤&����v���'�3���t[`g�ӗ�p6�yٵS��@�.�Jὣ�AƳ����$�G,xa랷��C&��?<u�;2M��	�dY|8�Qb���>޲�>�3��w]��bۈ^F�2N��HB��S
�u����T_}��+��_�N�a�
��{R�,jNe�H��[S�]8��S�)I�Ե���W��I	����<~��+�V�\���n~�U>�{1���ͩ���sq����u��݀�(��ް�O0�q��+[����9��e�Һ��cҋ�H�ܮ6�B�w�@�X��.r|�����}�=l��^��2q�����f�������=7�t��{�?�n㬖�V⽠d��������\i�g����}(@�31Sៜ���ۃ�TkE9��Lg�ȈZ����ۊ{JDa���`�j�_J]PHϙV;Dq
S0�I�B3l�${Ĉ���0`3h�"�����
�\CԈ�:�m?�����h�r�һqԋ^G�ir�&��ܛg��?�w�zNZ�x�+���Kՙ�=Ҷ�h�`.ir�OIt�5*!�d۸��F�|���v���}Z��"��J.�e�̾r�ܞI|Ɣ���Z@��iP��
�W�� � ��k<m��ZQ�\���4^��Rj%��H��c�k�~����'�Y���?I/u�L��vz&�T�L�᪟��f�(.�������U�N�O�]) #��}���H�ofֹj[�~���}e��2hE ��e�����h�)V��?�e���@�3 �y��|�b�A��\��0x�M�Wr_:ZER{�R��x�V�VM'����L���:����
2^:/�����V��o����T	r��$\(�����Ǒ�J����Ka�7�zE�����?�ms����L�H��}V�(Ѳ��IT{� ���F̪F�p�j�D�q�e�z;��^T]���l�ȑԞ9�X8�J-�@i@i�}5N�ߋ�ߋ8̙p�h���}�������5�3�B_vl<zT�l8?/���2�8p��/�15zqhjݎ�!P��noW���耭�g������,�s�~��|����h
>$���Orҙ�:&!R�3��P��g(�̓6ξwF��q7�
��W
�b��s��AK���HG�Uڲ��H8�Y|�um��^�]�W���x�S��lMu�>���I�J��y��\�FR��{�Ѥ +#kP�ۍ����l��5'��΂J6��:��1Ĩ�ؾm���Xb��V[՜Id��8:��P�<���k��(j�@���䵒qA�1�#��_Ѫ|��m�������efqC�D؈�^��q
g�=��d@@i�w^A�1c���1�+K�X�N@g����Vy�R�A+#�*|m�ܬ�& ���}n�X!^��W3�,L4�G��,0�K�OSc*�q����5] m9z�b���<�Q����ĂqÕr�,f~�.�hS��C�,z�؂5Z+#;(T�[	3')��y���F �,)��I���:��xD� ���K�_I��j�� ���z��z���=X����r|��q���K"j)��v)����$�� �>��H}���=�m~�]\�
rN��r��x�_�!��ͳ�OTx�"�W���l���H0i���������jޝ�J�v*D�4ٖ)�H�wB#�v���T�陇3��`5󯒓��2�O����� Ԣ�m��xn9͘�&��Y,]��-S*��q��!�	3���O���}������\r�u�NZҢj�����fr��$��C�]iMQ1�����m�9���{ٛh9P���r6�#�|m��N���^&�v�6#�ܖT������w/;A�U�{|��X9��x߫Q c%������ë/4�H4�x{eT�Gcf�����I�Lѡ�9�x�b��΂�:B���1�y@PV�љ{��,����r�O!Ju߶�'l�d(	$��~��Z]kӹ��;�G�@�`���^X�����O����ܥ[�q_wv1��J�8��Y�2z��c3Y��ǰ����AL�;k"�R�{������$V��7�pʺu�j�nSC�:���Ϊ��J��c��=�y��Y��7��	=�`�<�td�L�G�7p��O7�9�&���K�����ͫ{]���lD���.�-%�`��&���'>o���^�3KQ�˔B�T�4�д|��âB���}2�X�����('�΅+��Ԟ����̤0�i�`U8$05��+�*��w��Ͱ1Ԓ�[���]�r�Ye;U�A�k���
'��(��m�z� �n���u�$Y� �a^�_dyK���+�ׯ��l�6�4�2��X�%�����?;iH�빛�#�jC0ȣW.ă��3�(�U�K5��uo:ž}��C�MC�}�FP�ԋ8_�n�цT����*rç.�1n�u˭�t��p�2�W��N���[LN�e	�{ �b������|=߬��N�W]�BГ.�����=X
a9[�wW�V9�=��-P��
�쬝���b^��gz4��!h�.T{�P�MC��>��i���(Z��Cs6���g�6�pO0%���ZW��_��H�Y��@*�ob�S�^]Y�%SͯU�ݗB�*2VƮ��X����D��G���c���#���򫚳x�hk�OF��
�v)�Y�Ô�@=��M��<hɳ��%����m���B���z$�&����O��y��&��5�k�A�zq!�����OP�^x����T���*�I�'�,�I>�ek:	Z�(']��r��;���T�H�u�.ҭ�J�<
if�$�}x��\
��_5)d�YՉ��x��	�R+�*�)1��HH�E�}
�";Y�O����E[�3��ϧ]��C�G��"^04ϟ���� �4�>���O6�/�q�]�}����)D��x��ʡ�s#���C�K�S��t\E���4	�Ȉx�M�4��I�s��WM��Cj�ޭ5I�'�.^]*���Qį�X�0��-:6��&�+��C��w?(���Ē4T���3���;�e<.n�j�Ŀ���^o����1���Y����D����7�¢�pz#D������nљϊ�)�Q/,�^
�~�ݱ���J@O*[	��s?�l�I*�</=B�7��3�{a�"���8ږV�,�g���n�tC�Q��{��psM�YRî	�@��4�����can:$�n-�����Ûwq�纜5Ӻ,�D(�no���aaG�+(k}�_ڧ�If����Dv=�C}��H0V#�Ⓞ���
>UP���I��+o�@s�p$[��:x�U��U�C�u'@��^\s�E3-�\&��4���R�b����+�P�''�x��G��P*��6���9��2���������
�&W	�ƲdM8-�ͼZ�+�,
���m�q��0�H-�XI{g�5��9K�ʆ��dpX+��*��a�|Ԛt~P.���v�n�&#��g��)s�ǤdXh�,�ϡ@��Q��hk5�"8��>+o�U����#ݩ��t�Xº��8dG^��e�1}?q��+�"���=�[t҉�u�x��m���5r���4[[��/�h���32T��uإ-Fp���b�Q<}٤�<t�,-L�ʛ�$3�2�Aޱ�C,�6�ߕ��d�&�+D 5ޠ����H�j�l&�C�S��s��Y����2KG�.Q�Z���ځ�
���Qt�|�_��iQ.���6QdpcD|R�������E@i�y�T�_�E�CTP�h]:-��D�����\놵;������(���f<��'��!N�p��B���'Y��MO���"R������N��I�L�|W��N��G��7P�!��%!7�︹<��YrQ/�8��چ�+=���s=4* q�U���4�����؂K����R�w�]� ������M8����נ!�ԏ�:��P�_�z7��F�2���s�v5���&U<$-�ĺ�p��9f}��܍�T;�9�5�5H�mP��rԕʃу|_�������(fLN�����H�t�+��v���ˏ�:�`��iT���IO �T@V^P��h�7+>������X7A�[�Jp}����Pac��P�{�q��?b*J��d'��%S�5� �=Y�h".���Mu�����r0��+ֿ<߀��ۧ0dCCFj�� 2	ѼS^��b��ǌ��ɼ�r^������� ��~~.&�h�,Q�i9m?��Y�l㱬�1���m��96�2X�؏&����w�vo��o��Af�,�.�V%���2X ]�D���I旻P� �0���#�V/�a��M"��_�����&�~��x�T@�i�����<@���A)��h`�,�wI��+��w���8�@#���7� ��b���R�Ӗ����(d�t�t.=&p�2�H�}�T[���»�"W����S�!�}(\��ڝ�#)pm"c�P���S�Z�Xp2��^�^vk�K{VƲ��\��sw���w��,K�ϫ�l�ד_��X�"<pt��Ę���^�@�/�m;������E|q����~��G���M��;Ĥց�� �BJs�x#)���at�}��(0r�Ơ&����k�w�o�m&��l�P֡��S�Ls�����;�n�>�_i��|>>�b�3�O�R��v���/�ۄ�l�9����04قQ7*㞃Fڹ����yRgY��B�9���us�^����w��uw�G�	^��{j���%@��83f������k
���I�@��(-�J_��>[�����t��z�^W/��u4�v�j���ː���lq� X����ʒm��C�5Y�����#H������L�� �Y�;�9Q��~i�-�9�]���NVF�n��pZ�|gŝ;+�[ˌ�8���I���]���N�!D�>��4Ю��eWǤ.j�f���D��n&�Kpa���mݵi3)< #
�	:�ļ�AN�����S���zt�p�@��D���\ϋlO!yS���=z|������:�@,1:�T�m��:���*r�>2F��lLOJ 4���9�H�d�F�"�M���y�v��4�̑&�'x�3���g;��_xΑ|D��τ�M�u�Iّ�񳐶-D��S�*f<7ںe��6W@�%m[[�+��NT�ֹV�je�X���'��fo�����r�E�������UƇ߳��Q�t`|S���7d��@:?��6��yN���b���&��(-#QȡgIo�+��w���r�|Y4��uK�R��.		�(��.�%|"3����a��!7�`����As��RbD����q
Fx��Q?�B3m�g�Uј�� ߈���T��F�����,���C5g6��grv�5��@9�_��ӣ,��0�k�}C���2i o�m� ���h����-�YLbJ9�nR�����Pp_�?)�A��;"W�V�yP�]f��ͅ+ 
8h������m�����������	W T��7�"�k�ض�E����M�0 ŝ[�|��W$b���*�[��q�Sks�>N�5	�xR|S"f~�#l��8JD.w��KG�^O�/D $Jz@�m���f�.1���_�F�bW�<!O�\!���)�׃���ޒ<�B�g[��2�'F�����NLP�~F=!������R�[t��H4q���8�ư�,��%�3�k�9Y��C(�)�+�g4.��� g��xy�.�F������:'�ߝ�������������d	!���a��_ �!�&g��vH("�znhǕ���(��p��G1*nÔw�׎	�V��� ����L'�%E�j�"�������Xa<qa2��#���l��./s$��HҠK�I��fĀ"8r[F%�0�������*����{V4�����a�\"�p�0�i��hW��Py|0_�!���=�;-)%�T�z��̔;�;��a�w�r�3���6U��,xDM��ë3�}�gDG��g6������U�o餁3���j� 6SRڣT|���`?B�Q�Գ��߭'�6{��_-������=a���Ȫ�SK��E:���%��C��^Yο�!g$���F���7�H��o=�w�K�0��oK%��D���d���3&<:B���F�۳z�3f�?�u�{H��x\�/e�k����3JN� ��Q ?W���E�8����f!��-V�DbTMpiCL���D�
��tABy_�nB���=�N�'@�";��o�L��nJ�Dj�^҄`�r@F�� �B#�=b�f�J	����*Ue�1/�e�c��sx�L���H�{�D�Ց�Z�M΅�8; ��{��e�zJf1�@ʒ��[b�Ћ3DJ������1޺cp\���m�vHl|	�u�L�1`իL0�&j#��L��n���[�y�s��1���5��Rg�E/ᰲ�Jo��hُ��I(�6khO��焴8�˩dI�vR->y����+��q`�[K2��g$���Բ���e{�o����>���G.FY�z8��3���Ҿ��}'���j�fQ���o��F��e}����A7F��|>��Ѭr:-<.P���WJ���{CU~}u��\�ڭ�2$��z�,9E�BR���5�x�#��V���}��7'���Dnϔk�ow^������"p��+���-�C	ޚo��9bP�M������֗��wJ�hNR���W�[B���)t}lW�j�A���ي	ߕ=d�������ؿ)&
�� ���/���(E���bvI܆���T&c��C�g��n���~O�F$亿�G~�C��C�Zg�"�A6�<�㟪u5ޡ}�-��Wڿ�bgL�CDy�6_e�S���E*�L�Y��k�o�߅�/�<CfHT�j`�/��M����թ��:/��
�޼%d�g�`�JY�Z�`5������x7�͗��:q�A)�Y�\�P�Of��R�? 18�}�-���������6Tr��:��9�s;���D
4DV(eW��v��;�k8��㗞��PJ�pz��Tr�n��n���t��l0m�\�헗��v��0�	���྇���o�Gsᮕ�
���9�G.����V"�Y&J��~?᤿��Y�=��]e�T`6���l���]
�bu7r�/���R���|s+����wQT@�0�0t_+ԝ�RyF�E��I�[���,a��<i��Q�a��xz{��h}�h��my��e�j.2}je�艃���̑�$��:�����UwFJBi��EG�ꐆ�ͺ@��Q�.�-��wЬ��ݾ|�N�nj�<+����ErwU�e�R��5Jx��K���O-ݯ��I�ք�5U��Xj���`q=�d���6�@p'��pa"t2J�%؟!����J�H@�F\�\����G��L�ڴ0����GՁ�K_���24L���td|�fv�a��M`������J<@4����W�?�l�[��D^f���D*ǑՄ��̶~i�o�q��.�-��秛r	R�3�Ũ���;dq���}na6��u�\D@km)���V[��u������S9��M,q��pŸ@������ӛ4�}$�~U��>���R��yP��%5ϻ�'L����<rћ1,��C{"p��ukhb�v���g+���(��K<T��F�}Ǻ������c���#:S]qp�k�����>��y�|�+�*~7�*�O�mҁ/���}5�NP|�)$��5�����q>�3vŠ��k���p��@���-�!6>�K�~�@?^��4Cˎb ��b#�ׄ�����`%�aMa��� �j��;r،�j]��oQP��!�~Ő5��n�F.��� д�b �;���Ӵ��1.CO��V���>�;�3��{�ꯩ*��M|��s���2�2�兀��$(�˟���fK0N���Z��9�U�k7��~���RIk٥�K�`Ou<� ��54��d5�?Y{�)�����~�3m�U��=�w��I�"��<f��XC���<ϥw�H�����������fJ�g�Ҿ�µ!]�Ε�]���z���5xz�w�Q	}#ǮG�����\�%�?���u�'�y�I�������}`�o����[p�W:VuËd����G4ӗ�,������Ako��t���Bs�<��L�"1�ч��Y1�`P�	ԫ/���Fy��FB�!��b�̟��񚚧v��oJP�l��Ÿ�/�wR ��{dZ����x (����O�p��X��{f�L釥2�k%`~Խ���V��!\ޛ��\e��q����o��V)su��.��ZQ&݋9	�JG��X\��-�����[��\�]�y?8
�(W8v�T]L���m�{z�vl�]��ƾ<�. r����9�t2��yF�*��xM���cs�j�(DUK���B���:�s��|_H=��N�$������|N����O�F�`!������'���gj��7��텰.()�I�®_���K^�:)�ѕ�ʸɬ��٤��N灡Plih�xWg�[Q��:��p7���cy�d7d��;2�s7��åRTk���埸^WIA�v�[̬��!oS�ȯ���!X9�$�Za�p��u�N�nU���e�k	hd�=k�X,V���%�=}�7(�����`p�e��'�O�	Ix�$rX�u�i%��.H)���T���� �5,��>^S��Oa�� �$��KKc�[�W@��*�jM�wŗ� ��4�%ϔg����ayԢC�'�(-xS�F0mw�.�|����f���^�Ʃ"�V��?4mn��0�+Y�#����zͻ��!��\#Q �RbL���>��eܝiS��$ܩ��E�V9�c�{5�pi	6�!E�2�V�o�ec
Y0��;$���~)���s���8�QM�$����)�=ά���v��j�$�+g�/��
z&(�]��<��F[�Y�]�x?���HF�0�,���3_����v�Aw���çH:��-�9�o��gJ���3�q�ÂmĐE����T�Dݸ!P<%�dm{�k�<�e����q<��}Q���H
~)��0U�bi�e���̩�%4<��oٙ�ܺ��SӒ��,~j� �	�P�=J��`��Y�He,w�j��y��#r���mC����d�q�e�y��j��I�@��G~�����G���"䩵=�z@�H��C������a�h����N7�$�+v	�Jr=������S�n
�->��'[z.+�zw2�+�ʁ��n/�֌gqZ�бqn��
�\�p�.�0��P���E4�?#!��2�_�
s����!���PӍa��(�Ⲟ;�Z��G1�qD��n��c�ۢ%�M�b��`�Ty��"%�q�	:���J�����fWG �cgM��Z7�y����9�"[3ެ�=���[����yBE	跰W�],�&�@��(��-}ki����Q��`���X�@HP�M� m�w��l�.W��CE*�	��ē%�ds���!�/����5u����'r" �gM$�kD���b�L�Z�dw�8�q�E��	�z�_���4G���K�E}���3O���2�V���t7�a�ģbG��!���@V�D�ѓ����z��,����L��7�|di�j@G)���9t�,[���< 5ʔ������;��*���
?+0Y���$Vj\~IM�}��W!�A<���b���õ��o9�h��b�2E�+���×�Φ�{��vʪ�G��n�1�� 0�pg{�*���[��=��K���b��`�-�<�"�+���|����4a��h����3_�2Ͱ�%���LkyX8�i����-�$tebڳ3	�o��u�\k�Hr`�;�Z���7��4Kc���quĶ�4O�]��a�|P�96��s]�g�b<ċ����M"_~T~xwRV��-<��k�<	���B�|�w����"�����扆ew����dyXzϝ�%�q�aa覿D+@	#w����e�ҿEZ�y�i1�@��2���4U�z礦厼��L������]��Փ3�m�� p��[������k-��{�9\��~>n'c���k䑖�����Ի��C�rz&���&r_�(7��u�}wd.9gصe�w�P�Xگ.iɯ2��� ���
Pt��񝚔�b�2a�P�U�'����ْxj�$�=Sk5�Ϫ=e߬��MrQ5��nٗw�s�GFD@-��8�°�$eR��1�em�>��E`Ϫ7|ӑ��{���T�EeWo���L�2�uC��в�p`%��.�	�^����Ү ɤB��4���u�3)M�ÿy|��H(�jf��-��-L�gX*�ҜY�+@�1�F��Ƙ��nrEكO�B~���՟??�"�ѝ��ptb������B~ ��?�J�Amoj���w�����m|��͓��ш��̰@�-jW�q��7"���NG�ZM��5�nҗ]х�~��� ���PM��qo�W�~�����N^�<����Tv��i��w��,����Y:���=N~}#K�U�ap�_��)�>ڗ����~3��]9] ?���HJ�k�V�k��}�-�0�ބ�5���ONRQJu�+Ԩk P���N
�La��#�����?�8h9!�����f���?;�&��8���'�����s(�z\B��g��!�^sɾ���=�pR���7��~,�74i((�G3�q$�a0|�ǏiXC�	'��nt������^!N��b�⩎�7��L���^�A��[9��{SN^�%05\E�b�̮��cF�<��9�M�Օ�}��hS�Y���i�����k��C���z�/g�����)'��C���W��4��������P
jrz�Gu��aC`e
�V�{S1-�L�S(�3�2lcL�W�9�ЬIK��N���?��l���_�N:ND���NER�|�����1�*���i�6��fo���r�x�?xH��G�����R��F�����["+Q�E�曇�%\��4��2Zl�o�����Kd[�ʇ}�G�ԟ�))�*j:�t	�-0�a��)��赌�w?�!��!G!��X��DU}��n���miG'/������7�D�؆r�)xi��bx���2['	��v�?�ȓg��ۜ��U��)V;U�>��јԄW��t(t�<��v�`���0�O�����ʖI\S,;���.r"��V�\�f���;D��is�}Ue�2�q�vZ��g��*�kK�eT�.�8���Ie ��8r!0oI���%&,�H����l��F�t�K���1��Io���xӡ�`�|*m1��K��ȳ�"��a��=�(ٷFץ ʈ������p؆��-��fԅi
j��c�@	<h�ӑ�� �N����/ˮ�3Ɩ�B��dy+���&(K�~�@u�Y����=�vXo�U�Ɲ�  -�-��ўn����GD��Lۿ泸�_�-�	@6f�h)�+#Ҕ�U���]z�Ƈ���XA�e�,@���kWg`����Ӗ���j�QͶG���d]ϻ(�<���s4-�,5 �mxZ8.N�~�bX�=O�.R���F=���m�IE�*����`r%�B}�l��]������_���l��J5͎�����R�7L���Jz>�(I�$KG���Sp�Ϛ��Lk����[d��LP��u�����8N�%fU����W�b%�=������F,&�9��eMqm��.$�����yX����9�w�~�����^iھ�t_���k�T�G�O"�h�
���6��]w4�l��4�B�r��0T�ӟ��BN�d=�X�2�kS"�b�PV��bk�ƭJH��ْ~�H#���Q�W�[�s��h~�`����g��r�w�w ��U� x�ԺQ��f�L�'5y6���H�!%�.Q*@�|�3����_�Y'`Χ����ˈ�9пdt\������A��^f�_vG��J��s�Cunj0e,+]ɇ&�I�Ɇajpi��L`qs�dJ� T��Q������[&�ܒ� e�����fm5lP����DO�x�flɞ6V� \���B�T�̝�P�r;>����V�	��I���Qç(w�lb�$v3
آ�Mt�յ\�V�B�j�dI9}\��.���':�`K� �K�y[m�ܬ۲C��VBoZ�1��!<��.��_�޹+�*
������W*c���'ne7F��
ۮĢ?����bASn����y��@§U9�>��7��]�!y$䴺�7�s���;JX�b|����2���������V9K���j�ݥl*�	f����w����%�y�-���l�=1J��.���7?�"%�ؤ\���\9V����ke)���*����d|�R��¹��GMC
�h0�� ��_h��Ϻ�P�X�b3�^O��C&P�c]�!C�$Z"�.R2v@ú��E:qxF���P7��3�YԚv�ܜc~� "��OmZ8��l�|�w��_5��{��G9K����S�=�ںk"����_p޲_@'/gWhv�'��Z�W��WF��2t,Q���D�*���$;�"���;�<q(�Eh2j�j�-/��Pa[�h�~�U����;�\%�B�8�Z�qЧ��6���KvߊE��X����8�4e�vbM�,ETr��:�j���ˉ��5;Ow����Mu@`p}_�M �0Ն�"Ԇ����hxZ��;�Z�M�X����b������E��ϳ;ϖG9
  �G������U+&�P�ӳ�1��QEK9��t80�h�,2����s�a�B�x|,
��Qet��.�P�*E${�k��J9�r��9��Г��}�S#+���(��B�zM��3���F5��y�t^`�\ �����6�1�s�-��B$�2��� >��Q��*����05�����W�����������W���J��~��T9���L�Vi	}]��~�
q�Aw�6��ҋ���q<U�s@q������p��L*�8�)	?:>\:�#������{�1E��s�j�~AbL�D�QK�1(����3|��;�,���H��������5D��Qx�l3ny������ݜBK6�*.Xvމ���b�d�o�9�V�_
��I*��2�	���Ɣ/�&��+^S����^���@ڤ��x�!�Ц&��ˆ��	p�Fd�aa��yB��^�qkm��lC%5(Ӏ��X?8�I8�q�җ�*���Q� j��g��`�bJo�%
����ɬ�u�����a�ye#��M�����sL������}f���[��W����g:��4���M1�S۝����E��Ɍ���b��R����}X�#��͐{?�H���#�v��a<��A�&t*U��X��-0H��XiI!ߌ� ����fͰ���l�3ΤB�;���~w�{�>1��P��"�̔��S�F��c/�c�N��Sv���^d�{��L���'�Oc%֯��^Nk����^�1{�vFH��v�q��&�[0$�Ǜ�;��5�"�(̑���O��,�)�m5A��=�Dj(�a����t�_��:����T�j�Y�d�\-.�{(�����<��F�~J#��{x�|����?��zm����}��c�kV�I�L#pjC�U�^�8�SޒNIW$�܅�����L�U����%����1��IZ|!�]8�S���\���2��D�<ɩ�.�pj	����)�r�-�w1�Y�������>��|���:�5J�?Ѱ�I{yҽ�����j�!]�9J����,��8[��WŴ���Ff��*l�跪��f������T�E�W��7N�UBQ��w��MW��d���?����'[}���Τe�
y�A@u����{ܠd:L�F����⋚��rT��\!�z���%�jJ�F[�S�w����ř-8m�k/�	)�!^�Zʼ� `�rԟ��BI����l���e�E�Mg�bj~�Q$4��n�Ժ�}r��uF�?M���+���]N�D�*<�A��%i�{�k䡮��k�Z�.�v�H�@���[�6�n�-���ڊE֜AB�ZUnB*VՍ�����+zli҅(d����<�W�)L�E� �zh��|�(�Ȟ�l��f���Ɓ#���&/0		����+�'�fbN#KѦ�ĝ��{Hf.Q���W�^�T`A2��R�Y�)�&����F,�/Зޯ��5g�]�d�7̗h�-`�T8g��9����?�L�yz���직���$Ȉ�10��(TR� ���M����� �~Gͩ&�A7�.�8ֽ�Cc���e�mUl'�])̝�y���-��Rj�Aޞ���>'��-meaOd���?b�b9k�J���./�}����|�s�l��ve��m���b�ծ�gD���Ўߋ2|*6UW\��<׭Fy�.S�8�6�5�����|`7��)��B-���u9�i�3D�M�(,M:�pil�-HuΖ���3FN��ݽC�dّ����
�1<��ZZ��,g�e��=���;WZc��+���E��o��䷫:�ʑ�j`����P�_�q>�ގ�#O���s�gf�)7hd��/X4�S��f����&�̕��>�
>����15QZu㙅�Y�MNXV�j�*�����+��e�͟K�TI�u�� \�<�2�s����ώt�uI����k�7�v�,�H8�DG�h�&N$>]5���w�9otD��r���p^��;AϮ�hNҷ��r�p�?�	O����!�1<��a�L�g���  �¿�'q�*�=ǳM�M�"��.�$���νH����P���8a@��/q��Onqc�?� ��DE%c�8"����ݜ(���	�Vڋ�������F}����I�ۢ`*��-�dp,�F3p�{��(9������27��+c���F4Vh�5Ͱ]�Dj+��k�TG_b�ga(i�����z�݌���7!2�'
����<�0�����
�O:�F�;��||���и�#�G�sd��5�g~P�������b� V��t4˒�B§4%���<_:%;k����{|�z���y�u���`�ܲ�������8@�*R�����g* ���}\��N�Ф�=�ޗ�N����9N_,�f��6ڙ�ܵ�Y�ˬ�/J��
�j��م)��ڎE�*�: �'TAk���z7Ѭr�9�`��Qʇ����n���#L�R�T����ka�}y,+苫�(<�2ݣ���X��խik�z�40a�:>�R�ۺ�N�-x<�������@�z�{f.�L��i��1���ƱMhQA�Ѫp�v���]�ܯ��!�Xף},������5�����5Z܆��Y��H�T�a��|��s&h��j�~^���ל��Y�z�$ �a5YP<tR�X-j#h��'ŋ�W�\L9\7��C1��vL1���.�x�CŤ�PĞm�	�UX�d�dڔn��N��5������k�CԶ�O#�jϑ���3��t	R3?xfW'm��e�wi�byM� I�O�5)v۝E��y�`�*��EߠN���8ݸ�D��/Wq8I�KYJ��Y��Rė�}:4g�r�q��[����k=��)	�:�����=�+�5�j��"'?3��Q�˟$p_���ag�o�r{��+����0�L�C�N��#\�)a�d��� 6�i��ShHE���VU*ʈ�TĠ4L�����"�$�-8��Z����0���;�-!�ɱ�B�����X
�@�жdn��×����]�+z���^.Xp]�����$��Pc'�dX����7�qx��1C)��ô_#��&�s�Xd�d<��,BtUS�G���&ϫw˜1�L}��mc�kW��_~Af�T��d��آ�7h���������y�n�5|>��t�'g��t-��S���b5����29��8J��Ʉ=�ʪ��2�]��f_�=8%X�<��"�V���L�Wb����C��v�e� ���-j�?q���v���H��SJ��eh����>��������C|��4����f	�(aT��Y޷@_��N�׾��K���kFM�^�1e[�h<�۫��՘��U��9{N�0���\��@-&��ս���2�Vx;���k��ҹ2քn�F(�����n#�Y�r� ����4�:i�>K�囍gl���4���x�}y'��B�����N� �Cq�`�܆O�M�_�x�kA.�=�5��Z�-�/�&tQ��
����a����?@�o�(��A�N����S+�#T�h����17�*�3��K٣����ԩ:4�8�T8ݜ��h�2��|_E1�R7�[�+e����}���S�2���н���QÌ��ݲ��#���p�q��@��� Sc�o�׻�K�R���m���p�#?+%]�H�,>h����z��Qٻ�(���m�з�������W�
�k�
M�&K�h(ռ���k+��-\��L�L���ǲ�(�L�,g���&��owO�2�yI�Ǌ����8Uۙ��h��ME7�W��y'9�+	�H��Ro��7ht 3>�������-�eLw�Dho<����}��$��ܾU�(+������"����}p�h4B�Y4hA��D�?��@"Z�S,?-z���mC����� oG '�����nU�bX�l��X�5��k�jNБ�ۻY�c��n����]Ð�����T��e �R��fg�M(����-�j=u��u=�G��ܦ.t��`&!�*�\�x��u�[m[]$��k�t(=��͍�ޖ�m��g�����q`�%̆<V�7��&h��p�@0�1���TCh�l? z;�(V�Ԋ��TX��B��<*�IT=&�O�p��ߐb�*�&s��ڣ��M�C��v$�d�EMI�4Ӏ=xJ�r�MDt����ns�+U���r�0!J,^ �X=ͺ-�i�z(Ye��[��X�ؼ�2u!���hl�鼙��B'ھD"֚��E�=�ܳ.�W�@�l��Gp�UX�����0H���\<jfa�o�*]N��;_�G�¨ ���	��)� �;�����Ä�-,�׊*���G��/��ڎ���	1��1*V��Ѝ�Lc� ��M�G˰#��E��(gW�	�`x��+��/��}��~.�ɲ�LN'O1��T�h�=6W�K�K���.!����QLN���8^~���O�U��d�pIe������J����ɞ�k�b��8`�����VK��y
7�����,la&��8�{���#	����$a�Y����#�<�[����*�w��q���`�:c��]�����	o�*D��%�>
��� ��(�;7�@�Qq~����0
�7v��@��O$���i����P�y�p\��ީ�5��s�i����C\�ى~������[Na��yWb�^���Ts��R\��An6.�e��T��C��9JQ�����G{��b=�Z㆓�vq"��a$xe"Y($l�ս:���j��0\x9�}�q�Z�yㅝ�	�4X߮��O��Z��ϵ�p�����ꮮ�a�� &�${���k��⟺�eӶޤ��
��X�.������2�%�c�� �2�W��bK�۲끍�pc�����uV�/.t�3˾$o�����X��!��E�S��;`����n�(OY�{�Jf�1��ͪV�Ǐ���k[�e���2���	��o�#su_��0h��IY�c���%?�#��  O�j�A?Շ�hq���7
|ש/{a���ƦrmUڕ	Z|�*@��aVJ�$U�g�4*_��'O�@���9&K��0��4�c�U������n���#�(I���ؔp�Q�I��X��RH��9�N���]Z�&q�����R�YՌ�{�� �G)�}�S�>ȫT��U���NS��g_M�Ɍ��؎�XX�U��� ��*�������"���`fq��N>f1����⁠Z%-,o�(��(d���e-��gVs����2�$�SD 5�`�^�1q;���M[޴X��B��q\�b_�ц|�Q�z?�f�ڛKH���Y���Wg_�5���(y�ԃV��3�`�d�\���kB��(X�NYV�Q�&X�]��8� ���3fM�@����V�Y���]K��5���h�4 �x�j���0V��ӭZ̠'(�r�+�Ao���X� ٤�BB�4pu#N��~���d�<��,����<�ӗ'����~50>�j�h���Α��`���E9E� �v��� }����8�[��R�w}j�O�54��x��'�ކ����а��>����M���)�Ml\x*���m��CK@�ʹ�"���t��o�4�����9h��|����<}��A	�I�h��h���Pv��u�@S>���]{�pN oȝ!���jK���8]uR/k��ż�"��%���if�WѦqV"�m �'���
\���b����org,ii�K�����iթU���D@*��EK=�%%I��{���30?�8�z�o� �̚i�Zf�����k�@���`0��W�&(O)Kk��Ns`�	E^�RX�ޘ�+�$��/nƱ2�.������<��<�ĨAr�� �ʹ�'O.\�Qe���S�ͭ�v�3����o �\:].��Q^S� 7��$W���~���l���	[�^ k?� z��ě�g�s�IĴ��ܠ�q� y�Y���sTa��&T��*E+)2���0[יL8�@�wѫ�6�SW�q�8V��ڥƗF���NlW79��<�qh�ܭ�*@.���}3;�l[�=,��0kTF�T�4i��8�ơ�r�����9�������&y�Z��5��Op�A�*���,'3=���r��%r�Ŭ.K�ԽW1�r���DT2���u�W;QoiOZoXW��S��B��gL�mz{P{Ԧ��L4$�{�g��ke:NFt�p�/�.|�d��nr�H�å�#� ���|��f��*V�l�M�zi�UK�ӝ���͕�`�� �d��UW1�R���\Ɛ�/���Y��Z���~�Qo��]hTn�-����so��DTg�(@��פ�\�����c�x��;��[z�KZ6�����oıEw,�M֝���[<m0���oVy�/��j���v%UE϶�w�� ���p-�۞F�v�k��*�.N�t�R>)�
���}�k�Λ��F,�����5J4-V�ֈw8-o1a����8�E����-�.F�����d$6�i��;#� L�:����A���Q���6�' �:��G[�c���Wt�s� y�g��CԔ_c���W��r*���Pj�ʰ-���6ol�����j�.���$f�����fϕmL�ƿ�n�s(B�L��Ȕ�T$Z=�����!;��X����i��g]up�9P%5�53���J�1GcfE��1�ڽ���[�����N�S_O���Ӕ��>���D���;���Ђ���	Z�ã�1��8�mE	��]�kW	���+�����?�p���T��������ih����	�&�	��΃���4p��,������P]��@��z��ط��I��4�a>,���N�K|_�!^�˫�^�I���M�m�v� �\s��A+P��xF'?�,�8#0�����2Z����n`ZQp~YU�b1���T@"y"ސ*�?�T}��GP���6c�SX��9����٬UÄq���D�~=	�Pl�D~�C-D7}GAY%ԍ���h>���pt1��Рw`~]�8�L��.��[�b��_ �߸:�	���:�ڔ>W���/�z#0��	�n^UӇ:��{\PvGu, 4��J��REB��� \pҰ����]�^*y�R%�}"�ݖiO
'j��#���}��P�� ��h�D���`n�ؒК��������Q�[�W.��#8Y_ϵ���t�*�gK����
���}~[sa�zۚ� �֘�,BOR�E�<��B'}���~6&���%&*�:��@Gꘞw�+���A��B�'���F�p����x��؟�:���K�c�F�.	go4��&a$|q���h):�$�Ҏ�-���	�^�n� 70�|9�z5�� у�Mp�*�Ǐw�-!�#5�?�蜹����'�����T=mt��i�O3[ŏ���E�j��&��������ŵ;�479n2ξ]�`�;��La��n���Ƃ ��W��i����ûl�oO�4������?������瓟�jnt�3��-���B�C^_}���D���>ȭ��b���V��o��^�J�U$E!��{x�.u����z�ku"�z�	Lg�	��;�R^e����ڵۧOuH��?}K�T����B�$�����8�(�~�lŕ�Dc���"�w��޶����nt��|�
.|�s�az�:ܚe� ��)��Y�|�����s�\�I��N/6v؁T�>U�P�r��w����Ór�������0�A��ʵ7D$꯻\��X��JV��{�b7x�����۠/����1�'!���kq�ճ��+TP�H���Hat-�'��@�%�;��tN��ܶg]�d�n�V�$�\a�'�S�tD�7kK(�[�A׸��$w�%��x��]�eN��dF5��h���]�h+�9�^��O�4lGB�Y����'��n�fL�$R�s�����0ŬOG��@ $��*
��f/��ꀔ<SyCۓ9���-�uGO�ϓ�<}�%�_�,H��:п�G3 �5�z @�\��)�&ZE��c;��������E�8G�}����\Qօ.(��a廒��m戽j�n�O��B]O�]��PɅ*�D���X!�<L��s��K�Fmds��S�� /�.}p�������"�@�v���?Y��	����p�˘���;�kb9�e~��?,3�%�P{a$�P��6���qE��	�l�Ή!�x'
G�����sQi
�����w���,-V�i�|̫8Uw+����OUi�Ι8=i��a�B��\��X�c�R�R3I4��C�~��9��Z�T)��[z`R�<r��X�P��|�C��6-}Y�?pR�J@��who\�4L�?��OH���� ܨzNn��%r������[l���=����p��H�-�V���_K�Z�)��I��D���O�G|���v�����R��0�oB�#)�f�����N��G��#�C��*�Ω ��EM/H�o�kkH�����r&��ȷ�)wz�%z?1��u+R�CG��j�41�C�]�p�$�L�d55�{�2�mX��Oe�C�ε�Z�.�Ok����ʙ����k�qXʁ0[��趇�^'�0�����F��X�b���V�E�"�E��F\=2����!�.➪�ݥ*,���?���xG���8%�H��z��7SR����l�9�>A@xd��G�o\��7��w-��_�Ϯm�\��DP�Tal���C�H�J����Fğ����@+D� <A
�&N���#�l吡ۆkH�Z�׽4�l1���'�aq*"��OO_�d~#s!?��`J�kJ�PC@,Ę��)M�B� ��~��1��V�LTp1�ۉ5�)���.70��2r�NaW�βv-�W��/x���F̕�!]��u�W���~*�FmD���iKH�S*��V'V�ƛ�[Vx=��Vsl�fy�0�k0IPؖP�f����Q�ueT��U�^�%�!|{
閩i99G��S��=�>�D�Ͽ͜�Pg��&���xQ�R�I�s��M��������th���NoժH�2��/�bI��D���9)���}�z�1��-�e	�������ƻ���Jv�:҃ɔh�E��p�W�n�L�C]�6%1��xK��L�>~D�1ӎ�,�/��*�ᡐ�]�k^�`��ڋIi��f_y�G�B� n?aF��c�&ȹ ����1�FO=�a�J�����)�55�����8�TS���t��f�N�'���`�c3�ؗ���<#W�v�~��,�E���IiQģU��D=���Ho���'l����9�_���"�Z;_�Zz��F�j��cf�M5tlu����zЏ�$�[֦Yk%��@�	<�V3/��}/�Rw�s[Q�>��gtwU���=�@L�=�{�rD �u�
�3�%��c�5)]��pO
�V.o5
�	��b�diZ3V5���Nm;-������lЉ
 G�697��Zv��X�c�SK��FL����Ex�}$Ɣ�@m����7H"��΃rV݋#b����O
��F�F(5�N��2���1�K�];;�GX�T��bK^x!��Wfz稜�{f�U�_�!E�Zl����621����d]6JD}m�"I�0��w�vKV`���y��<?!B�����7/6C{���3�	a�g���m�Hu��@f��L��&tYb�����
��x�S�Қ�y|�� �Lt@��
[Z�/��;���9���A}y�����:Z>,L��<V�<��h������D�T*��LZD6������Q��L�(띉��p/�*�N�ā�K)S�ͨ������L����om4��0��>���M�:�WtX����K@��L�	���̖��uEc8O��Kp�z�v�0�N����I�1qb������o�s��LT�JO�豏���8X5���������]�B��Gcu|h�N��L(6�����6�&�{��y�[y��V�8�E�>{itLs�B綒�k���k:��5�Y0�7�ďhA��E�x[2�.��ó6Cqs~�y��1�[O1~H��)���.�;'���WFʆ�I����L��s3`��Ճ��>�̘����30�����e(��cz��Bφ������6�H��(.�龒 ���|���h��.��0ġ����wu}V�3_��*k8�gej&�(/p��A�ƲuLc���?�`4թ�k�9��v!?��*	gp���m��|��h�d���q[���o1�s��d_�o+}qw7K��p�>����WP�����A�1?�]Xd0���g��	����/U[���{��a%H���Mt��D�����&�����0�@G�@����v7{x�w~-��*^��?��;����21?��bY�$53����j���h@Q��)����D���s�p�K]�t�����0��5UД���,��oLzk�F�W"m�#>1�Z3Y����`(�]ÛQ/�D���I�����m d����h���$ǯ�@�M`h*$�ax�
ꅇ%?�s�qEw��uX����xG�����C�[;]*�n�?������C�~U|Eg<�=�+Yn
��)��F�˹���h�v4��YAB�"�=�[�YO􌥜���A�쏑n�%��9�A�s�7���6�Zi(+nB%�-���|f~R��3�W���Y-�GY��0o���}L{��唲2[��1B���o�l�u\�W$�0BSEa����������>d����,]ை�VvE���7�/xN�h��*�v=@'�I3pՃ[0�!m�Y��v���K�/YH� 9*7���Y�!c���3����K�4��b�$=F����>�A#����Nk�5[Q7��u�\��I	D3��L'=��8��K�3D9k��ݗS.�z�J���V4R񫅄h������6�k �J��d��p������;D�����;w6��	��A%��K�����C��X$��:Q+�[����큱~��B�J�����.��+�9R[&0,�MLl[^�l���+2�<�7S%�onwi�8pl�Ye��˒$?���{/�l��z�i���7yQ��ԣ}Iꀊ/�������A	E�N�)L�
T@�����^M�2ȿ�GmJρbe�Ի��߆�𜈯���![Q7�l�8�܇�c���X�enO��t�H����O�D�2V� ќ��ך�N��9ߒ�cm`N��z
�F�x�I�{V��b�_�ڤbP��]~�A�F��`^d�Yv�<�J�tE����m�� ,�0+:ʺ���r�sP ��z�DA;�*�+m
�x�� ���ë'�$Hj����(5=�����鿊)��e;�>���RD�]V�N��|���8�j���*��e	�����c)jK�����<��$E`�7�
]�߬$X�GDn@��h�g�,(�S:Ob�"I��v�߃ӽ�6�{ЗX�:/���oڂ��Y�h�W����Tʰ�#?⾞?���Ox��WD�Q�SH���a"&�F
��04���J�`2�3�f�:�Bӿ|���^=���c{�P��=�-\����T�K�P���U�=d�ǡO]�Z��>V6�Jf�V���h��=�&��o�oG�'�!�3� }��J��#�x��,�����T�g_a�\Ex�7y���d��p��f&��ʜW&TÌ;.�Cbp�(��D�G��I�2{ޝW�qwf�tu�c�a�Q�c����#A��1v������]�F����ֶ�>���1J�D�B�
#�5�3��>LA$:ýJj3�a"��&� �<9����~�.�_�i
�¯}�4�rF=\����S�8�j�� E�BE���T��Z� ���E�sW����Ԝ�Lmݿ�4�s��SM��[��n�����ώ؛z��}�Ĥ��~F�v�ã�:l��0�%kU��m�a�7��ʉ�e��gs�N&���$%8��V��t���W=k#��,3A� �%��)I6��{�����ʌk��,��*����W��r'x�(�u ۹�
p���"�!�D1\?������TY������1/-��MP,@��T��I�$��݁��ۻ�H���tʃ�[PrG�|Fu��@:�\���צ)nֱ�4���4����OW�~��f%
�C^�cg^�"�<����Oo�m��tl)�s	����/�'71��0��Qrs���9���hV����X�F O0B��]�ϳ-�%A%��l�Ή�����JI�����E&�ê1=z�I�(�Z���v/w
�J��`�X����8ۢ������0�bފt[6SI(+#3��:����'��5�e� s�p�J_=<������d�z<&(��z��-h�����B���R8	G���Sf�U?c?쭊gv곷�b�W}�72���P���-R���gk4bn1�{���"0�Gl�诸?9&
�'����������}�XHc(zL٤�܀9������~�}%�xnS���P��]�
x���PG�%��mM�c���N{�~4�V���=�SGF���B�z�rY���R�P��YT�h�����|���o>��W�����w��l7���!�Up*Ql��H�����J���CV��ǌ�)�l��gRf: �W��Cxq̎_��VP�/η2���˦��a>�7a������Ab"���b1Tg��W���L&�r ��_p蠼D_˙�{��_V���D?�i7����� w���#�3T6�$P�ؑ$D���������$�9���8ƿ���i��3�"I�����J�Nn�F�DLGw�Μl\��A�G>T��쯒Ha������i�@<]�xs�v�s�Q�kK�=��R��U0[�}��	��a;�V
]�8�E��=.`
_�?mt���F����~E�Ƴ��&��i�@T7z!�%.d�����>s֍����$�����B�����&\�V�g�Y�X��Ri-���Ѣ���eh�]��y��+K~���8���}�Rr��}����n�h�l��e�`�G�N+�<lW��h2��)n����4��|�5�~�iS�>n+�3Y�'�s�Zz<�F��0��Ǌ�
�����xF ~�z�����>���\��~JJ0�I�p=�I*osˀ����;O3.��S<&�pT�5�UƧ����5MI�1(������˖��k��rG8��g%3ؕ�d�����7o��$L}so���+��ylR��Ȅ���g}ٴmm��_�qٕT��q.x�&a����D~����; �o�|���j3��l����e�5�t`0����l��_��)�v�<y��MS(�^��K���SRD��?�pz��H���wJ(��&�|���KȲ��?����+�i�(����:��@�u��tt"�y?uZBS�ۺGF��}�.�ip�rո�7�Z.6���'U���	����~�@o�c[Oc��y� �~;L��n{r��.��q����wo_��>�2�l-��.���5QB��Zf�=�&/TEa� f�T_$�r�f�P\�����6~��	�+|����d�>��K>��#�9����
a���w�&��]���3G����YEN�S��,�H颂:�/<��1��=F�;k�n!X���ߧ(����ۯ����h3����K]����L����	�|L��D��"�*��A�ğr�K���&��b��cayS�<�hx�y{��0�dj����r�����T�&��T�"va���c� 3�ݙ	Ϲ��̥�e����Ư����z��+#H�\#���Et�o�sed�h�oщϪ��~��f�IZjҥ9�R�y[QN�#�a�љ�v[fu��=,?	RN���z�#��R�_��T�O
�V��L�ك^G`���]�4����3�V�,k��a3-�D�P�*ϓLr0i��إ��OW�ۛ�苌���'�`������j�1��6\�w�Z��bUn����F�i����T�|�!��e�,�총�9��h����� )
ٹ�v^���b�ouL���_C��/d�	�N𖷸+M4=$�x��y#ɊrZ�ϛ�~z�ώ��6` ϩR�V��ئ�����]��H��j�����y��b��%�hս�&{��f �v4NgwՕ��'��%zf���y�>�\O3en?�-#��CL{����}p���zf�H������~h�q�\Zh >�{U�_G�3W}�O=�����G�� �O�z�ʣݹ �?��_�_{QILO���M:teX0�-`G��
+_�u�ɵm�-��V8d�61+|҅�(��CTT�/ϥ0�	��w��
����+�#�aTf��Fp���t�x��z���@��Ẋ�P���=��F�F�6ndL� �*_ݵ��K��ug��rXj�{ ��89�ig�I�������:�(�,�A(kʣ�e�a�P�+�cr'���x/��\c��4-v�Ry�'Eև�%�-��Y ��=F���?NB�߽�/s�Ym�
/mR匟�)��t3�<�m9����*
QY~/�ߔ�~��d�&���izL�WR�2�x��z�.[ �����|���$��}1K����.D5m;8?bYE�Ʊ��N�Y؞�Bj��g����=�e�S�V/D;��"�B�&�,�|ѾA߃���tg�|�5�c��fH�g�Lw�ՠ�Arzo��p��l"ʞp��n���oad�_��;u�3��JT�u��^^\�ӹ���l�v����-��.�Y�~�vȴڹ�e�\��y���:U��P�;Y�Ov��uw���Ѕ���ET�My-�<�5x��%C�t�AR�{��'fd%�E�LY����Ox�ޝ�l�i���6B0�[����L�*�iP\�� P�G�|�f�X)�Ku��E�o���7��1��+/�(��$��W_l�����$���Y�/�[���b�N�<��Ʋ��j���1�8���-g����,ۓ����Z`�!��!!��DԹi�Y��b��MN=W{�_��[�� ������((�}  2�I���<Z��B}�>�ϨY��LhRq���1%ҕ 1�0n��v��7^縡�Y$��Jt�5|j�肔WQX ߙ*x���΢%x�э����ے����d���j�w&����b�^#<E3����W��Q��C���C�ee�������W�X���v`w1{ZզqoF�Oo�8@����F���B�fQ�c���
R��@�������$f��N�Ùg�h� ��H�w�<o/�]E�K���/�9��3hŧl���f�dϧ��Asq�#�Ƣ&���-��˫����[-xklEP]��iG}]��ZT&v�2Ep��M=Pl0>����.7V��,�S��m�ve��f=]���V��5��5�+��e�!����(*�#b;�A�_�s�
��$C���L����A�_$[
�)��I���^����g _�D�b�$a���MΤ��\'���G~]:�7��w⫍�/F�� �����j��v,-�|���RJQ�6P3��1��Un�����V4�.oJ�FD��]�>H�^NL~�5{i�t��C��ΰ<�_CU&��pod����i��[\��]�n6�{�g!l�ĘAQ�]:W{_��0�}�:���\�k}��	-v�E�K�!��I�"�Pn��P�c4"���ՠRJI Y�[]^y�@-?Ct
��_���(c9��Q�h�ն�`Zf����D@Oݱ_-8���'0�ʫbD͇?�V��"�o�ͺ-/���
���ŷi@�{�e�$�K�p녔a�60w��c�Ę1��+�~�l��5B�z��'����f)�J�ezQ���`a<9Ъ��=�ƌ�|�v�^xW��UA�l9.�  WS�ߐ���}�fo�������b�m��7�!T��˛��eѴ���Kݧm*|�e蝙��vL<��(gI!���V���n׶+,�Y�gi�}�p�m��C�<���,��f�T%���Z	�Гl<�rR]��~�~o��x�պ	J2蓋H��t!��U:����6�M�h��ׅL�$n?�u;M���.'�1�Z���˾�a;�0p����V�D<���<��Z^��-G;��m8q-��W�:;��ym��p� ���$K�v�Ȼټ�G�t�uIْ�|��#���A���e��N�ohGQ�h���I�?G�窦�?B���������i^(nB�B)�� �H�7���|D6F�H(
�*\x�͇A��3�Ѥ��Sh�h^����R�����CB�<��L��˽�;�ӧ���X ���߼��E�l�|�L�>��+J�r��ؕ%zHY(���#8�@�4���w09-�L�1\�9LL��Ar��o:�[Uf*���$���I�Z
ʠ�k�shD��+g���R¨a> ���v>�<6P�uLoܤ���9)����p&q*��-VfAH�l-�[-JUəd�F�DtIfh����r_�g/3�G���c�N&��8rD���(͜
m5���ik�/��l�:0��W�<C,uu�ew1G
�|!@VG��*,X�>!_�)E��eQZ�^B9ڜ�3� z���b�<Z��b��G�� ��x.��M�#ѝn��8�NkY�ږ�C��q�w|�����D4����D��gJd�Z�B:��%�	���r��&�mf$���=5:�b�R�^YY�f�؉P�X:1;+��X�oЉY��IJJ2�T[�Lh3�qPj��[TE+A��-���"��$���1�JN;��h����بHQ�I�3Պ�f:j�q��f�Q伩kx/����p��~V��Ŕ�t:�&����Ml�WL&"�Z�P�巎�Rt�wXr��C�S�?A	:?6�4�#���6`�@`��Ԙ	�J��[�����̒
����בm����t�M���J�--f��޼v�y�D<���Ep�j��d�-U�:�
��u����\<������?
[ʩ2T���	zFA����vJ,z�����/XL3*QlAna9m� C�;ۥ��?*�X��91�0)�O��y7o�jy�J�vF��
�`����#A+� P���#�tu>��cI�_����	�|BZE�x�|%����9y���f�`9���}���\��3mo��6:o��7�r/�Ρ�%8�6�{}��v<t�`�m�M���}#�|{�\�QEm=�)yt(B{
�oz�Y#9xm�K^VcleF@�����p�)'\o�Ґb�n�����%��������&C����2�2�'��ѿs&���.%p��18w�?n�1��πN�����Ll���Ή�)Y�X�Q?�e�:k�_�4�
6C��Ӑ��談�!w(�+v�0�u,4�����ɸ�}5ǈ�3ֿ߻�ϴ���� &��ޡ���X�@bůk��gm���r��*e�%��"��J�
�����h�:�}w�ž�����ȄNpN��;�(�z��T6 �S�o�ɁMrT�|���5���������<�VlV��4���u������0C9���{-fY�����"Ļ��*��רeA���|,M\��6`��h��L�x$o�:�5iA{9_�8�T���"�5�J�r�(o��=K/dSd�B���K<a�oS��?���J|Q�v�ll�^�	��{w�ؕ�����hOE�Ԇ!�@��4i�/8e�Xs���JX�IN/xª%�0��e���a���p	��@��]2��<ޝ�X��p���=��ضX>�V�}��p���g�F{���aP(v�h���q��&�X��#po�C7	���P޵��`��/��ˌ��IV�: GL�
E ٥�b��^�0@u��374����	�t�-�c�tbd��%�J��]�jbG�����<� F�r��z�cR���zBQ���SK9jO���zMa�f�wQ?�W��Y�s.*�{
9������K������k��R��2�fb���U=jػ��8[Lș~�m�f�R�汻�;�#+w�.H�.��>)�kWв�p����(�Y߽��U)��G�	�.s��2J�����詶����2X�����h��xJ]�벡�/��N�-�=_��$#��W׼9�K2�3��e�~G�dQ>�ݍ����I��gsq�b����l7[�,��P72�o��2^?�H���Nh�)y���t�FJF��:��R�w��eN�8yh��Q1P��es���3��
��#��Ô�C@%W~ρ�Z�:f�;:pvj�+�S����1{;aċ��U�AA��`�'=��XO,�$,�q}��4�͠�EW���9�t<���Z|�N�E�y�	��F[�
%�]��M���O�Lmt��=yHz���긢�WE��ᅕf�� ���ҿғr��Y"2Kc�*>KA�����v���o��2_�������.�Օ��m��m�Ů$��
���ʉ8��� ��B�~	y���}!��n:���@�g��x%�_��D��y6l�P�E|�^�2��� 2v�EZ1�B`�jO��=Q����� �I�#����!H��3?,��ځ����7@9��/�'� QV�3�|��^��pyӺZ�)�i��_�N�� ȦW�߈��+=����J8l}:�A��5��%��W�P�w1�2<���U$�gD2^z�e6����9g-�cq����<q�"�R��N'A�g��3�xǞc��!�]�7o�Uʶ(��H�%�;�Ck?��PPs]8j ΅~��u��a%�~�׵��^����f��xHno���@�-v+�W����>'���v�VI�,�{�v�D�P3r�Ke5&�ˋ��i�H�wôL��:q�_�B��p�,�w�NmV��'���T�7��Dg@C)�߸����՞g����� ���tݪ�����5���ݏ�3�k�˧̹�=~�k��-���_#�7������?��k�
h�#�>І������eK���3Unڢ,���-��V�H�ټ+"����u@�/r�Yv'E7��ű�`�;W��*��v:�c�|,6� ���"����7�w8���^"7m�@z�q=U�ު�i�T�w�*Z�L�5xJ|�kJϵ��-8��1�������o��n�iقY�������pB�B2�IU-�"��Z�d>���y�LTǦ]^`��?�)��x����N��2���ȳ:��6��XJ�NT
��FU? �]<��ߴ#^��Ik��^0���bf{0��r+����萧<+-�N�@2ʶ��6�&�����	�ʢ{_�V���AV�L0��'��pv���^�N�@���<��a��r5!�X�\�6���ei�R��|�Z�n��VƢ�c%�R���7�����9�#8�RB��%�W���~�.J#�,��V�cX�D���U#�n(�m��ʄ�P�(�a�D8�.��������h�*?j5dm)��!RvcZ�r��u(��rc�-���&��B���ֆ^$S�oj�8�e��ENa���x������K
k	�l�.�5oS�sr��&��A�����`�f�-��8�_�l�	T�a�e��k4D�%"���=^(-3��v�/����E~9����|��p����z��T9��ǐTPh:�:��y�B�%��R�`�,�J�� >1z��	����KhހV5Z�KW�]߻Ǵ������=��Jt���iue;?~��-V�g�j^�4�i�[���V�/e�1R먡U�C�L���@�✽C�Y�~��gÐ<�u+���v����Eb�	%�{�3�Kg�Y�;r/Po(�=x�og�KĬ;KX~qG"�96b.��?v���И����$�'S��@m�,�=��(p6C;�!�8��L��*���]��X��-��
�Ϻ0,^\��<`8X���&}ئ�@��K�\�X��ǜ�6XvڦCj�ܶ����ty�1��F������W�P/�"�q ��������e}V "΁���'�]']L�s��1~�_)[wa&}�����ΈD%h�徣�k&$`�1M=��B�6�&89��j\�c��Gtf(��h�!@]QS�:�����i���{XK̫]�Uݺo0$,#9i�ur�d��������K��
K��fp��\�#Q9z��8��\A�6B%P�i_��˿�Ra�����%%e�-	�|���4+#��M�~i�iH�[�·�fG�p��A1z/��r�8�H��'�������i�Xؓ{2f�9�g|�u�����Pw׆ۧ�z.�����R��V-Y�ŏ�q��/b"*��D���*RI!Z���ۊp����Ǿ����1�ZR�d.)3's��ku��)u#鞘[9߶tu��(�>+q�+<^-����+��K�5�F���^KK�Hn�MX�X��ҧhJ[�������^��;���M��#���'`�B߀�]HȰ횀����τo�A]-�,���������I>�A'�t*ԑ��h�����ۺh�wA8������	�U,�hz4K]�(Ҭ��ⰰ�)��g�|٨��y�3�ϰ�ѕR6�7x��u�:�\"�!��+�	tX���DL��i�ݹ�O�Z�t��;m'9v�a�Z&UF����t����*D;+�_1��b�02x��P�!�;ȴ��_�1HN��P��d��~:��\���ou�,1y'e�9�`��(�|,1c���]]�����|1��(��ЃOȒN�fx}��=y�5�|x�'V��,���
�\a���-���	޲g#�FCLlo�Of�W0ў�׮�%���;p�1��@kj�X<a3�)<� "�?�6MA�z��a�<�=�5)��Ϩ��'0��'U@����+<�.	R��w�������7�n����*������s���ZCժ�ػ����wB��RnJ��r���.3|Y��0���c\�f+}�$��8��ĨW0珐�1�d�z�z��m|��<B���J!qv���	�����tG�������~ć�G��Xz�#��_�6��$��>��t^ Euk6C��O]� ��,aɖ#[�.ڧ4`�4�!�y��7���Ļɘ���z��2l��y�DH���5��o������:�c�?��<�T�Mutr�I?)}��v�!�Ú	�GYW�:���#�â��%8�-x*Q�ţH��X9��9���؅���0INhM�gb��%Y�O� ˙ Dn��8��n�/�gY��=�"Ǒ��MS���gt3�(�j�T�v��گ�FX�>t��iyJ��6��h���׊�^�k�籁�Q�����V��n�&��6�⹪���!"ã�ɛfP<{�J���_Hǈ����Y`|�Z/p��H�������@���N��ˆ�'`'�C,��gb6���H�(��a�V��z�'TY��׉���Y��E��%�K=K$�+�������k K�����5�
`�~�Y-��$"s����>ٗ� ȅ� ��eT1���.%���!��Jp��>/���>��8!���As���K[��g�U��{"�����'�2e*�]>Q���<Y������x
�(}LH�5��ۡ�$"�R���aᤖ���dL��	>� �m
��s�?/~�ĵ��!ba���ɔ i|��V��=%D��3�MC��Q:4t��?_�l��f�E����}�E����H�~7�yE䕶U��M� �V�?��x.�&G�3p�p-e,G���l���UD�-�w�Yh���e��%�����_���8\�eĻZ�#?o���Nw+�Vr��t���>S�IԤ�@t��a��}�-,"����st���]������M-��g$���%� ���E�js���}R郓8�ճ���8�Z)����odp�ct��J��y��ے?4mq@��d���X��[_{q�X%�݁;:�X�(�_g���U5�������ui�*�`d�(���>��*6ǧm6A�~��Lt(� �*���BKJv*G�y�ZE���+���$�p�e�T�g#�wh�S�D�47]@~��6ؖGZ�>��咯l^�$@[��.�����t�J�Z�c��x�.��K~�y���"#7㞆~(Y�0��M�}E|
�T~E{����^�_=�(�M��N�_<ww�[;"�#����m25cCn�����]�cG���qԄ�&��WA��O�fѳ(g�|��oa=f�o���kDIl M�~��.ěB�Hj�6��!N5��*�.��A�z�:R������T�5�I�������E��	�C)��4�%3�����wb��$-���5N]�t5�b�Ē��&���M�~�~���ZA�7q�k���cS��,����y fŠH���>�e��Q��8����0t	Ew5�^�/ �c�@gf�}�5���/�N�74�N�֋'}$���t�s1�9$�.�ΐ��`�	G;'j8ɚ;n�4HG�2p����7�.(���<���WW��t�V��n�|��h���
>�[�.�0~�j��tm�h:�&ZS�fwb^t�l�Ok����i��58�9�&�}ϧ�	XiT'SP�|wȿ��e���կ���;�5��%K�SW�q�������ͺ��.���u��N+��!6v�{ ŭ���u�LVs39�)mK>n�B�Y��X
�('������N82�6�kkߦY�c�*&B�D�
ˈ{��ls�c`�F8&����q� #���K}ٳ}j���z�m���y� o�^��3~.�����~�Juf��Ƥg���*7��3f��V>B�I�}����o��^ �D��5%|��Σ����\1�3��	<�G�1�����ʋ���D^+\�[�+RiC_�O�<D'6�e�ꒌ���[�W맕 �r�Ro����jO����E��秏�^��S.����1M�o�e~_y���̘��P�ms�t)�r
#1Uۈa����XG�|�!�j+1�e)9��Y�CQ��D'��0@�_�� �{�_�[LPJ�T?+�˼��k8�<ѻ_`.���<�>~7зf�`�
��@�Aq�`F1�O��b���k��P{�9��eBA}�g������~V�NFt*QC�����!� �\�^%#�RO��Z����#vuIo�<�<�ե;i$+]�ā��}�>1`�'z& uԖI�S�3f���^��OK�TFU���	�-VY�(s��m��z��I{Ge-���!5�׶-0dp���߶��M�π�m�S���L�F5:�r�L\,��@�[3z�y���mօ��;F�m��d�8	�S�h�E��jb���
	���>9�y��:rfP�{/��/�>1��s��t#�g��M�&Ë�s~�^_3$s���3�Dz4q�2��F�/������v��������W���::I�w}�������G};FQ/*4�X�=]5=o��/%71m�������$bN��@����➿&h�\��?,cC�o�F�*85>%S&�U��nã�%�|�Ҡ�"1x�wA<��v���3�&�Y�V7D7�)��m<Y�Q&/ˣ-�h�I@�-�X���L;o�
�2~�}ޑȵ	�1>�����Fb�&�<)�(2�N��kE?E�s��X�V�l�Q�_�V�m��'��b�22���XO_�[�N�ڿ�T�U���@�֗�Q��F	S5z2I�	1W�x5z�(��E x�U�Y��_fB�V9���ί�vS�e���;����،�jZ����#Ɔ�SVi�gԧ�e<<��=�wJ�?ޛ�z�tK���dP`�M����V�kx|�H�c�A@F���׾�g�2��,<�z9�����=��A8��v�1�-5xF�+Kff���7��I�UICWV&cDz'�9Q�P>���yT�v�z� B9�uc�F�c	p�#�b ���iyS-P�.�!�W�XmFv�v����8ҶS`�a�ud�r3-�3>肄�