��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�]��Xȭ��p�oȡ�;u0ީ�^�)�>vys���2{�L�~|c_Iy�K����-��9!��\�Bi�D��{�Ԣ��r'T��NjH��ဣ]��9��|p���4dտf+����ؐ��7&Qa�z���m�ࠧ��3`����8s�=L��4�S���J�7�h��J�3�_�������p�t_3�ѹY��S�!����_-)�_�3s&��������0�:pzj�MG4�6'1%ٌK�93̵�8~��L�\��T�Da^@����i�|�\�) W�T�}��h��ЄY3����U�m�ڞil�@ƶ�K?���_7�<v��DVZA5�k8�+����m'���9�v�ɏ.|�]{�[���&G`�T	�~��L������C�
&�P,�;w^E�kJ��^ hz�����+]��boOm՚��̩��Hb(
��ȹ���Y��Ŝ�ޅ'eHZ��jh��܆��`>�>t���	r��s�p��q֥�#�����|�C&f�7q�0�o�?��Şd~���;dk'��y�&,�ڔVB������g˨�',7p�35���x�޶�9��4������2�Ɏ�H���B�K�f �@���0�7���QӨ�_�6�qNJGV�� ��^���o��:����ق�`����V�W�lJ�iE�/*�L����g����+�]��mZ�_�ia��f��'	�q�,�(G�({�>n���+�Pϕ6�چ��N��aX��`�B_��"�CƼ;^�mJ���0	��l��xqjP��;��w����;��σ�iu�\�r]{�%Hxn�������y)P�0`^RfF'>�k��E��_(��H���`�@���o������o�X~�y��':[8�.�nW�;�X<���N"�4.��.{�����nŘ����ҍ$D �,�*! C�I����%_����6*�/�Uk�U
�#����.��,�f:-��W&��$;�s�Á ��_\58uRM�f1ڵ-���޿=�"P���Q�$|�e���ͻ��Z����h��O���w;E8��ѝ��e	4�����
��SF|�j���'3��,�w����CW!NI��S6d{����춀��(3:��!!���&���Wf�u����fl4�7�S�7���B{ZYL������{��D\+���p$�?ϐq���q+����tq3-��w�2_"�$��J�Y���h�Ve&��P��
>H��
��2i7pC���v��yg,*J좝V�营�
�p7�� &J��qi��=���s�+ZgW�:�*�����m V�_cj5a���hl��	�YDp&��P�k�'0��J�J~�t�[�.`�ki�]�����$�J����&��b�lOh��u�s ��r�N�8Z�ǁ�r-����[#��aO�=e|�r�F2PmƉ�j���
w�v;)4�,��$.��@���-bA�Ec��+��������E��7뱔�H\�\�%;���[.�"�!]����gtѕ"m�ꊥ����I�j<d1W����GZ��4�S�5JY�qμ�d�	/b�:=�k(bS������
�P!j
�<鈱��sN��״)I����=i�ƾ;~��%)�к\+�25B`��8E,��U~ϭh;����G�EJ
K��wl^�?���F�(����G��l�MYQ)��[�?�����hO9dBaeHoE��= ��a痎�b���0* �����&��,	\i�K����ݥ�3���̀��-(��c�b�J�p�C��
�B.�<����g�"2^}*Ҩ���p���$t-b|�a��61Ğ�n�h���s�R��� �>�����D�����v���0'#���]jp��\3�:���`�N��Z���{����(����qt�`��Hj�Ξ�Qʧ�qz���J[��s\�xt��|+jr	k���LM�h7��/J���	ԘE�{&�+�f��}�>�)�b�j|��K�1��Ob)��)�I;W�Ӣ��:	G�����+��4��B��8l��U����rgKb5�����P��Q��(;�&ibV��I���$��a���N�lO��,�P*��6g.��}�挓NJ���D'�cM�D%�	�UJ]�g������6��%ƿ��e1�)�-ݦ[W%���� �]-%Ӛ�5~	Bd�h�T����8z��7#����]���&w	_��OW�(D�(i`��Gzm*&F:��C�le�x���,�'u �~n�z-�����樹ʛ�R�:#d����k�q�����G:����E�����T��u�	�1 ^�^y	zlc��f�`Q�$���>��V,M�v7�d�����QP�Y���K�1�M�=�ô�v�3@@Y�OIR�t'�̿{��9���]�@g�	�LJ @>K�%
�_���^
��zY3���Z)˻X�U_����2��:��H��ԏU��s'!zP
�@�.\46K�|y���$K��j|M�3�:����q��3��L[u�Df�l�Sh��1X"h}S���N�wh��u(O��qM��A�G��CD+_������m�*�cVKT�'+�v5s����>
C���?� ��_��V���� ��1cL?6�}��Pp�6�т
q��(d��;���G�U���
��>|���+�y�����6 �ݏ�`�Fn� ~Z0Qt�����(9�bnRm���.�2��W�<ft�a�;ޱ���N!�飧@�HP��Tw��@�+�@@=uW�`���+��N���a	��Yd���G��Ko��Χ���z�n*}��t��	Xy�u��;���EiA<W�ʬƃ�Y�� [v#T��#�2E�	����l3	���%3��\
#ӹ�p��Ka�0�� ڢk��)���C�,�xGT��\J��X��K4V��򿒗|_�VFa�
��ZkT�\�������jſp��=�l�*)�+;{�JL��v���v6LlI����q�x�?�����Lƀ��,'
�<�W|� j��KtsB�.�O]=�����$\)'�v��S�g��3F[�p�U��KY�{�?Jzy �T�wc��L����i?�m�V[�V�,��V�0���ֶ`ɉ~KZ�m�h4��f������������n���%N7#�P�q|9�4���`#v-ru�Ջ�@sP�\�x���I+��6�^)v2��x��E�5��iĿ��?��^ǲn��ۍ:Ig&���~���۶����S�S����o� ���jS�̚����հ�\�M���I�,�Ԥ�^�ؑ��w�qz��T6�psNb��d����%�cX���{q�Q�=|��A;��s�q���΂E�e��Wm��α�`-�c�.��d�aT�TW��,O�8ΩB4լQ���X��[\��+�����t�iFƉlF�wQI��&�@]��t��k��"��2�v�g�%��+`P�f1o]����SI��f�^��2_����) �1���ў9L9?˲k�Ϸ{$<�}z!H���{U��hp��]���^������E6O��c�OX�O4����۾@{�b{ʰD�����+�I�`�d�î�_���wD�M�e��?ѿ3yТj���9��W	��'�{ZM��� �b
$��:�G��
��1������J�(����wG�?��$i,�%�4$��1Z��M�x�Ex<F�R����3���S�=�#��m���`	���g�$�Iߑ�fu5���)b6yd��,oe̴�I��w�����Ֆ�9)L�7=�3I�:Z�p�cc��� �	��L�U��r���n5g��B�Tt}�״)��I�\S+{~ +��F*; Rۦ�	��ߡ>�nbS�<n�U��b�cN�79�� [�2����h����+0�}���t=�wk��lm�£���ٴA���<�_��o�Q��[~L��ԗڨᯞ|�4�ep_QZ���Z G����n���j{ǭ��~^L�+�ou��&�~��Pl��X�6~�7�%*��3oQX�.#)���-lC[����W��	����.*���u!� ��X,G��Ž���骬��>�z6���0�Eu���U�7`r��Q'�p
����*3��O���<'���E�����ط�eҟ6���7�?�G�:"�Uw:&�C���f�~o 4�~�Í]`P�h`�]�(�v�yx���+�\�d$��+tM]�(�&J���H%?4�f=Jm35�&ܩ��Q�Ο٪V>�'Ֆ3-��ʛM��V��)�������Qd�f��OH�dR�)�,�r�i��|�"����\��w�ғ"&�>nj�7��S��`n���q�BD�(���s����T=�8W�@�W��΄)7]��$5���|m#I�W�5	��,<
��U���U�1QOui=C�^��H���rP�%E����tB�M�rC,����@�yL6n�'�����9���i]7���n�p0�s�+�&�c����%o�H(m�_#��y��`d,�Ҷ�8Ga|����1��7(���h{��ߥ5HX�2id`���`�����+]WKy�"�l�zS�Q�£k�͉IN��F�՛{�o�'>�.ƾ��Ʌ�(-ꛮS��Nm�OV'�h٠�l�v���v"�-��ߝu�.��sDsȲ*�Z����æ��v�'rr����3����{]�z'6�;�p�1����R_(	"��� =���'�y� �"�Q�a�D1M�˫!��¸a{��c�11��4����I9+�O����=\q����n�>�N�V���i<�ɛ�Ol�2���mA���{a�P�D�[�D�i+�?[��