��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�k�۸�m�i(b[�{�㇌�]�i�5'�`;Etg
<������H�W޵α���N-�`��6����ݾ�FF��eF4��_}<�ےA�[,�|{�?r+-��]n?���A&Q>�Mx�E��K֎�>v"wTD)3�2C�
!h׮X�L��,�_��ZS�}Ps��7�F�=������>��=�.G�Gר��6����<u�ot��7 �ǙI�QK�(��%$����q�k?/%XF�;8���	�6:��'(���k�Nh��m�G�'���G��GJ���tX���ۜ�(/%�Z$y|�`�*ݡ�E�$��T	""I�z�|��Τe�9���=���0���  ⽈��6���"O[��@�㿆�����m�QԸFO�;�� ��\뎵+�3#V*pm���Lc�\��I���� [+�-����^�ۤ��GU�ş�'\<ZS�OX��տD�b�M9-J�^H)��\eo��V R����˽|���u��åf^��Ar�h���+*ێW���m�"+��Y '�"f!4�,�k�l��z�B>��[������H]7��GIS+�?ny;�[�%�X���
"f���T ��6�C�=1D�x/sY��`Dj�ȝ��{��l��D��ɍ�����N�J房~�S��b
��&k߳�rC�9��X�_R�����LKu���r��j.�{P�yA�+���1�׶���� ����rw1�G�Hf���s{�r��X%Q��]#�ٛ��S.�j���^�)jv�����*������U��)mӥ]�P����0
p_ͬ�{��P��&9�sJ�J8x��v;��ZU���+"^h+���h��k�{0�d�W��f.�R�7�*�4tk۫sm��J�B��;��
��*ǲ��h���#�r4y��?5O�Z,�t�,�T�Ǆ�������6���8l�l�9�+/V�I[�(|#3j&~�(��VYܐ#�"C���p��ݟ.�۵9��k
UKnf�E3���we,րC	o����'����[`2ܮ��Rѫ��b������0���o�K�(.�l�i�Z�������^P��3O��ɡ�B�~�12�������G�Y38\�K��3܌���J��;)̩}��� ����X1��L�4���˻+�N������}M���t���V{
s���*���1�pg0�}.P	���������hZ��E�y����|��<����>š3���^�Wgc0���Qsh@�`0L�C2�9�ȗ+�PX�^Hv��$U��%,vv��CPd)��*hE%�L)����d��~ͪ
��K/u4��$�^Z9�3������=52��e���i�7e@<o�~��ƴ�[ED�_��φ���F�Ӝ��Ɇ.�	��,OkرEw}��	 �/{;���I��fŴJU:�Ⲙ�ě
�W����G��|v�p�䕘�k��	�Bb��iL���!UR��Kd�����w�`֝ڲ��ǐ���_��F��ܹ=/�k�3Z�Ia5��R >�������sWm}�yn��"�8��B�҇�FDE<q��3Z�P���8���k�N]�ب�$��u�'6��3���G��
ʝxN�^��8�
���"�'