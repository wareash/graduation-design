��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jåا{�\�u�?߷�dn@6�zf��r������;�O):�l��f_l�y��H�8��kM�cl�h!�p���w%,�
��`7/�y(�(|�0(|ӯt��My�AG}�f��NU�,��\��6���������.���x#Bw���7=��-���N�e�}1��h��>y��&���o��Gz���������S�+瀒D��ƙ�9�E~��Wt�~
�H��Xŀ�ɔ��l�G�� Nwh�jh3��I�xk��&���b�J��}�q:\�J�!�H�4=tV梷*=�-l0dk0�56C�4{�^���*�q��-1u���W�������j�*���Co5�ϲ����~��Q�H�G�L��	9rls��t�j'��8w�8��oD�R�uM�j������逝��+�٪�
�=99��V�A���v�^9IԄ;ZW�TQ=Q�`�i] }������B�^�=����EGE�G}�垞A`a}Fi�$S�%� ��=b�/��$h�`���~֦{�����z���u�(�B2*�Z��/&�[�l�4�!�j�Cw��C�`�	1�E&]A���f�A���Q��yV�Ĝ9�֬�����-��z�3����X+�{,�E�9�[�Ў�g'P2��]�fb��E���6���8�&�L��Q*ם��i��XrϹ��#'/��v�L$�p!:��}�k�n���$ �(BMyn��s�@�U1� \���ا��j߈LF0@U��NC�+��� �l��w�C"6Hfl0(!H��b�X���rm�{�^�1�Dz�P�R��o��L��.�aA��y#�S�=O�Mu��j����T2����jE��fM��x�^:S9G&��oݍ\������h�m)w�␊��� �6���UN�M~G�4����_�K�ȍ�[����*�xʅT����f���9o���i��ٝXL�0`�tZ>�PD0�������n~�=�_�?zU�/�e�'�πv-���Tg_O�Gg�Gu�����Y~J@XG��$ȥ#1���u��%�x\X�׍@�mK#����u��0��"�:��㜑��^���$�C-#���!]�A�����8&¯�	X��֡d$���]�h������ŦV�D\��kt�ݏQg��R��۞7[��y�
P�U7������:�6y!�e��	�:�����ח��_2K�|�xe2^VK�I�*����	h[�������XY�0����'�K��|v���h�z�/ w���:�w�O8	#q���n=óY��u�J��Q�
�������_o�9��>�����e��p��7�r��^��ͤ�!:�%P��*���kc3!�� ��dg�OC���Q�	�ˢ���8�<�k��{�p_o�ϖ@7j�3RCXpe�|?zN|pg��uC#ـ���Uc X�����o��WY�~�7���f�b��� ���Oߩ�����Ώ8jU<E��V�v��,���k�#�����ZUsy\�@'O�6����r)`��%�ʆ�h���CT7�d`RhI�/nzñ~�J�t�ui�LK��W�F�-�We�a\�:_��[�Fp�t U�Bd)�U鑞�ǘ�p6<R1��}>�G�S;�x�{n�����<����f�8vP��7��4�uӐ��Oh���`x�ԉk^ڃ����c#�1�C�ݧ?V����a�f~]i��!5a���6�� ��ۊ#�\ptł�F�u�%z����ˆUs�w�3���'�_���0���޻ea���\��|�|��W�'��l6��##�^�B��6)ލ�1{/�Q]�n�|K�*�Z����1�i��-��������,Dpo��)�`Uϼ��	�f��n��gCb��A�3p"�J#���#-��9v�Q	��d�/KoӲ�"dX�V�_��Sif�z��@�M��
��Q��0�@&p�s.�"�^�o�p���#��|��i {/�H�@��:��J�p�xY��0����=�/�Q�q�?��Xr.�kp�L���)Pv�C_���D"�p�c&~�R5h�v��������ϴH��}��T$��%�qX�W���\�?����=3�֗%�$�
��u��"J��1ն�?�;4v� �����p�F��wlw���FA��b�9��
Li��@��2�T~�M���1�M>W�:�3�v��O@��z6�\/�C�H��)�w��^���G�������Y*9�ɣ���7?�X�%�p{(��^����&]!J��Gf1��w�%�_)���r���K�d;�2*N��{Ձ�$x�i��Vw� ���p��~Uk!�k��O�%�8\"ot����.S���b� ���6�-'1qE���i��tߤ��b\�� ���絭��ǉ����(����#��O
�� ��h7��B�
ZҝĴv[Ў��&��	�,�v���hYH��# ���J���|I��t�R� �����#������nKc�Fmr'`U|%�d�PX+H� �+Ɨ�e��L��t���dl�L�4uQvw� nEv΄
��/�	.��s}�g>Y�;�nΞ�A9��p�ji�[(��	�q`�̊ЙZ�� �^2^��!���&UV<�21�b�̀z�摚9Zf�ж�c4��IQ��|x��B�f��9���Y��)j�p�}�"mz�]Q��pMA�C}0�z�'��X*�7妥h�?��
}}���$�{��c��YQ��cr��Nn�Fz/�C�AFʍk�����hFm��c���ܫ�$�A��}��\�4;;��}s�\�P�� �iHW6Je��fJ���4}��̮nc	�ӇѬ��-��^msz�P!��x�|�w�5��H�������B�	Mf�AɘU�9��7!��8���JY����d�Ww�7-1Ђ��o�]G.�V|����I	�br��nMSC�����S�g��Y�y#֐`���p>�W�b���g2I��z���Ě�����g�ԨÜy�We�5g˕VjO}V�FM�E	�:\3É������a��m��u0�G�L���_�01;�����j��C�5��._�5�"���en?����IQN4f�bi�9p��<�6�/w����6�잗,1������)�J��฀_�lN�E�@�	��� �5�_�7��uz�5y ��s6=uP��yX!h@y�gb�������:?�kr�$J�W��jC��~�^W�s��<�U��q��a	\V<h�w�8�7 <~�p�R�I����[?AS�0�X��`ye��W�p��N9�La��$:�V[�������������2|e��'NQ��j3w�3䔰�����i�r!A�,������%�
��@D�/(ӷ]��N�(B;yv�ZB�]� %�2�+�u�D�X�؎@�(��������Ü��l�L*��k��/e��R���[�6�~y�̷�ޕL��bc��7���i^�d�)�n��q!��x���缘Ғ���t���f?��9_W��-9o>�&_ܲIGX+�Ñ���+qyr-���h/į�"�Q����L�l�e#&2��s�8[��Q&���Xk���C� ���)-KGl��v�,�U) ��Y;9[6�� D���}5����}�S'�	rh��{q��H����9%0	v�H7��:�Z������i{ d�6EU�n�>��y%,� �T�wn|x�:��l(�_�|7����h��:�'t�䵍;bwA�Ү��n�%�5;ý0��G�"��{@��^���Ա?F���oC#C�Ǖy���q>����EBd�-ߌ�rw@ì�ߝ�{ShU���Η�y驸ݬ��|||"|��3D��UqV�W�ǋ7n%r��I�X@�myu����l|�5�Ԏ��}�Z�|�f���`�o�H�dο����_kl����)�ܠ�&��[6�6?�]����d��RB/���o�je/�,
,΃A�H>aT�����"��p�G@��ټc���u�����LS���1F�i�=~2.����	�����h��ƺ���z"�i��˶����Z�O�b9�M��O:HW"*Ạ����rt�;5< ��l�c�F�0�<�G�O+?��m�O��J�I. VI��N� �����!�٪c���/Tl��;Q(_Wǳ��lХ�p#і���#�I�[�d�#\o�༴�	�(���]��P�b�k)\�\m��[`�v����qpN5�ϟ��#�C*:D:�vp�,^r,C�Kɺ�w��������	���_?��G"�>�F��~�+��W���L{�N8�LR��LR)�!6��.T7"�92R�o��/V0->FF����x���'�NjK/��-�C�b���ux��/s�r�Bl��˜��smVTG=�ϙ(!p����S�ċ�2���"U�B����2����8DR{[���z:�J��p�I|��5�t<~�Z�N��i�F�e+ĺ#-� �/�jbѽY�❏�޿���TNwAg�T�	�p�����RT%�?h����tF]3�"X	�mk�H��x�&��3Q8ł��d�h�������[����?w�F�7o�z����S~.ȴ:s�]�D^zp�$O��Q��M�|��{���^��#��T�3�T��WKģ�~�5NutN�Q@O�y�7���Dܧx����G�X�0�ۍ+�8���c�ͷK���r�LIɻ�>?(W����Ox�
�������8���I��Y����:�X�5(�v4H�erǶ,���g,z����!{�I�)/�>��W=��Ҷ����-UH��D��G�V-�c���|��OIj���"���!���������܃�A��C.@�`TOC�#��kr�q|)��[d��$���θ��~:������eB�	����B2u�!�%��������<�@2D#���k�B;�L��_��hчtXLA�P�����(j��䒧S^�� 8����g��<��<�t�˴H�� "&��ь�$�KNx�? HQ���$�E-�IHS���j�k|_�����I�2�[>,
�ފe����p��/���m����J�{�c���=��@�z�:�Ϫ��W7RIv�Z�g�z}嬹ɏ��<4����W���s���޻݃~���(�:7�`KB]�N5��O���k�Y��@$pd�W����;]�Y��O��N�ա��[��jr(��x�Hѕ�{�M/.>����hʢ����EL-;z��SM[�L$�뒄��q��0�0���o 26?�5�TV�g6ڈd�tv��)2����	L�B>a2����
`F�}�$芯��ǜ��Y�o�V9w�ϳ���P�DK��F%�����-7G}>		}lb[�b��EnS}�9��pu��?]��u9�n5����X�2?���d��Vx�L�/�5����[9�@����ə��d����^�>,�޼H�e��><�H&����U�Kj�F!m9�:e�+V\�a���� X.=��%ʲL���ޣ��Ύ����xZys�&l4���ɮK8f��:�cWm�\ZnԊ	�I���pD�!!��!�ZA�����[���C�U"Aݘ(����fĨ�X��6|�xUZD�X�m�x0�#���?f�g��g��*�^1�Z���k1�J�S��@!}	s�2X"��`5�M.��yc�Gh@..|�i��W0_&���{b-� B�J�D;!"�[n؜7�ެ�{����;��}�E�r�����d��!����>pj/�x��?���vD��*.����k�	�����x
U��.�͞΃��V�W>z�G䕲'��
�=*���¾�*G��f�������c �ܰ�k�1�I�3��Uj�F&��*Ѓ 9xH��Ѩ�*�{�����y�m�<�ٌ���r�R�o��߲N�d��K�a`۰!o�7����Y�����7l||�f�f{��T�|�(W�bY�mvP�~ӂ�aلķ�A��c�'@�!��z7I�o��z�����ac~x�y ��-�BHk��,�w1(���0�q�?
-_�8�ʠQ��#4�g�f\Cx�% �+h��q �����6u���+w�V 9C�n>�+$V�(�\������AY��J����sS�7hRƧ|{�,LvD�Z��kl#� �%�7����%�V�:a����� ��|8�h�.�J��"tCjT�<1�Y�#����A���U�*��/F6|�(=��;cٙf����b���8(��g�n}��n	C9,}���p�g`����/Z�f��#jh�V��tm�M�c��	r�=9�-r�����2)=�����~cH�*Qj�*�Ά���Զ��,��|�����p:�	�@j��0�=u�}��x��2��.�;c�"��p��zdq��=
G�����%��;V�J%I��h���E���S��Nd)R۳�>#iw()u�4"%�g�r��u��ڇ�r(O�D<9\��1��Jn|�uxa6ע�J
��l���z0\.�_F��bó�QD�u>�1#8A��l��fT��,�V�k�tAQ����tp���;E����G�@���H�P�0$z('���_�����Rb��IE�ؿ^����H����O�"���^���D��RN���C�fB.�l��Z��VA��h�F|xs�S�яk{��S,ӗ�z1��&u�ݮ������<$T��_��L	}?)�v�RΙ�I ���g���,ul�e��C�TA��M���m�ɓ�qt�Lu]aS2���&�X