��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jåا{�\�u�?߷�dn@6�zf��r������;���:B���k/Ï�K7���)��0`��]�P@��BH�kCgT8Iڋ<G�FO]:|��:	(����v�`XH���r�	�e�L[��ga�Yc�#�Z�5a@w�����=ٍ��n��	�+>=p���9�������~N�k��_f�x Nk'�X�!9���-��]�.�����^�׺@�/�P(�)����Y��$��Ź�t�g��+S-��R��(����K4��f�������x��	G:J e=�u:7�~��[����Vh�N"���ܲ�Iw���#GFE�c�m��|~
~�Ǳ<�jCɈH��f�͛p�A�	gN,�1t����Z��5�H7���
�8�u�f"V���ce����1�S=�#����U��.���/��iptO�!�7�E�e��ly�.����*�Q���6�u��Z*�fפ(�`�������*I f�k?�����L�Mz���qL�&�Py��X����z�����z�f��2-`��͏	b����m���k��έ�~�R�����A��uFas
Y�]�sA���]q�6Vp@�z�^�Χ7XK=�{~z��N��"NB/I��6�YVѱ_IȈ�ٵu#=�Ԣ�$��v,�����]� B��ܗw�C��O�Ÿ���_=>L&������"n	@-mmJj��r\9)�d�r����N�A��rO�d�5�پg���êX�xԭµ@j���3��(H�mvn,�+G�8�}rt��s@o{ZL}����h��Ao������:%��y�J�f��Xy�.���1K���5}<j���|>ĵhr��R?Z���m���D�{����m��Mw{E�SFw�y�&'F��!����]���e��-�Cc���|��Tl�Z�s��\�2!�.��[M�+�h#�L��"�2�2��#B��%��]ȷ��Q��o f��H�f6>,kt��T}�������# �J[��W3���|^�a����� ћ�Њ�`s�%a�"���T]KQ��@YKGُLnO_��߲z�~I�g@�2?E���ؼ���ueS��-2$�C7;2wR[~��	د*N!>�i�8��gړ�5�ȷԷ��Pr��睉�Oy���U��c`����_7ax���XV ;���JG`ۄ�g�d��\>��3��j�?B�s
�V,�}���E��x�m���<�f�3��ت�[�� �1D��M�d������߃��H}�%�h5�x4��I�� �õ�b%�7^Λ�zn;B��Ͳ���V9/�&A5�	+6_'�����=+4�Sg�K��~�mB�O[����$@�9J��\�}���2VU�q��NG}�E�{O~�,��� ra�A���/�v>�RX?��߂����](e���ᖩ$��)�,����tW����#ቈpIZX�N��kW�<�D���fa�u~�yY�rp盹s$?�Iщ3 AK����� _��=���q+��j8�u6k�ȰV�]��.2�ܪ���k|G���lj !���3]�Ք�oK"�j@,L�N-k��%	!#�u�����7f�,��E�a�F����_��,��:x�"������	D�諻��nvM>�7:_
q+�.�U��~MI7t��&>��`J���b��Y�l�/��	��"�,8D(7^w���0�73��'��S kEK��0[>L�}�����NB=b� �@����,��I%ޚ��YN� �LՐ�o.�����$�P�o��%���k�-�S�>�Ђz洧y�����j�Z#qJ�����MOќnFr��̿^W���m4+QoI�}�Vh ���b�ٟ/��~e�Rj�� �-[4]s7�N��<#5l����i�l���Q�5n�����J ��0pm��	xd�fIF��U���G��-�)!�^1�j�Ԇ��.Ɛ�S���1�b+:�\��Fz�bT��)�<��#���� �o,�Bk]~�t���q��D��tP��Cd��7�}��,�Z�:�NE
`���J����Ժ�޻�{��Ւ��)ś�AJw�`(V�9[��OPg����P�6yv�j�s�s�����\�&��|׾�X #��r�p��sk��+ewEeg���θX� �N�5syѴF�\`�;||��>���c�p����!&��'��4[Qn�9�۷z���J�L����&(B:�������A`��?$�L���~��Ƨ�_ň8�S���D���4���8�������}��`$����%L�>
��{ļ� ��S%�/�y��|�'6�y�]�"�u�����P.�?�d4w�~�Z� �[f�j��j��K�>��\_e렲	���vܹ��:��(��tC� cut=���Y�2��^���#�r&w�8�Ogp��S��#ʨ��}p7�T�!+����-��@dlT�-&ќ@�Befz�˽��ܸ� Y����y�:�h5v��,����2��elq{z��LC�������ȃ|��׀{�oU3ZE坙Vi$`\�[P���)m�-ɭ5n�gN��0�ly�]�W�?D)%.}W�G�9���R��%�bK�Y૗�\��z�@ne[�!�o?�TS�SO��
7C�S�0��`ɉN����<��è;~1�}�Ԕ��燔+P,�2Ex�_���|�a ����O߻��C�]�`����p����	�8&��Eo��΄���M�j�~�
� �\��4�Y�>�֬R� t��u��؈V�B��U��\,݇�&$�4�Jzeu\�<�Q��f{Q��ђ!�u֗H���d�Vy������a+����^�?yp�x$#l�6���Ғ㫟��Gn�Z�:'^��Ռ���uUd�R���2".퇎���UZe�u�Y 8	u�֣�q5���"��z�!?X��tI��>��Ә�B��H �L��R�f+��?��&=� ^���UUUO�W�>tㆢԲ;9��`4d韰���4Ú�z�ie�{��ꨍ�	� W=xUd��nة󅢬�]l�jN|"�0�DF�F��@,o*�Ⓘ������/��־�Ng p��Z$ZO��_��%&������Z���b���Qz����ڞ{�����
┅�R�:;m�J]\�Ϡ��b,��O8UڥI_�,?��>���^�SP���qJʐT�(5��||�&����롿�S�t9\��AF�zq;��窺��r���I��E�c�AAȇpC`E�;�b�ּ�7B��[W�xǊ�'GROeFdĵ��Gð���m��;^Q�w4[u�:�y���c�(�%��h���q��tp�u� H漈�:�W8&,���E�?�fO^���s����������i�����i`�n�&c��B(tpw
g���ٞ��k͑����&5���)�e�J��"*�go���FgX65N�#��1֜Q���!�ޫN�z0�Re"�gq
�A���u����N5��1N�Ȣ��+�o�ݔ�TM�u�+�:���
�6�*���T�C��W�.U�]Jtϰ����3�#���y�oJ�����IR���CY L�~xK�K#�	o�r��A��8+Cs���NV�,�N�P�f��}��ñ[�u�x�&�2;�k=��+�}T�3��`�A��;��Uy���K�8��Uͅz\�����!\��������ģ{�a0���k ׏r�Q�s#I�>��a�E�$�)x�AR�m�$N;l�Ta��	�Ikb�C�h��k����R�N��S*��ڰ�6����g�y-R|MJ!Pf��Y����6��nW�AB�f<��?��p�Ea8��#i.��Ќi�,���*�S�;vh�hik�	k�Խ����Y�>�t����8b�y��UJs��[[��J 4�3��Ġ����Zx�(�g��x�4�ꦮ,�7����4����mJ�/�<�T���O�9$���zV4��!{�}8]>_�:�B��^�ff�q�ֽz���ׅ�oܮU�1��� �8 i�W��oH_S��6h7O#}
J��ޔ�@<<��TGq>�q�z���(Q��
^�;1�	�ˑ��yJ�HF�Ʋ�'h縨a�ui1�K�4�0�b�տ�0@�t�"+S��U!�m�;�Ͻt <���{'Ц>@��ő(�k(@V��є/�=\"�b�%�!o-%��MsIs�2�{��(X����U!!ã����S�'��h�m��>Kg`�?���V2ɲ��>�%���}��2���dː�k,�_�h��7�Wy��e��Q�%�	��"'�Iq�4eL[f=�}��7u%ZH��y�v*��;7i���&��2z�@����7]ߤ�Mz�J�4:�(?��ID$@+k�=>Kl0�w� ���oKPK��؊��]ɉ�2n$�����C�6Xѽg��Oہ��;��/�A@�JbU#��4�;0&s1!nIj��.��p��汦�}F�g���]wt��N��̈́R�m�'	R���ƥ�s���bK�'*����o�6'�D;��.�Fe�v�D�1a�j��~��pMh4�Ǭ8�'ťҌ�~�f�a��%�o�:��Lk$��clSd�k���bs�����=+�=z`��~��P�Fi�B�,�s;!��N�߸� P�ɨ����R|L�����a�f ���dR�D0�.��ɾ|��x�u��=Z7��{p�[2�#3�mY�\ퟚj/�T��i�.N6[�A�L���eOh��eų��/ϝ�k����U@Ke�n�~*&�j�o��?��v�(a�SdU�����wL��b��k��k8V姄�K#�4��T�E'sR�~��*5kO��o@�~=mz҈V��Y��+�q&�|��Ɂ��ߏ��$'��J#��&=0�(q�N�(���R%-�3��N��q���
�����Y���m�(���x�9�8���G�,L�i����ڜ�+6�לk�f���#������I$(Z.K��&��Dr��sNI~���u D��J���:��V{.�;�:���K-:�)����ErZ������	�F2�6�R2�u�%b�d(.�rp�l]��r�F�)���?��)	�`f���u0���4N�XG��W�����\Y�.m��3@���6D`a�&Cƶ�ul}����:���� T=M����b�@�i����c������0!�^��<�@�����r�������ɾ���QF%��62� Qs�n>uE�o�!tW�8ҏ.<�4"b-s>`�2���gרJ�l� l��j��q���Q�XӍ�eg;;,��l����c4d�cmJ��V�(僇��r�ˏw�zϸ-2�02��O�!ݏ ��)�Mta��~æ0A��bV�����w�яByy�(�偠�[u�F��WUY�.e�|Ѩ��I������xD�Z��3{�泄K2�zq�hz�BE(��D\q-��G,�
:�����8�����v��*�J�Jztʯf���.�T����@7���uc�ˉL�h�[ٰۘ�l�����qC?(>D�6�{��2+yX�L\��7�D	����
@��Q�����O��K���Vƞ�c���&�)��c�OP��r�Q�G`�]��������iс�(Y�ᇕn��}{"΍Š��_RQo��zYA����l�ܘn�鮄T���z	{���0��"V��ug�I]FI�!�����4TVͣ'ĔX�A������9ۮ�^�����kl��G��z�+Eu����؃F�����Y�&�d��N���&9�	���?JF�44�wy��*eXr"�:�:{���v/k�-H4:���s�/!��M|�e���X����s�2�#<��<���7@�8��^잏-V�� "����xA��i|�B��E:"�s���i�VCY' G��a�צ��?�4�bZ����q�A�"�ɾa6j?'1m����c���ܚ�$���#�FTW�nJ��L��_��jʷ~�/�3|��6^A�&�>'�l Rs��5:��]���ydK�q���p�I�J$�|��O�!��e-�`�J*���	���~��o��.q��qw������T%��\2��32;d'�x��ڀ�Q?�.���8k����Bd�@�����$�\}D����&�-	y���"����Ť�3e^�cO�|��:�XPߺ��>Aj�����e�y5Qa�3"�6�u��� �EoM�_���G��=�4O�
�-5b��߯ql����|�`�-�)QJiT�y�@:(�hV)��2��c�x��(������{���kA�\ҭ:mJ� �L�pWZ�>( WK����8F��M�y�&�g)��+0����	o�Ӊ~3w8���pr�>�&$�Vٓ4� 5�����>�+!��,�e��^��wO�xI��������W�+_�:�d��~p�'�����6 �O�p���t�/�zP;�8�}ջ�c��>�U(�&'i܈Ie#�h�^ǂ���.�
�$L�ʰ�g���]��E��$���G�| {���	+#�� �o�D&!HRa��B��:��#��1�2�~��l��òJ��+��/�q&%���7g}���:4w;���α��0�Q�x�2C�](�y�C�bB����	ӻ"	��J;�]�(�7	J��s����W�u�,��W|�Ѹ�?z��F�E{cpG�AwYM�yX��c�v@>�F#pNf���O><z9��;�w�v2��ٮ�ntj�{�p8�8w#���vp�>F����Q=�]{�
�JN�:x�d��P�Bv���֨3���L��^����wgT�2PD��Ҏ���bAɴ�`�~��Q���7�����B�`���C�������#�Q��8r��<xG�ݢ8�e�r�6%:�������$���'�&Gƻ�m���)��[%��chEw�[�o�@^�����i?A�&��{�s�`�$������:�X��l@"��!�p;3U��LW�f0���i)���N�S��5up��S	��h��b�;lI6fV�0��ɐy�Fl|%�c�NZ�ᮇ���|Lס��-�����l���T㹰&��r�B��('B���I�C ���91���J������r	�����|4~�ߝ&B-���}�LeR�˾�tf&�/�/=iڲ
c�
.��X�8a�O��8�ƫ��x�7�����Y�EugW(b��.�z7�n���bc{���� ��Q!��Ұ�Wl�+2E7t�MS���c�_�-M�KKS� 	�׬�>����q�ɣS�)r�o�hi�{�Al���g�@����F.t����t{�78,��=9�)��'�Wc��
.���{���ϵ�-���bg��>�肖��NI��1|�lU1Y��yN��~����`f2���͘gߛ�!���=m��f{b��E7�n�!���狓��;_�B��	�(Rփ�6c��X���O��j%ϫ )�-�����a�0g������[���s�p#R�4����f
���ߝ]R)���z+?�'{D<��}�$����&��+����0{�ls�;>`��=7b|���w?�1TD����;I�^ϯ_$i{�F���b3�x�X{.�����Ъ���9�.��"�����5��6�xrI"M�u�+���u̷�T)��[M5J�.�}�ȴ�^e�T���_"*��`�[�J��V�+�f:��7�_�µs���ocF���C� ���⯢V=������|&`nP�JsR��u�s�� O�i�'Ѩ��`�d��f[��W ��8u��H+��/������`5�ӗ�&Y��xȷ����1���)����<��*�8~���Ia5{�m�%��s���.�f_��+k�Q�6��/�k��{x0#c�n1١�c�[�$�1��w�P�PJ�{���b��SԫY&��0��[�&
��*�7�oTGvJ��[��N �G?��-q^�rN�]l=2N�B�3���J������^��)�'ygv5T�Mߌ�W�>�g���Ε�G>�m�9�+��P����K;>�L\Mo%Aa_k��tشZ�*�o���qܙ�v��EW�je5F�N�h�M9*g�.]�RV8���:Cu�;?���"��U4��j��͙�X�嗧�f,f��􇮪�����ӳ��ٹXd`�5 �����Cc폑��pq�˛�����Tkx�oC6�O\'��W�Pe����|�p�ZT<Nt����,ާC��'/����:��uϕ��d��U=��Hv�;�E�ë�7�PW[pʓ���l]t1��GfI%?�r_�`�����#�������2�A|��Ö�2�̜��V�v57I<�fw�^��d��W���M��Oǚ)��fT�`�w w���<����xu��=Sa��G���	ī�VtL���M�Ib��iaJ�][� ՒA;�|-���ɴ�o�;Ҿ ��f�q���cl����8gW�E.c-y`�K�DR�h�1��bfO�w[�T�:<���n �Q��s��Z$�v�$w�	jl�9������&na�@؞f��طqy��Z�	�9�nD�'M��^q�v��CIR�u�"�o�O=�Kg���U�1`6�����;ʎҴ<93����z�}���|��8�%����TBjJ# �Q��y�߳��8���MUڈEІ���V1�䋄H΅%
,�v��*f���s$��P��o��+�'N�l{� 3�L���Ķ�e��t��o����|]��b\�W�D�Z��$�@���vg٫$8������Y11�D&���G��Lk:ڒ�c��ؤFH�:��C$�ߑpU�������	���Y<�G�Z3��.�9Ŧ�X�Ic�