��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� ��5���5j jQ+���t��-�/����u��̩�Xc��R>G��$b�xA�Fn�z�F�X�Ӊ��q	U�z�qG��f;���,-vl��� 'J:>�V�	��0�7"�%�˝էo%���7J(]�7(MGw�rL�R���<c{��y�y$+{���k��6J?����ye�@��\��q3�!6���J�9�I�ʋ����K�e��t�f(��oǎqz':ݶ32/�.��.N�
s)��9�<�2�B�	>?�����V���c�Kz6]��0;YTHܧp��VS���J�0�L���<�0�q�j��`��Ѕn��-޾�Q7�z��׿�<SP_b�
teuϋ$y}�U��4h!���'N����F*9� z�[�����B�'6$���111��>x/�mD����_�X�5"���B��h�`�I"+F�8 3��R�f����<+:�5����]�-T̖�ߒ"���|�S����'l��]{�`!�к���7��*֨h��3��9v�w�'F��	�;����=6E�EfW"�UB�t ����Å��KKY��Q�&�5�c�Dv��7X��񋕲	+y��h�< a�D��Y?/��Mio��dX��vz��{[�BJ��?qq�:۟�hF���X<�:��/��|�5�9�_�'��0H#��丯����Ҭ���@z��JwHy���F ;��ʻ��ÛV���Q���>��{y5H����z;���Ǳ-�a��!��m�V��Q�J:p% ��[}���*�ֵr�P��ݯD�/�Q���>���ʜąïI�MH��V�"�HMf��$�o��c�AUl��K^�!�p96;�����Y"���p���_�a^!�M-'W�[�r���pU�w�i�)G��mr���l�����Ə�?��X8a�o$�P��L���'���_�H�4�>p���-�ޛ����Xyw'�(�ha���7��j�4��<W\���d��-Z����8d�Cb�Ru�'xr/�������h��E�DF��C�����N���paS܇�H觮��bcz���a��Pa��<�J�W�XM"!~�{�)Ͷ�(�T�X��rȃG��s�q?Ǥ~���1��������B���ޚE%J	Wx���=zI�6�����[.:�L0�T�(�g(�Q����*c7��Kz<"t��,��ʚ���k�|�i�Pޚ�餎t�=��|�����XG☺m�~��vZ���UV!�=��Ϳɐ�複�N08�Rʹ�N:uj3񋆿�#hH��b<Y��pn��:���(��x�R��t�)�(3�0�V�h�-	�?r�K��-��F#d�YD���p TyM����\�x*��9q*��1D�w�xƾ�N���)������
w�M<ɰZ��uGA����^:1��ɧ� ji�=8�;�s�p� �1���/D��D�z�;�*�T�KNN?ʛRrR�D�R���Y��&�|ŧ��N�m��\�Vd�/��37���*���8���^����@%y���=d�ǋ�)���]�o�>����F3����]e9\P�8�F�t[q���l�[F�'�x*�`�q���t4j �j~O�?��Oo[�{6}.������M*��oU~Z����Lhώ�߹�GUy�[��:����*����SC�Ѣ_�LN|�����;����t��%<6��z^b��6ѩ�8���*��:��FW"������Jc��'��c�^�&;+�nv=��H��o�{y9��}��Ӷwl���T�7f,G �������9����覫jS�{�Bi���`,>W�WZ�@���2���c�A�fC�~O��~q#���b|�ŀ�A�#�v�MH�aS#x�fI��}Yy
^]þK�b�I'�;���\pq�
9w���hI�|]�՜��U���j|P!�z��������jJ񏩁�NNM�(VS�r��¾����<�]�NhiZfX��x�&t�~���~�����B��Od}=1�_'��I�/i\"��W�����o��IR˄�9NDN�0T����p+S�rye���a�^m�:�o�0,��퇹<��a��zMP��G��'51W�G�MS��\%��d�h�gs�/�"�Ώa]���[ �n���L�oϒ�\@w��z��U6Y }��O��A�쩤	 /IY=�Έgy��J&`E�n��^�d5�0���Wa#�C�ɰY7$��4��	i��W"[�&[	n[4/4n-3�u�/��'g�G�K�4c�׀0o���1'U���v�9�U�tTX�A�!�?�I8��1x�t����mV�����:'�]͗oH����M��nG�wY�\�M�O���"�_:Z=�,�~����T�T;YЈ~����S��,}p2�OlR*�������N�o�C�NC���3�1��ӑs@�}��F%<�#CH)�����E�K^\�h����ׁ4�d;���n/ګ��c$1:��k���iM���Kz��?5�!������}Ru4��F��K�
� uٰ��]�i����Sϰ�n~[5�s�n���4��;�!��X���s����}j�t���r�4}}����K޲y�Z�ᲜZU��,��~�ʾ�ǜ�Gģ�[�\8��C�)��_|���E+�]�ۓ3w�l{JO%X���Mqw�mr����g#Nz�C&_I��Y��+\}|-K���!)�����>�����=��:g�	fC/��Km�Vz��ee$�~�:�c�k���2k� �@ˬ�"��٧de�y�$.W\J�D$C�1g�W{$���'ۼn�(-;4	_-�c���./'M��J#��I��_~yzƉE��o�Q%�/�IY]@R_�e�%��v�=@++����f�$�u�R�BM��0�H�Z=��P�[�w��,�-����"�/dO�KsM�O���HbF����\�����a��GmgY+�������#���͜�RKCb��ztv���AkTW� ����?�o�TiƤ�du쁗�5�����d3�39ep�ǯo-��X
�|Gg{t���ir�ƕ�Q�Z����S�h�Mu-�l�[\���h���P�[��f�9qyO��
 �W?0*6�Ԛk��k��چ���i��{t@#l3[<�+����Fq�\pq�:��Iɋ�O��?�ڼ�G�L1�r����S�H�ݱE~����F7Ӏ�_���,��~�bH��D!�����r�W��u언���8ЛW�,=��By��=�8�.J����e��@
�4� XyEq�w�w#��ɲ�p��8�G벁�29Φ�xG'�% z/��T�?�$qY�"��߻��!6Ť�C>2 @��p�=3��c5����y�fNJ)�۫��(E &�ڲ����P��.r�h��mg��kS�VNhK��dm7����͝��Y�_)��s��t�m��q��Nm��EXh�����x����R�D�� ^�'�Oa���@wo�Z���Q.�*3�$�=D�ǓV3/�E��ֽ,_�m��o�KmQ��`'�ъ��r�J�9pu�}�q+��}�����R?L
�J��Y�(C5���,Ȩji`��ǉ1L\>!0�m�k�}{�0 u�hH�m��셝�>��IJ���������ei-��ܯ@�ۗ��� J#y�^A�5��-�N9��.ԿJ�-��P�30ܽ3�rM������푥{�rY�=+��n��̞%��n��gGQ��=A\�㱸~s�>lj�6x=�p���S��1b�#��BE�%&Z5ۤ�D7=�m��+1Gt^P�W��[�2�ܴ6��PD�eb����QT�7��9V��_�J�bA��|�S�I���a0@�5��"n�-f�3�������ՒX
�f�����VJE%���{|Ws�pka#�����9�`Q�Ǘ�\Ԫ�r!5�b���#��RF:˹�=w;�kb��;���TDD�&+�/�lS
<�p�>��{tՓRKD�����'����?���}Q`����-�:��R�@rW�uե�M�+�*�DX�!;`T�u-d�sTwWƂ���(O���Y���Y%�%p�m�w;����%�Y"���gtbG -ٓg7-��.�Ӹ�<5b�#��.�Z���+��2܆*)U��b��_\I�j��{�`���O���u�v�O��p���>�9��'^7�:��*�