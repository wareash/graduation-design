��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e����d���f{��@����S��>���4{��ת�AO�Q{���v2�������n�yK��l6���z�X13nדF�1K�\��فH�<���Q)�[ϣn̿Ԁu}Z?��<V�Ժ�	����&g��΅c]��$�>�K76 �o�:�5m3�?rG�O����0
��*��`V �^���I-�C��$�w�	L�z�*�v׳O�!�.k��${�S[���P�+��'<�af?�g��D8��Y�8�jP�N�cJ1?]� �$Xt�^4=Fn��L���j�e.^P�<p8[�+`�Ű�qQ��nh���#`�U ��$kN�� P I�՟�U�h痄.���w���@���:'�w�(�(%߆�2q,�%D���-��S�mʭ���ף�G��|�s#���������`�\o�v=� �07����M�fhtLs2(�)G��?n���B��SU�0��gm�Z;l���8���I-��Ă�l���j8}0rC��E.�(���WCb��%ɩB DD��$�ga�P'�q|�I��㇭y�[��&(L�>{Pb�f��p�.�Sx����iK�"�q��쟱k˓z�vs|$�S�'�7g�T�p��1>ͮ.�!z���Q��k�>'��x��]���zY^�{�f�0қ�#��-��=��5�v�k>�ϫ��]{�9�d��.���ూ|S>q�6�����ՃU�W7���Ȼ��oh���b���a.{��_�Ix��£�Υ�N[��|m���w�����M�� %��	�������QT����BIx8T-�SU% �����ڻ�3!-�!]��e���
zdm92�8&�@`�S i����EVG?Ȅm��%�ϪB_�T�E�/���M�-8~�����,LHx�d���xr5�,��ѩT�Q{��3X<F"ԔGJ�b�	٭��1��Q�㗍���J1�E?x��[`�d$��vjTTA�Ӝ�>5aoM�d�U� ��.�� �0ng�U�e�#�V%d���C\����2GW����ǩU'�c��$�,��sVZb�Q^n�e�El0H�� ���������D����������#���� ���m����������6�u*�w�s����V.���C��C7�Y�q��Zj�޾�sL��z��&Z��;,�b�_�!M���K��Y��ES�n���ǐ�D]c�~NJJ��I��'�=ի����ax�;�������_F��?c�G�X�f��8й�hg��,�˲-IW>���nf �6:e>�z�����P�N֮!H��i_S*k�'�i�O��w���ȘQ�I�^e$d���2���E9#~�\�[]U������;�Ʒ ��/��`�r(4k�5���$XV�K' ���`^-^��U�!���aJO0H�c�?�"��&ll�DV�E1�r���0�|	m�B�a� -d	���F�� ��qg
rA�Ήzس^jn&����g\H�?�9$bP�Z?�i��PDN,�K�wxRw�ƓP����Zd����C'�P��4i"қ~�{z�T^_�=<��`ȩ��tc���ݣ1\AA�i@@�������uE�ރ�Y4*�C=Io�fJ]\���B��×�d�FU4�8�7of���̏
?�ꕢiN��hڐ�6S >�5qcc�c������v%Y9�X���X,��z�C���)����Y\��<f����!�'��I�w��9"=a����?�]E�t���{��\�o0�,D5���aq��o�1=�+y�ԙ��D�-��D�fP��%��ͽvG��WE�`�����ya�!� l�c��n��6�,L~3;����s\æh]�����y���y�y��U�A�7��f�F�0�o5Ӗ� fκ�ҝ�3w��O��џٱ���^��Ax¨ҳ��;��}���I�Vb{s	=+Ҍ�T#Po���+�8�}��~�l��D�ӓ����7�������@������Q�uc�ܶǤTp�|���O��ZK?0����\�/ڟ�gz(*��ZQž]r��qX2X�kJ�����;xTQ�@{��u4�� '�=z/��<N|H#������8�Mڻ� �^\J)f�ކ��N���]`��ׯ��ܾ9u�5杳�YԾIFF�p�}����{�z��)]��}�;�Xh��f27�ہ�|)�0�9i�����P���`�N^lӇ׷���Ec:B�8f6²ϓ��7�+�O�3O|_ݐ !��A�h�P�����J#
e=2�cA��3i��	�	��7�u_���X�����	�^��~��n�?�,.�m
s�t,0�<zwT���O��q���}1�]�U.�:�� 2��	��T���{-�N��%����P*N���B�Xn�'�Іia
�V�e�S���J��U�B����/&MM�CJ�՟Cg�k����M�Ċ��5�2H;>��������)9M��!=�X4�����tG�0(G2��Q���[K���M��%��u�pj�kS�g{��P�mU߰����4�@W/�@ȹМCئ�׆s�q͂6�N�ޮ�	H�A)��77Wǟ2�>�vn�I�В���=m��]��Ev�a�sX"-)�ůVX�+��4�c�!�&���Gyeu4�Z�������)��g�M@�"\W��=�/���
l��%̯@�B[:�(l�o�?�:v���o��*�l�<��׌Y�
�'v]&\�7+-�&��Jf��}a���w�s)�t��s���+�]0�^>ɿG?aA���@��%m�a�u��c)�f	�.9W�>��E���a����v!�w����+�3���]ӯ�����%G��$���F����|q�\�rl袇n����??��l�۸��g�����/0����{Y� �)�+6���0�q�ǽ�~��xT8$ġ���ǲ�6f� NTUhwi����r9W�­�Xv��RC)͞+��b�;�v�ON��Vx��� 4p^O�����꒣��"c�Nd�26��A������Ğ^�Z�:���ƗM�ʡ��Ϸ[9h�^�X���<��[�D4[aP�BeqӰ ��H.O�d����K1��B��F|��.1,s��P�f+�zM���'�R'#>Wu���j	���zؑ��[S_r
��AߘK�+<�t���f��)�t�nWb�����%,h�u��:/�dx��6�q�2Aˍ�z����U
6Q�2���o[Zؒ\�aǁ!�gy����A�I���`�:�{B.	әLϹMهAF�.�}iWΕ��J،tӆ_���
��c�D�.�HjƺX� fXO�p�Ɇ�9%�!��R�Q7(�v�[$�<�.�w�����do![q͹kk�V�H%��Tƅ��ܘe�#qg��%�cZ���z��$Gd��+�'3cZ�r� A@
�m�8����c��*�r���
潙ʡ�>y�{������_l!�Hk�vHhʶ��a�i�iNsvT�+���D\�E�J�/�s�% ����0�8iw�xj�e�Bm�=52sC�σӾ�e�1��y�5���D[�$&h��J����	*�8�.ղNc��Z�(%�x?[WG�)=�7*�ב�R��a~�_�CP��.!)���������w��М�93@#o�	�ⶤI:b��g�e�?��{�VA�i<�ӵڝ�s�Gr9X+�L�e��_	�!��U�l�|-T�ҚlMfQ��p٤�=ӥ��$,��e�o�v&�Ap����B�r'T5;rϕ�0��-RS�{�i�,n���.�:!���]�D��?Ѷ�#]�'ߠ	�q%߇[�0 �e $	_��]<uc�>=�J�yh����s:h�Cm+���8;d��n���!X�ҟ)��{�~t�^�x ��J�Fk���$���f��Y�׋ �<��}�]w>V_���0�U�͟��^Lّ��w�:Q� �E� t����3[
�͕�߳rl}�c��&��o�t���-�f
�̌d.�>eP��A���B7�3V>��osm��ɯ��O�\��F�_��Vp͜#�JG��џ�3������v1��m��C���	���m�,���ɋ�Kϯ��0Ƨ�JerR�4�;���keW>�N6g����F٥�l5���[VْR��8p����Q�9��"��3?�ݙ�h,s��R&,-�P`��a	�h'��A�a-��ի}�c��J��|�oX7L�V*�72�5Oͬ`��1�~��7i])����u��`�ܛ��F�i��*%����"W��a͹L��_�Nj�e��?��۪�=BD��1R_�R�=����d%��X��0���P��qF& �m_�B��hih�L(����$�=�c�����r����5�vp�S�������L{���F!5�8��Ӊ�Y�ީg^�̴�4����Y�cy���a���Û f�?��u� �V6�HW���x8�8(��%��La`'�nOOI�/Ӑf�c4�p.;��i�	��!i��X]Jw���ǔ��>0;~K�0�W��?�]�9���}s<*,]>P�	���{
rj�qX�H�>>!X\Fq�m�s햤{H��ɥS��n��_u�Z�aq��c��J��7>�(xף��z�ekNf\~L@�dԻ�hr��0���rD���6�.��ş������	�Й��^!�gP��4g���g�M�����E�E?Z����B��4�3ܝEr'�w*������"��������Z�5vi��B~�))aW@�WϏ�)S���m��ll6Y��+� �hi�~��#�zz�j������NeOK��4c��T'�G6�_t�I��s���
�|'�aB��?�t9Q���}=����ɲ��tB��*H���S�8���M��6���$Z/znT�͎{�f��[�A��G�%�ʮ3з&��;Z�"r�&�z�8���)�[:#���]!��.(�� � }��c��>�b��<��夿����1Q͹Ȩ>=�o[jq϶8�%8��Sc��l��V�	����jh�7�̣���B1	�<	F�KCPb�r[��f��(j3��tf���-�E��P�k�Vʉ����>4���>]D�|�n���e�*K���GM�b���X`׫σ+Lq�R���!���ĀL;�qP�� l�3����/��b︱{�l�&W*�8Xh$k*���C���Q��\�颹v�K����*O]�%˩�� O���Lv�W�;��/��q�M��ɘKP>��"���@��ߢQ{R���6�oK}���9z�p!^ib�����وHN�im�٤��@PڸU��HR�qE��L}�w��<�B����+�S_�{<���.�}�+�jJ�W=ˤ�05�?ӛqna����d�ZU������Mr��p�X|�=[خ��������޾�ݞ�Lp^��,*y6G*�,ߗ3�f�v�*��
��k�Tӷ�v#ru#��Q�1��~!4	8ۮ�"��p K���Z8_��K<�e��%�/z���L)y=.ѹ��if��<�ۨ����0$-p���,�iLM�Q�#a,�מ�C�\��غd͍�d�`�k>8�щTK����	ͺ�B�=/�&ML<�.=K<t�f������݉�L0_����aO���\Ï~��`*
��.q�҈lr{�A�.|��e�꪿q��ru`���|j#(]��%w�J�i��-�Y��e\=r�(��4-�L�v�pY����"���J-P�_�"5�/�{&/}���py��i@�ڦ?WoE�0[���@��d�����oٶ�[� >C���q��L���T������	E�i�ҳa��Y����G��^UdI2��ǖ��np>�+����� ���7y �����9u��r�g��q�fdv�vN�:����T4�-�{���k��������I�����$���c�(~<�����J�#n�&ոJ�+�G�0`�"d���*ݡ��fύ�}'<֘��Tb:�E���&�pO��ci/��嚙��!���*�}_y���>�G(1�np����b
�J�<��H�z�.�#N�@T��ߘ�����w.�#m���%��eY�Q��c���畋�#�-^��T��=B���e+� v�lkGp�k��j!���IT���/8�!�,'a5�N�(Ҍ�T��':l�ȇy����MCE��L�f���	c� ֩�r��E�=��^	R�=�a�n�"Z�V>�5o�%S�(�KԞ�^�g�˄u��|��2V��xCꑬ2&aC{�>,���,,߶B|�~)���+�����C�#K��%G|�+ƈV1��j)vD(�=���:�9����a�Q�v�"�O������0��1�l�ȓST��K��Z�<�m���:���f[R��s3>7���!���	��͈����_&���Fp��Ẋ��_\Q��2T?�o�qV&
Q��:9]&S-�LA�K�.4;/�Z�}$u�Đme��
CS� ���=�%lk���7 Df9�=guC̃m�b(��x���31�i��F]��ʢ��K ܭ��w��nL�J3_�m>�h��+���A�:椤w��NB��o�EH*�b��[��e�n���I3��d���%��ܻ�v�~R����.���mf+s3p�kh0R�!���,��)�*���ī�r�nc�����*h6G1{�����:i���@�����ز���1]�ѱE�~ �]Xd�z���~���t�IC1𹪤ұ���מNǪ��-h��gS��pq��V+�I\8? �����Q��S�E�6���2(I��*�ʠ�Ǵ_���)�,�j0�K�R��u�U5a�t����i�tKw��j�D%���.|(�W
�c�L�%���d@�����a�$Z9�A�v�P��QgT�ķ�CX !���o��\3�>�-���=�(��������-y	O�vfP���-�!]�����b\���م2A�/�>�r�>|7��$4�P����&w ��鹬Tщ�ÿc�P���K���4�ݏ�ҳ��U�C��S�-U�A3=���E���`_� ã��F��x|�h���vP��';���g\m	'�7E����8=dL�㟥0Y����3S�yǦ	^��h����J�R�Wo�D��"��Y��`=z<Q�C�`���=Ѯ��@i7�DO붿�z�]�--E*N����NH8iߡ��S�ꜘk�����w���T���g<D�ѮZ��m����$��?��h*i��1
�<)�ni�fb�:Q��K��<�T ��\�u�	uJ�'[�z�P�t��|~,����_9�σH�{�CPH�T���xC	P/����������?�����B��d�R�'�<�Rbc��������_�b�']�~�T���s�1�O�S�O��N̩����X>�1!c=>�SrQ��y�#�2��{��DbG5���T�L:J3��8&{M�y� ���x�-ʹ]UMJ�u�����������}QP��9\�R����K��or����i�u���)�7�)D ;{`]�n��K�n[{�3�G	�F�A;��Yh�\G��ld����>�>>&BwS�]/��4� #�a�mSN�g�b�VEnGJ� W8T�������Ŏ�T0`��)	ӪA��ZQ��fV�s�P�T2;e�AhͿ�.�h�M�D�G�Î9���m�S;:홾鶪/ؤb#�i���`��W��@�egp�I\�u��pۋ�P�,+I�-�~ԭ�.�����@�#<=8��(E�����Pl�����raxR��WQX9�d'	����τ�]S�i�kPN�&�&��P�H�.)�i��v؅9
��24�X���a�!��@7 Lu�M���"x��Ő��O���i�7��ZO�:���C"���烩ឫpB�|U�^���mI~�
Zk��H�n�v��)���B1`>���7>S����[�� H����T_�O���_�eY�G�*� |V�F~�1��������eL�bR�B;/���rRz�[��M����xW;'�\&����$2�=����Dr��Yד�� ��xX�]b�_zt �����䈢]L�a�w�:E{ua��˭�e��`�o�"Ҳ�u8j@1g0G�C�Y��s='F�KT���� f+���'|�P_Jk�' �Vq_�a�&<	��:���.�i��RgG�O�r���W[G/�:hB���F��ZӞ��W]&ş�)h�'_�&w�I�O������Q��)��M����y����6��@Q<�߯��W\޷8/���p��!N��Q�:s��'�o��6�%�g-^(_�l��Ǐ�q�Z�`��-�`;�ۙz&+.��lӒڷ2����b/����IK �6�/F �֙����iӹX����ow|U����h������p_�y��Ɗ.�Dbڣ�<׵�Ƀ������I��q�,3�`?��IhAp+�g���Lg��f�؟d�q;��/�#����i٬��N=�~�|�!|d��&��T�q���EEw��c��ȣ,Jf,Oʔ�$.>���
�T������Ƹ�7*o�p����ٖŏ9uڭ�1�x�pL��_`Ȣv����&Z[���5y^�i�+� ͍
="����&�Eo�sS`��W��%:tf9���w:)B�Po�v�:�8n�/&���>�gX����%��Z}����-��K"ZU-i�e�����fmѽ�>�
bQߎ8\�n"1W̨���Y~K�����?H�Ov�!�t���Հ��Qi
�3�{��vI���}�gd�D��h�W��1gQP+[$=�y敠����i%
���	ʚ�/߂�����&��ʺ����%Ғ��y��k� �x/	���Ja�x[�b��"<P0�`$�@�"���T���5O��;�/S���7�&8�괈�o�7�P�f1ߑ�l�EOi�?ۜGޡ�^�)�#�4#������ٰ�,�
c���ezgR�1����G\�^�c���r�KBWse͉��z.v�Df��Pi�h��T����Y!�\y/����r��~3�?oT�Wc�k%��׾K<c&��(seN��yk�o1j!�@,A#�>iZ�`�\y=C��7D �1'rR��ޯ8]��KJpY��eo��{�so�� �C���g&�!�[�"؎|c�ٳ��М ��?"����!�of�������>j�:���`��.V�������x_�7��Î�yi+/��Y���9�����O��!,�8����_�y��yD$e�����l�6�V"+ �Qi��J_C�7�]��0H���05�B�Cu���+�҄�+��������>����o���Ĳ�Te��m�vG\�F;���`��C5���a�nѭp #����9��nC���b���:���~��&�3~�pg%@�1鋋���T	>���t3�Kɤ̙� A{��Q��IV�t�u5{�t��JeA/���FE���pj�ߤk�f�]��T[�99DN�Q��x�Ўn�^K�X؛�X��a6[?/����3٧�'�M����q�D�XrZ��J%$�q2���Lൟ��޻�־�m������d&^a�h�a�_Ŭ�q�r��[����9��5/�@O"y^�볱���X|H_�w<�s���|q��b�qk���Y�OT�E�2>����
��ޯL�َ?�p�E�z�o��fϓ��߱�����껋2[P�5T�4m���{�]�-�{�fVFj�Q���3�� !�Ye�\&
慚g�>���\��!!W)��#�$U��.��j��J#6I ��Z�?ŕm^Y*}�]�i`R[IǮ��uZ���f��L�F@�y�j�˓uuTf� ���R��m.��I�ǉ�!!��#QT��%��ݲ�D'�&s"&3���X[F�%��^�ֺ�/'F'��¨슁���qN~������!i,Ot���}��*1u,��#���M�%�Bd��+�U�d���2� B�����k_)|�G:�����Vg�����~���4m{d��l�������kꀠI�`8��%Q
[�{�@�����?�6���#�p�WHO�F-*,Te���{Ӭ�B���A�H���f���?�w�S� �Y,s��ޑK·~��������e�N�Z�!|�֟Y<����&�+���	�@��x�쌙(�(L�������!}?/P������ %g��e�+q6�f1t|%�����ˠ~߼�/'S퉋̀$*W�lo�& �&� �Y�\��&�@h��<������3�z�ݦY�s6�B1�`�K�����E����?�ӳ�B��+�R���մ��?0'���,ͪ��T$h)Y�"��k'�F%[�3���PrؐG��<4���/u��}^nTG���h\t���a�!�
�s�K^~��J������n���w�����F�H�ogl�^��Ap�\��i���,�=��A�����!x������S�	<M0�ƃ�4��P��y�a�����|8�f�!;k��n�s�lZL�0��\s�}�
7�?]O�����������k����SN���O��5y��"\otU�aֲ��G`s#i%R���L�k���|�"y��$����/��U��cpe׍/���p�]t����{�7�b���ώ�<��`�^T|�y��MYo�$[Fa�����y�$%q+eoi���l~4yY����ڲ�a����\EtS��0�'������s�� �B�Ɂ�ނ�$km �菮�g��g�����į�(	�4#A��6ǭ��x�;7 �O*I�թ����k�����cڅ��Z-Q-�r�)a$x=��#���.7vK�P2mmTr�����B(T�{���T��\�M��>�P�]4I`�!5���t�����{v�'=�ǱT����zVb
I�V㇥a�;�m�?��
���vY�sZ	'j�{4�h�_��m�����@���]�̈́�ޛC<J	Z��2!��y���۲7��R'�S$�9����?Ք�W���Q �ĥx�ac�"�L%��C���z���
4�޵����u�N8�����s6�������{[�\������������>r��h�K�7}+����e��Ý��ڃ��ǵ�]:Y���+�kڮ+�+��m��QE)�«����xr-o�n�jNt�����B�ǎ�i����'�����=����odb��Zq���k����8�dǣ���z@�f!�f��,HEz���l�z���!I*�ư���L��I�[OT�5!����o���jdYP��G�V���\����k���m����ċ|[�H`믿�8�~����<�b�^���>X��@pNH8�}ʅ��~�?ȴU�S�6�!�}X��g�VR��r����!���E�t_�T���w���Hja| �H��d�}���E�b;�RI������7B�w{,O���Z�H2��8��UE��t��G���)�(^0�-n�W�B�,
�-�=��j���C(%��h1���7�R��|��8���68�xQ�}�Ymw��1�be��l�;��3�I�"�e�Q�@U=�J1�*H�@�$��z� bo�X�-Q{b5B �Ȓ�J�͙a����WDS�����~�W��&�]Z��B�V��0"��A������j��yKT�{��L6��+��j�L���IK<su$��g���0<���w����8,q�9Ӵ���u���U��xw��z����qiu��J{9�(�S`���e{�&�M����W�Ao>�s��n�8�s�1LܩNa�J��w����=��ߑ����mU�G���8���*���6�!�8�̒2(d�Ȟ��x8�
��?(�p���Ii���$��;D�c��ፖ����5��*���Ѣ���QʮMS�\�2� ݝb�(�,�U�	�խ�w�wGM�S$%a~
��5ү�es�he
�����;�{ؼ.D��n�`&�E���?�]�X}Qm"�k->1@ٽ�Wg�H�i�b�/�(�1Yj�S5�hW�b�Kr�,�4�a"`��QV0���ʡ����xQ�|B �d[��R�	�[:�`3��]�O5�sg��a�;�[-���{~IW�vg�ֽӔ;��֤<u[��Q�=�Uj���
S�<�K�l����tSO�IX��?߳���dq_�:W� �R}\h�q����e�j���mύ��<����A"�f��?e���c����!z�c>��Gx�T�_晞�0�?�c�{/�B�,6>P�PS�3�G�����f���O�Ɲy�n[�
�o?�X�>S�`��%�����"~'�l��������gt/6�֟��2���:	
����N���J� ���K7{/�|\���� ���v�=8KUv�]��<���#����.xɰ��+-M`�R����M�	�q!.�R��3Q�h����*�s�~�e���H&::I��g }���I����F�*�qVM�SK���i����,#�����`�U{��ݗ�j�)�Į�7Y�n���}�N��� �#�J��¸�*�Pߺ.�9]��"S��RL��F:���l3:~\�Cs��1�G��v����+It�:%����YɅ�]V� �m�w�ȫ�[�{���")
5'�ns#�5���v���/�C���?`�-�OwR�<Li���F�t��)��~�m�0i&����УV9jO�u�����d�=\>%�IR3�0�W�ͻ�^���-�7���Y���1�O"$5^��~��~x�өi���Q���;���^(�U�G��*��%n%����������{�C����M}��8��z��G�cOo	�w��?#i'�O�!�bR7��\��IP52�MWB��㽋q�ӡ��~H�9��Vv�G,�P��Z
���qQ��Bn�|�0U����Cf E�4���`��g]=�����C��y^�2P�e�V�s0�\�������<]�*`o�����wL��F@;������U!�4������y�q�JސHS�(^�N ��7����8�|ߐ�O�K��-��r6%����<9��T����́��Cx쥁�)o<Q];;�wȎ�9���:�c��(y��V��]���Ac�H:�7|��ٽ�	æ&��0+@g$��a��"5��0���MQ�>a֑��»c��&�i�<������W�٢F�R|��8R$���zs�ٹN��c'���z��A.C�DZ˽#�_�|<B�@ �,�Z���.��m�?�B�q����D�l�7�����6�*]N�Ƈ���?�G(�΀_��8۶噹��z���.��������,�-#9�t����@QA�Z<����ˣ��r�:�UB�ٛ��bf�&��G%7ܫ�:.P�]S��@ِvrM�=���M����$�s�{�_�zt��g?��Z�O�ٔ �3�U���=�����t_Ι"�6�������/df/������5�W~��Bc���"�-m���R��A)t���������	J/�4.��8��y����;A�������G��-}E�B�qk�̶jת%�yL%fq�6��^��x��T]ym(�q�4b3�����նt�Z�_����x�ߦ�{Z��V��u�(��Yf���Z8'i�؁6��Z�ÎvU�1�l�Y�`�*}�����b�|�V���8�D*�A��:�pH(:Z1p�Z��s����#�|)i�V�)H����
���bIRXO	y��J�l�mʫ�UL�Y�Բ_���)vzv0�cK��g���I��T���]Pq�#_�Sp��+w���މ!�\Ϣhg�k��.�_�Xw��Qoc�_�J��st}�����q4S�����E�
q2j$�q�U}�!V4�T��lQޱ¯�����*����YwVf��}�����e��A(���xATD_�'���\���#�O�-|AP���R~�l�.~2->���vɍ���.��,]�O�!N�u.?��n����Ed��l����ٹH$%oY���4.k���cu�u�"z�g����t�g"�����X,���I�̂����Q�������>������kF�V7��2��j�
���E����P�V��T?}A�SߙY�t����`�˯$Y���ű{��{�x��1���C'�Z��G!��5�'0�'+i@�nH�Ň�,
32� ���TlW�m�*9Q���3K�:��C$/���������&:��c'�v�_wg���x2I�L�|��������u:���&T�妔�y�-\
�k#6������DX舃���BK��ӔV�`�8(�1����2M����º�ɶ��,-]w���6���./���D�&)+pҬ������]�8�1S���U����u?����a��ܵ�mR)�4*��n��`A�u���z޿Z������<}�t���i"]��f�%��P�@*8 ����>�����T7�%�e��L�1���Ĥ���p���#y��Gl�H����!���!��_���x�&y#�9�h��N��҅�I 4��&��?&a�������FR�h����l�{l����7ZE���j@�.�n�!sgs9���U��!����F�7MZ����:���T#C%S�O�h~n[��F7�~�Z��C�M�1�z�~�;�))?3���H}tsi����)�{��Ւ�~���e@J5�zK�a�,����-3I�bv�����U�kj|��
����B�{O�7^�sX�mAa�T|☧�����Ș�b��Iˎ���D���X
�nF��Z�8�QU����f'��gh�v�@y7��@�$:��qz�K��e�-�S%��yT�5M,=�)�����n���K���ڌ��Yx"�Xb��,���T@A��"��f�˸�@�ո4ԛӷQV;(e���C"ԵTؚ�fXK�Y��+��A"�+�s��ˇC��ө�������-�k�~�o<9��a����څ-��\���&�?�g?��!�t������
9%�8�X�{@.*��(�W�yךZɔ��j�L�1A���`��@){Xa��_��<w%�Z�(\�f�)a��M����%h,�!&�|�`�v_�U�^�1��ӪA����3a��=D�m��cl��u�Wj���M�6�M�vYsvy���Ѣ3R�(�� �҇���/�(4�T��3��}&�s{���a���M��+4loKngZ����{A�����ڈj��Ay$�ђ�l�h���8_11�jy�v�M�cI�_>�\Y�VL����uv�|�i�l����e=����Lχ� o�I'č�h1��_�7*�rb�$k��;�^};B�R��j{W�����<�V2��}[:��JS�L��+�)�@�[e���i�d郍�m��fv�I�b�텪��;�a�K�ۭ޼�ID'�(�������u�F��M_.��g�$th�j�m]f����Q�ޗ�5Жg<�|3LuĆ�R�,��5�v��ʍa��ړ��d��ƚ��?H�&�5E���G��l*-����H>Ss(z�)\1�Ȣ��BI�x\0�6�L�'='h��Nc}��9W��֣����PR(����n��)��v���̑-��}��;����$���.%_�d���3N�='���vy��f�,W�����w�9���u�H�!9��ZױZ���x���Ʊ����ї��34K��l˕!IoxG(���Y���Me%�rJn�LS�Q%0w�����D�nuڵZ��Q�/�N�abInZ߶I)���I#�4�`�atW�| 6�<L����1�ڂѪ V	�X���\ͽ���+��(uX5�f��@�럷��}�"/���gs�OS�V2��ß���˱�ה?��hA��)��˛�y�Av|�O݉g܅L�Sd�l�R�h��~���c7Aqٶ.��{���`�Љ�6�H\.�Mw����hG]�����b9�=u~v �K2��[�j��]��YR�a��j��D!=I3�$1=h�{52f4L��
K ��L��'DȤd(���D�Ős����{�T�m�6_hf7�v�~�C�rF�eE;��-u@�C��rz�M�g>��}@�es�׭�';KD���1G)6��=��g��9�Ոێ�(���y�eU?ݬ�iJ��U��h�}��ku�^։ч�ͩi�{s㵱���G0a�������SK��i?�Ba��M��BG0]�)}N���8K0�p�=:�3����ڼr
[#~k�Q"�M���"��<�Y7T�&�k����f��8G�?� ]�g�얇�q���V�]A��y������E�S��3{�|�;<�^�_7���̳�a���W�ܾ�)�b�׊ψ<�w~&��$�D��sK� �f!+\ܙ.>C���j�5�r呵��]?�
�w���3�$#Z�}�������5��:kly���|9�wo6�qwZ�o�����NUA�[V���t�J�Q/�F`��fcX�:�����@�uoԛ�d��v`�Q�0�W+y�d�P#����B�Τ��ZW�%�vz<(ubք���!%`���
��ȆS ��/Nf
Ef����;�䁼��O/ Y����B���=0<Mj}Y�䂶�Z_�-�ʤ��oiu�o��Lﾘ��B�����E{���KD�*��5�r���#�Uߵ����<6|q��!��#����:}�|��������`����N��}˄��C�Ժ��ܒ��mH�.��b;X�DqMzW��)�X�+E�o��;�3�PI��n��I6��Q��������s�9����P��_巳x7���~>��{�PF��qt���~(0�N��n��2�F-����S���w0�kNw+�m2T���4���& ����K��k�Rcc��������}`#����UI{pSXM��<" �D:�@����Ҁ�nd��rC"��2'�R��߄S���#&�
�#s����{Yb}襜0gk|�Z��~lQW}`�a��ސ���P�m�m=�e�mO�����W̑7Y�\L������C{E���*geC��g��I!�ƿ�t��Pȭ_����d\c��	�O�G�0�"���� Cd��R�����;y�����Q��y��i�r���W<��pbA��I�h��>	T�0>�e����@5j�����4�-�^~W
�����.�-:�a��Y��#��ck�x ^B�H8`3ɂ�Χ�}�w���CT��H�l���������4NcL��5���<��v3V2ʿ6��}�ڂo�Tݭ}+��1������"���� Va�jR���ȩ7�����o)&���>sqqϪr�f���J��P�o��AgT�x�W�q�JÜEL�'��n�?����ܔ����q ���$5���y���c=e�d=�m5��Q�Y�t܊cJ��fj�~'��A	�$Ѥ���<�*u�`̦EZ�L�WU��*-g�Co�2C>�4�A6󮏷H���d�ҵ�8UkR���p���k�����V��Sιb���7J��]��@��i���ڑ���~�����{��u�S���1�$I����Qla�9��O�_B@v%B�i���n�κ��K�*CJ�feo�T	_J����G�o�����U�&�)�t�j!�18�t�%R�EM5Ճ����9>�8~���D�t�cF{h������� t�5eh��n�B��R<�� ��V�#k�l�O�����.x[e�����f�� Ȉx�3ָ:�%܅,�ӫ�I������ʐt+�3����������y�ɽ�f�ׁIP��l=���~?V�|�M�nYK/��f�8��v�l�b�A���RA�-��G/��9^��KťZC��B��=���_�#��J��n�&�E��n�`V�9��37���@ ����A���nE3�.a�3����S����_N
��ͅ"�a[:a���6՘��$������z)k��i`+�X��^9[u�%SηuJ�����,� ]u�]]]V+j�����7��m^��ɹJ�&^�6�zԢi�7T���>8ji�n$�4�g Υ+i��M����ewǗ&&`���Y�b(
O��f� %��I�K�����t2��}`3�I�vB�X�?��C���y�t~�N�!?��`��̤�V������:OK��۔����i�Ep7�7��h���2���������T�keCM[=^g���(�9�l�|����Vy�=�
R�.����(���DY=��u6oʗ�I_���Q�i��Z�I�����h7�1��(*5�y٨�48H�<�ꀠ߈���4v�4��D(�	I����8x��	҆M��B��8E#w�斶���iEQ�O�Z|��q�B��N� �T�����g��ӖS�S?z�R*i�\\į�qIL�����i~����.���o#�z�J ڙ�\���P9�ҧ��K�^0��V�u3Fl���uz}9�
2ۍ-5�����N9�Q���p�C��Ne�.`Ǵih�䆀���Ǫ��_w�0�"$�~�]|6_:{Z�suJ�.g�x�I�K�s(Nӑu�i�F������G�F߯Rw�Ǚ.�u�C���n�n�'���<��\��%?�4s_���XZ��+�Z���+k\��7C��,� �L�NN�Q:�8���m��Lw1�h�sJ߾�%�eISJ�t��>5}�gc����04\ڊ�bqO���1�Ab�#vL����2��T�����	�	�"FP�y%x��QSO�OX��T��YxO��پ�s����Ȕ��Ac�6`����.Xy��d�Ǡ�틑�MO����A�}i�X����h�Z.����,����<U1�G�����vxC����*��%~��ů}G鞃�a�U&^�]�p��P?$D �#�h��aZ�� �IJI�F�ɬ��1]�Zs���^@��{�ʐ���~'?���t�\���ӛ�}kQ����0삻�[h�"���B�>��	�����~4�j�<Ke���I�d���ܪ�����+����;k�wRG�_w�4��5Lȟ[���PCU�#xV2ҸS���  �E����3��P�n�Gh�׵���њ�8;���.6H/(�pm��eB1�9/2
Y��P��Xx��y�oOy�B�ǌfNyv� 紤���aL�1�V�#c�t�}%��$�Y��1�Y�Q���Y+��rlض���1	�2�w1O�����e�8gP'3�aH�8��
h��om�=Kr(Mtr/�1�J�ԛE�*���f!��jڥ�B�tk��DDߥ�DC^�ȝm/��a��°˲��P3�Ɵ��&8y������!����?�KZ����|�u�F�IC�z;�u��%{�l��A�@{!�q:a�@-[�K��SXܦ61[�������Y��"���� <˔��q�b�IUɠ��Z�;�tx2ѢX��n�ۯ?�̉��%����8���$���g�1ba�"#�����;Q�J�7x��m����jEU�]�����ݒ�PB�P���\�D4����X��w���P��&@��
zJ�{��ۈ{���W/���)x>��.�SP���ѫ� P�H��ߺ@��n�-8�(�gEcDǖ��KF�&�C�3���ӾO�o���1��o�y���]a�pJ��.e������;���E�G�V�FB�?b��?�Ǫ�\����?��
��!��_W&���.��"i�$<���7\�,�r����DV�%3��'�L!�񦽟+-�!oV\FA�����*?}��rUz�Z�
�[�RĢА����uqwPam��y��-�@(�fC2%�Fy�����O��:}ڶ��V���(��Q���a�r�؎�u�ވ/p}�w��?)Ah4Y���f�_2���3J���;����Z�X�&ŕT`w�g����{�W��3�B�.4��7>�e�.��3!��ކ�h�����!ۚ'
���-%�An�^r���!��qLYH�%���D�Zt:�ք��+@��ѯ��F���d?�$�ӳ8����%/e8y�v��Ȝ5�&8����	F"OU�1�:���16�l�U�u��1�4��Q�b;sQr,o|���h܂�öC�)�&T�Q��XI�3]#�X�N3ϸζ�F5L���yx|V}Ko9I�.S��8~����� vG[ރ�\�g���ڴ�m?�m�2��}&� {;�t5�t�O�zAP�޴�{���Xv���>�5#�s�&��R��4�g�������Ҳ�+뚭fp�C	��9E���Y����x"��yF}mAD�/�����Trs2i�Rm�C}�y��PF���.�*�Uǽ����
�s�Yw�0$F�Q`�)��v��ZL�#�G���h�<܊��Q\��S�	U!ŏԠ��
�K��Ȕ8���팒�@���/���s�]4�d���d,��;�è\�k���]��gi��^�#��.w}=�Pl�������~F'���N�n����x��@#���n�=d>*��\��@�w��2o
�*U��i�z�[C5��Fϓ)��Oc�kYD���I�(�������f��� zT��s|����@=x��j�3��Z$-��}3Srgy_�^7�*qw�95�{��x�?�����pz��Jw#��|"E���>&B_���� ����)���m���Ţ�G�4�����Xy��������Kn�W�y�Ǘ,	7�{��qsGcK�S��(��(�B�)H_g�G�z�/5��"	*PF��k*���k=1�<IN�Ő�����U=Y�_<:��:���9���DY�RG��K&0�dy��[�lX�����2�]a�%���?r'�5ǋLF社F)_�_=��`H2�a�G�.�(o��r��<P�=
���r>bo���C�\o`Є��2��y�
:���MA�[C����Q�\ؙ$����h=�������yy@���F䈣���rDJƔ�9�=��x�%A��w"y��F���,  )[6��N�9��^EW��K�
�h�b�OB*w�2��Дr�bB�̔=��3� @V��jT���=�z��L���[V&6��LP�d���� b�rh(��v���_��<�F�܇�fiɎ-�B���s�(yD��'TfE�i3!5Z�`�o�#Ll�Ox�G���c;�Ɇ��'W��LS�ףk}�t9Uk
�N�bW�����A��*a*� J�մ��ΡL����R3�΁�ل.���%��㮀��l��;a�U�e�T%��#[S���jG��F����������[�]a�8T�L���D��P�=�ʀ�����:=e�'nƆ_��b�n�$3j�é��2�z�.�{�胚�S*�� 
d�t���w�H���^��V��C%��26�>��m6�b�/�vj�=I�l=��(]��Q�yrK��\� ċ�%��u��S w�y�����yx]��<�q����̒V���_�N
b�W������pf%�?����������G��UY1a	�l�<�`��\qbpx����a����j�ܳ[`eR��*��핇 �ˋ�=z��ǻX��.�)B���L!�
c��->��"\�O@����j�(ڐ� �ie�y�=��,��t3��!��^Z�H;��N���8M��Br�(�L� u���0v���]5]}��f{>�M7M�S�7���F(gH�k�4J�=̛�P�K(WC��,���=�%gfp&#��4�n���e�Hh{��Ϸj�_'.l�#�t�VV�6Z,�E��p��8�3��}z�q�c(>��#�C:�\XE!
[�$��jN���D�H�7;+��=+p��8=H�腓b��^v˳쾠=0� �Z�2" �rO���~n�Q�l��u�k�$?�
�*���ʮk��>�����X~�އ$wAsuR�?���	���X�&k�<�ߙ@]������9WO��v;hb[1k��\7eӔ,`��PW(�ށ�Vt��0[��h#�H�dxK5 x7y^ʱ6�d�%�ȃT��,���
��$�E���a|���[�y�h� ��֜�+h��Cj�Y�X��W�&5�8(����j�����m�YV�Q9Y)��̍A(%X�B1_�7���BBx��iŖ�Y|��gH���1RS���@e�<%�%M')἗�S{��
.�h�Ӊ�)�ܛ�Z�~��RQݽoMLJ<0�.	=�%g�G��NR�_��$L�a��$��#\6 ��΍�[J���`��^0kf|�31juXB_i6�N���Z�}��/K=����[f�Է���]�ft9:���a������,�efq���qEa`�6G�r�Tvq�@J�"��q;8�
l.m��{=��K#v'�a��x���B_#�4����tCAu��8���j��$��&��|�(%�&M������Gc�0л���r����~����m��s�'��xT󏃒n�X*�6H՗)�Z!�n����!(̚	f˛�q��20&����37������_�I;'h��^^_��<��\yPoWM�	c"��N�w�0��슻6,	���D�j`�?X�1��,�@h2�CI�r&�%W�2v��4���|��.��4�P���� ��H�:ߎ�rR�����T��A?�3���:�H��������\��V	�;��˱���*�6S�t�5t^���<�.چǯ+�V���J*�7]"��}��F&.vD'7o�5/`�����ֿS6���gG����_�"1��g+�rb>A��C$�|�nɍ0f2��o�k�K���Ȥ�ž!�}W����-^o��%�.��� �q��겤 �8�������4!������@j(y��=�!�c���$�>"�v�m6��(Ue��u��X��Є5���r�7�(AZBP�Z~�r�뒩�L��k�A!S��;+���7����G�|Ax�C��������YkR���62�r9���t�
�g���Dk���������rt�T�����8q(�DZ�����eg�=��[���v�F&l6-!ңLO n� ���-~��L�J�{��\#�$H�'Qe��q�_
���Sᝤ���?�x�lt#�9G�|�8��C�.[4 S9h K^,!e0a�,��T�ҵ�������f+�F��vq�AbY�7�h��f�8P'���L�1R��q�S҉�7�X�k��N�
V7��<�Q+>X^S<n%���;K�5q,��#�jsJ2��a*��zLv��
������'�[S���n��� ���Ǆ� ��יDm�A����RT�+,1���"չ�x�|���
.!ۮxZl�� �?���ς�8�I��Z�ٰ#Zh��x�hU}ROmL��,�%�u@I������^\gMǏ����dB���zTQӈ"`��FRv����=���M��?�P��Q3r`/6�S�,���żY����m&�x���l�!),���$�����������A���w��Oɲ�+�c�J�n
����3e�ˊ/���$��+���-��?�����i�iǿIK�[��2�
���R����ݾ��J���4���^`���z�^������Rg�n��Hv*�F8IO�����a��N����,i�K~��R���q�K��EE��58�E�C�4����vW���E]i����	8�+C�&��Z��*�ݱ����:d��{:q}H�x���i�����NRM����Үk�}g���Z�ˬ��e�f�x�4����r}���ApMP���8fH5�2UH�y� T1���i�$uCZ���� hh��b+Wv�K��!Ϟ�ŎΞ�k�MJw�0����	v�^���7�v�"�G_�e?�������ߠ�Sd�C
��dR�|��πH�ݮ́�څ���ۦ��2��"�l�nđ��1��-յ_4>��?��&�5Ķ��wq3�W�����%��yω����23;D�h(w.�� jA���i�)�J��Q݊<��܀7�Q  =�a��j��$�F!]��k��8<���,E�SL��ٖ���6�o�@��"l3�����{"����p�)1���<�R]�����5`���)�Iӕ)��@bc�6!�<���;���c��WN�aV�=�����^��FTH"m/tˆ�3��D�Z^ڳ�\E��epQH��ݸ�	������iET�WB�?!��4�y����xÚT>1�h.n>��q� %_*>L�3-��Մ,���^|����I�����@��l�
�7�����=�<M��N��&�ɝ�m�`ޏ,y���3/=Y\�7�kڹ��ؖ� 
���5�A� �4��)��+`(ENR�u�#��w(�lB���픙O��.��y�Y�f��Aڄq��a�[���趀J>>�3/����5�ʿ���fmVE�E@F2�Cȶ��Ԏ>�5�x�V�h=g"/�L4��{#7���E�QN��q!h��ņ]���1ײ��Pi�1��9|�֧����%G�j�#�[���U�q�\'IN��<5?��(M�f�n��j�«�|Yנ.���ڴM�7UQ~m���3QR>���	���՗�g��Ӻh��z�n@<�'��đ��ʰ���Bm���Y�7�#Ƞ�"����̄�~���1Y�Χ� k l,Ԃ��˺iY�{M���sr�mEiJ#%/u�r �,WqU�������LC7� j��7�=:�
������D�=���5���#S��t�J�6����X���`$
�q�f�y����Y��\�a����;Ҡ0���B�F
�S�x��j� ���u�l��Iy�Ø�Q��S�J�Nka=ձE��*<̨�eLh6���}r��S!0���r�͵q�!yF�>~a�O]���wƬױ�a��K��t����'x�@���!���^���T��*�Q�z���j����^�N[
�=�h�|�3�E6�/����t�N�����s*�E	�Kj�\�k�|�y�K!ʁ}��~|8�KC<I��P��m�߈������~�hl��خ|<�#GB�(T�~Y��2��'*��EI���-���!�	����Zh(N(� �YI�"�@?����N�l��sD C�8~����0�dv�߾�^"�ۮ�]ᙰ���p	�-��Ǔ���f��"$��b��X��|,`��AuA�B��H~��N+yw��J�ͻ�����qL3�۩�>l+'���[
/d��O��(��%��p���\���2�|��Rf� ޫ%�fM�sQR�?E@�ht	��yXWc�G��p�����]U��r]MJ�
Y�G�I/)�,�nU %�?������ݞ0+:�d��O�j�u�S̊�%`ʱ�w=�ǔnn��pA�K"�� o�3����P�6E)�p���%��|i	*�|���C<�f���,�]V�M��69�;�����[=м�X3�`0��5��#$�R�y�ϼRL޵tm7AL���[W�kVc�F�p_�Iܜ�2���{Y���.Æ��>2E)�@)�z�����(�ƖƖI��l ݐ��sLq': 	mm�讵��ye�x���@^�7!{9x�2�1�{����3m\��^��8�U�V嫬���+Q�´\��Ym�?=+�3��w,�F����U,�jix��,#�Ip����H����YU����2j�)M'�v	%Ԗ�yT�=��/B�a��y(BF�K��&N4�($w=O"BU�m����ڻ۩\�m^`�O�r{�Orq�c��ʋ�2]��R~ԃ��L�"0|`�2屫�C;�/B����&���E���>��E�m6Λ$9c�?E���x>���Vv�W�>1]c<h_GaV&��JP�r>+�f�)��x� ���`���Kk�����}%l�W�;�A�!�Ru��ݭ	��?2�%^���BxG���xfv����LYU@eE�U�w���J�\с�9��8]#E!���?����q�h�y�I�,�d��GjM0	s�
�ۼ�U�yn5��tgص�r��[����svN�oT�����s�-�5t���7�?�:	PZ��:c�:��c;3��}7S��^�܆����o^ ��o�A����:����=zX0�	�m��@;8��FmYgGh��M��$-�	?�%BU�����mȀהG5�$`�}���'��T
_am��ˬfp�@����H�౬=I�U��Ln��D�����$`4���j���+0;fou��U�u[��I��.35�N�-� ��}оn��2��3Ys���,!�a8#23��g���7�ˉJ�N��U��u�2��t���\��UyX�e���胞뗎M+��;Z�� ����j����	��������!�+Ż����-QT��_t�1�HĚ�/�F��CgP	`)�/���D]��:m �f	4�(��Լ�liɓ`�s�gjucF���U�ķi���d�<��5�7�hj���7��.����Y~`�l.*,9�����մ�F��K�$@����[��_��F7{=��:�U��x2�ۡ��tV�@]�ں^z�T�:����,�L�4v�Ԗ�S��h����ؾ��ri��1��Y�B>�ä�7��r�Oj�X��7�m��yc��^K%�XZ���[&��\&��QA�*�Y˺�&�k�<y��k�Qez.�+�s#�Y�;�2Z���L`�Tu=��;R�/�ڇƧLLN�}.�F6,�v?�r�ҵ��+Ӻ�{c�v�(��<�J|����!`Ւ�ựk��k܁�5�{s�;��� ϶��B0gw��5�s-��e怊��^ 8�;Z%o3	E���p�LN���U�X�Q���b�,��E���;��Iפ'I6ro���y���0�~s�2����Ջ�v�s_P�P�J���!��cL�p�U�Vn�h��Lm?r3����Dy�;��E$A����VB6!�fT�~\�q�;�Fj��e��(�^��G[�Ä�&`�����"�҄�%$,�6{|���OL�;v���i����������俵E�|eb��F��c1=�_�����X,��n5�rFe`�G�7hFq=}<ʔ���shZ�P+�\Dh��i5�?�?4Ɵ#��d�@�W�+Bk���5��O�w�-�����E��΀4\I�*-������HU.�g�mnn?�0";�zT������4�Ml���b�ъ|�;G�������!��:��(O�j�,�W�^��nO���]#�;(	�ԃKpU/J����Ey���R�,�T�U�#�-����yc��a�?��	o\WBT��f2VQ���&Q�0���v�A�=��Ň`���7�@�!��35�Q�~���Nj��@�M��$x/f"1BA�sQ{n�C)���ӿT�T����V�,�iX���FpGͤ!��v�j�(,��Dmˀ!Q=�w�)��b
%�<o�Jҧ�Wښv���x����ӻ"Af�wUz�_cJ`Nq�c����њ����lKX}���uQ��p:#mPF0Df�/�ì���X���R�kZx��d�z��d:�|���}��35�Dd��v{�����+����Ss$�ԓN�a)���y��ϒ�K�B�!�0w(�E�� ��^�$x =�L��r ;�|�v����\�q?�)(�j1��8�F3ӭT�5 }��FM�A��"��MY�4|�v�a�:���j[Ʒ�`��V�9�7��FC�fF,��ݝ��鴮x&�����8�YYR�>�!��Ҡ�@�Ry}���B��̛����\P�(�Y�+ѱ�ZP�>����>���*�\2;�"��Rp�驜:g��gY�xJ��hACo���@� �d���:��f���խ[��w�%U\n���a�c��y�C���?^wL�_3�k�㣤�7(�E딘�m;�w"_�Vпo4/�C�ѦC�w;:���zr3�)�\��M�~��l�T$f��7̮��E��[� 3}��|��6i�������#�&^��, ��s�5ǔ1!1�[O)�n6��]�7���Ѕ� {2�ڄ�l�2n�R�6˪hz��<�
�!S��>3��&�`��m�=먵�	����Z1��ZUiH �v�@���A�	s,�b{�cR�'!>�9 � s����TnZ���t�{��)�f��'2e��'G��vvV��fT�nA���M��+G�vB&��L
ZN�K(m�.���5�������~�b]�m��4��t��肢���F���<�W�KZ�~S����C2��G�"��bg��`D�ЗC�j�|�Dڿ�[�'�w�5�|S��?��f��|�'��;ML	�&K���R����ű���|H�5;p�d"�A�v?�=�6,4�4�G�_@�r[�a�s&C��ʫR��� ��&9�TI���*�Gb�E���b��ȑ����R���'޿:a�"�뚛�ھ�f�uq�<�N�8����P���Ip��4J8c��E�Nػ@���a��G�֪�)@�����O��,�F�7na�ݠ��H����Q�g��	�dʰD�	�Ne;���)��}��?I����5��N���JV�s�az�̀�v.�~��<�:��䑵��P<J6ޤC'7��Y;�p�b��4�~��gI����{�n��
)��O��Nn�����	��1x̬��ec4��]���?M��}9���ω0��:��6PuN/d�f��H�m�tP`A(��Vs
���9���	��n�ɉf��s2>y�?��d�神}��غ�P)��AmI�(�:;#@� ��YM���A{���WgR��ѡBQ1�\��YרEH"�8��ηGf4{h�h"���,�W�`-�E[ދ��T�\؎������ɢ��GV�tW�\D)��F)��L��4��XNi���8������<Q�X�������/	C.�W)�U����$㛌Ss��(����GdW˱���K��-S�wP)�,�Z�5I���B��ϼ1���D��)�k�T]��tx�I��������x}P]a��n��Z�
h���̻_��2���$�9�9����ySlR������Cm�� ф��4&���>
�0��$:a�J*�,
��w��Y�d]*�#����p� 7�Z������LX$�+֎�Zs���xy�f�6�2Aء�gf۹��|����WT��o����C�q�k�*���#%{�����-G�N*_5��He�����
�[I�*�OpT%��\+9�{A%	���¤N*$=��Kd2��͎� ��ޕQ`^��5�F�
]�S����)��ӓ�]��'��c�%
:��V�p<`�M�*u|(?6h�,�r_ -�g�_|�w����7����9����}2�/�#̻?��HcB��b�7�X��
�I�p6��������?˗7sյ��)B�-��5�����*������R�A;���f,��s��jS;L�p�W@.a|N�|	^�����U4���UKUs���Y%G��ꈜ!�C��MpUڹ��"���,xi/�S������t� ���f��l,Y�Y������P{u��) Qb��q]��N�P���F�0S�Br��y|/�P*�*��N�px%���B��-]��#�lw������n�����%L�.Ϝ��Z���ޑ���>3��vI,��>]i�p�t�3i�K�q���=�]��-���4S��"-�Z�U$Py�(����9��Em������T��4F��L;��MF�!{��a7H��1`x�X{�yQ{.�(p;�N���X|K��i����6 �$u|�W��,j8�F���U��՗�l�u�2�φQ�3|��3� �b: �5K}��@x�4�@K��/h��I^��_�?~x%m�{����Pjl>�?Jŋ��]Q��)O�C��S-��9˫�\�G&���Up\���ƛ��w�P�i��+����;��Ʈw:�	