��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�]��Xȭ��p�oȡ�;u0ީ�^�)�>vys���2{�L�~|c_Iy�K����-��9!��\�Bi�D��{�Ԣ��r'T��NjH��ဣ]��9��|p���4d�#尭�ǕmpC��՘���z����m�0��X�fծ�+oa���}˗!i�v�:¢#�������Q���*Ӽ���	�<���������VRK\	���V"�(��wG>��<�4��ԽB$HQ�U�޺�gN�*̣�������&�6�\���O��MIB�
I�,��R�XT`���ׇ���\��y�`๊�]&�1�4ɻZ�S�u#��5eQ_���͏R��"Gi��� �)�
ǯG�0�V�Bي!�=�����Q��"[���c�o2��0�=�!2�3h��5��H.*�>dMP�P��ަ��~���u�s�f�UQ9z<J\����C(�C��+���r�)+��/��$� �3���;T�J���O����X �K&���*�@1����0���]����~��;k���R� ւ�NLũ�4]�f�����4l!&s1�M��!9��ߞ�]�䷬���dҴ�̣��k���$��d�~�|)�P��I$:uJ55|W/�?|J��Z��M/��"�Wz����l���)]U,;�F�N�
���O�o�-Μu}�}�܃R���4u�d�y���c���Ǔ��/��b
������S��_�;>��E����]J
���CE��Ϫr��"�����[(�O�D�ҜF
�W>�V���gᩴ?dѓ��ͪ'!J���V��a�r�ω�l�5qA�/w��~��@�n>7��h;�������}��O�ugj�Խ�	��-�e?`5m;�u.r�{�%3X���|+����P��Ӫ�k�Ig�#����$��D��r����<Of�4���S�3p\�����w^7�\<���TI	C��ȭj����h��q,Ʌ"��ԍ�5lV�\%��đ-���O��\��� ��o }� cw�Հ�����:�OEK�=՛�<{���D��g���P�0���&;̀��S�(�W��;hzc�d�������]�H��0�iVqȟI�m�Ƙ�2��hW�4:62����؁)k������U��";[�1��!��@��ຖك8r��MPA[/$t}���%�%d���o}���=:W`au�p�'��6G3�L�(�E�
��A��2�ں�#�����*ps��P���l�V4���g�-�O����ǹ6p:���f�\���ā�	q� �#<�F
z�����/�,`�C�����r�\4����%qhV�	Ϳ���+��G�#��d|b/�F"��̒`�����w�c����U%�.RHנ��@l�(ɕ����n���f�:e�_�)Lcc�'�ٹ91�w�A� �c3[D�A�w��\������Ő�k���b���A�5ju~��-%bakx���<C8�n�r\ 
��e��7��>T)�ψnT�^M"����8��N��B�<�������"_����f��:(_̨Ir�,��}�7{��lq:Yy ��,����2[�)��VzX�q��B��`OA��xi�Ҡ����� "j�=B|pT�]tlO�k��c�Z�Q��F���O��9��������O��&�)��;��q��qOr��[Sp�X��5,���ޫ|� ���!�J�_a�Ҫ�t�¨eQ!��^~s�0PѺ���H��@�%FWb�ʈ�.|�v�?
Ԫ��5&GFK�G�sH���ߝ��uu���m���̶��[Qhص��g��~�yT�Ġ.��=�r�����I�f��x,�S/$��N��4o�J���yxE5���Eiw4���Vfrtf�U�;�@�7��B<[�䃘����2܊��������LU�87���Q���z�?8b\5��t,)�p2�����R�r��\��[�J2,�^�?�s���g����_� ���&��o���YH��-�qé�M��|;o�� H~:�Z�K�h��4YZ�hG���3疔���8�:��osrmb�8^��r�H�[gT ]ľ�+�	��C��	����`/�P+�@�:d�[Թ	8�(��B܂�nd�>n�X)�T�/���=�ZI�\�΅7*J�����91�/sd�+�n�T�E�M ���tyLa��X�8ZH`��I�$��bS���1՝]���n6�2oQվ'��6�l$��������so's�Ѐ_�i\7�k$@�\�y�j+�YV9�w�0�K�@�w���`2��+d�ӑG�[1�H���	�B��T�Q���� �~��m��,�W�#T����� xF;=q<[G��,�9�:��P���j�h|+���A3Z�z{�9k��ʹ��O��+"	}5T�:���|v�q��XEH˳o33ɝYJ1�^4?[u��O=w��"��"�HaT937w�_�(�8wD0Q:����_.ﶈA0�Q�l�5�\����S@����
���W��f�ד� �w���=V�μf�����.?�Q
7u����V�B�[��� �z!�"VT�y�OIR��<|��`d7�\|�E�[e���tuJ�4�dg
|z��n�{���K�8)�ڗ�c���N�6�p z��\z6��N�~�V�����A�n�͸"�!W!��,�)��a{���7��_>�����5� <1�eo57�������q`MΆ(�ݪ�8�c�B+��x�	��Z03��R��r��1^��*����Nq�����Ir����U5z��4� ݶN�`5��%�Y�yV�j�$� �o�xnu��v���I��`m�OY�"v��-�Yވp�{�q��1��c��X��Fa>&:�\h�pOa��Y����Q�z����6;��.�C���h�rzi��Kb����6���t3�랕1r�Iy���1�Xx�h=3�B1(��2/9��zQ�s7d+(��J�4-3٦�ȋ �����R��$����A(�X�@C!�O(�����?�Yr���ro�
��S �!)�(���=KN�K��n#�3��˘ռ>4���]���_P�������ܟ��yⷊ2�� ����r���Ԅ_�q�$���]@J[��K�%3�����P�f��<
;�Х�&U�+�$�&��G^�Y��K�@��5�<%R��c��Fk�6�#�� t��|��A���II�S�1� �{�j����<�륋���C>�$�n0�0�LA�96{�,O����nJ�:���q(�1��|a��<���ܜ���n�`D��MH��ܾ_�tP�g}��F�u��z���u��<�0������@R�ua�RWG�05���LRO'[Z|O(���2�R���=h�v����|�ä��sp�-�;L' ���'<�\?�R�~�J�q?�D3�pq�����*�L�H�� �Q��%Q��P���l�cůHG�=�H�6X3RO�J��:+��h��Qv�C�J�G�/J0��Z��:�ނRC#??�5�e�@����߱���y+�%�#�G�E6UWQ�N}-NR�N};u�����z�L��VOI�A=׭f1��3k×�Ո�Nh|�f3�?����)c���ƆlgFwQx���)G|�'D0H�\���}D�?Gem~j|��dkg:��_��@D���l~m��>�Gwk�2jW�]�ud랠j^�0,1{+j��8c� -��o�͗�Ӥ��;J�Mc>����|g��s�~pˏi��`�����ڬ�vq�I�Z�}QL)�n��h����uX�B2`���!"ďa2�O#Q3N�&Y��_��Ό�Oz6;\�VΟ�$�"iU� ����`�,����M�:ճ�*U�T�I�L��~.�JWR��1	Ӑ�}ʰϊ�� �@�e�kΪBJ$�j�ñ[�e;�Wm�Dc+DwR��|2�SސB�������3�W�~P�e�e 	W�G�m�M���f������Y�rR=�p�.�C���s�6ȅ��d{f��a<
����8���Dmd����YK~�J��:L��|H�S9����V��U��z8%@��Tc�q���z(\i�`��Um�����q]Af�$ ��A6A�����I�W	f�^�e�+M��	���a?���
�<�� A_h~�;�gU�(,��G� �O&������K&�� ��6�r��i�Q�-�<om۝s�>b��=���6OyJ�����4����x��D���b�3�O�c�����'"�z�������W��������e	�}��r�B�O��r@�� ��+����ad�s�$��}���������q��j`�vEA.�}�}��b���*m�h�7X�&��\�Z�o�l�0� �o,^$��\�^�6�l�}�1"�����Y���ƨEi�J"�����#-���b6��D�@�d�}�Vp޶��G˓24oC�-"��L��̠ؑ%����h~un�[;i��N?� �e�{w�O��DIE�*RD��7طҦ8��,?~����l��'�_N���Jk�sx����g��/�'�r� H�Iq�(W�*�����F<~��b���U����J�J��~�<�n�[�u��T^&C*+`�������X��}���$|ho[�o�*�?.b�5\K����ͮ������B�Ej��m|ϕf��;��G#�%��պۿ��և��; �>��ù7Rqԓ��:���� �;:s���aȻ\��!�Kݎ���-[l��ӯ8Y`N���s?�
�1��>�y��j"���ܚ%P��C�d������ט��
KS�wj}�u����$���\9���'�"���W.�8�����~hj=��8��q���Xx�b\E`^�[wT�V�4)� v�HaŔ��jQ.�Yu[mI���v��I����u9P���
�Ӏ��*<zF7��$ ����J=c��u<|c���բ�d�ؚ��<+/g�vK�zG+r1�A4��E@_�#B�yi�Ks 7���	ޅ� �A��X���v��]S���;7��m�w6xL�ԕ��B 1mNgj�8š�{���>E� :w�j	(4,<>�|��v���.�>"�68�M���Cޱo$q��J8�!kM����v`�k'1`I]�A��G��)��C���6]vCgN'����bI��-���틐@������:�6N ��%]��9Rq���Pe,ʫ�C���6��2r���
�rn�1{�ǒ\߀#7�$�aہ��ԊQnؽ�}M��vB�VOf{�4a��.��h~���c�DH'x��W$�@�0�R�e�ޞ��yv�玭o���P!n�pM�h멏��xM�����ʃ!�H�P�T/o��c	�hl�ڂ>�7T�$�{�bB->M��C�p^&�+�H�u�F�6����a�,�]ކ���:��ߓߧ��`
��22�Vm�u�l+"�E�~b�2���`�"� m�������X��
c�s�;l�.C߈kԠ']���F�����}J�`H����V�LB��$�z�z���:����8�U:r�.��qgf��EYes$�%��I|	�P��@����gx�6��@w����D=��% ;�/7�͉�3"m���a4<z�!�3�y���Ri62=�q���N�(����z��Y��K��XS-o� ��A���)8o8d?D��V�q��,�nw劼+^*M�BD5�@��+�R,x�#w��g�sߑ0��h�F[���H�2�x����;F]��v���lQ1\�)3Ѯ�4�=���?�Z�k�/�2�j�R� ��ŢA6��8	<�L'���jÙQ�-�@��[?�*����I0�n&���!��Ӝi�/����0��T�$ekx����1o$��-����0�{����߶��*��'\���-�}�����J��{3��5է�?	ZS&O	��n.��P��2�?�@��]Nˑg�w1��z%'��^ym�Φ uI��)��k����?D��+)������`S���l�/Uq?�&��T�}�h�#F�:�! ��
і�'�G���U��m���r)
�%ӧ�"(�z�hz��F�uPX�sj��᢯i���U���� \�L:c�	rW�f)�ZLc��o��~��?�H�_7G�z��ų��Of��J`@Ԉ ��!&i��r
� $ކ��lK�7~����E��[�Z�w�0�՗*1u���l�R�0�:��>��Q+]1���a���fy���� �# ��`sǶ�B�H,���#�y�N���T�؛���)1�\ɍE�����ƼE��84������b�3M��6y��[�|ݬ.�@78
��ƺ��	K҈w�W����k��������́$�L�A"Jq?��l����#�f� ��b�ᐕ+�G4 w��Q�iB����>UJs�N��[1U=�ZE�QM��N������~��
H��{�zh�;Π�#'��1"����Θ�I�V���ië?0�'���`W�Z�D&탕|S�X��h��	t�y=�a��3_����w���ښ���.GH"ڑ�W�3ꢕ�Y���qA�V�x�^AH9�P����;rBnU�
���`�ϯݵ6�H;�JI�u��j((=1�W�톦^Mm�R�(�v�������4 Q���ڹd#2wr`M�����őY��f{��|����{ا'�w�c�Ԟ�[���<�y_� ��`0̜Z�
�w	J���d�Ʀ�]�q_D��1L��R�`G)��VTؠaJ�{I(9iMt�;LpvI5���ݍy�O�h�Z��t� ߈�ùԼA�E=@r�&�=��%�����P��{�G��拋"m���$�:�d���Af&>ڛi�CN�b8� �f�Ҝ5�v@�#QG�� �c�S�GF�����~:?�a��$b�Y���N�f����^i�7v�$b��-��m��n4�%an8�B��K�G�Q6!0G�J
Lji�M��yZ��BCP������{���F�y,�Je�������C��J�S�����5����0�1-��2�z0� 7Ca�&+�����@�	���@C�\��]D;]�V��$�tn6��k�����9c���]yo���n�d׃Z��M=Z�C�AxO�5#����H��q���!�%2u&�TT�;�����Zo�A�mn9Q�k��'H�V��b�D�τq���GH$v��'�"*��b|�a	�:CP��#�a��Q^a�z�*�|��T�͡�ЂC��Ea��:�A�V�ڒ7)dtو����7�8�IjU��5j��Ք�� ��N��}�s�#^r�	����X)�?���ʻɽ\_ū�_q/_q~� ��?Q�'1��Q�Vq^IJ�z�+��PʂҬ��T6W̻�S�~3���)���#7�?�����(��8�kڬ@��O\�8���+��&=|��a	��*����Ҡ��~Ld木���8�*iCsk�f$Un��9��v��o�X9����� ]�c�%g�C��܎�J~��J-�������=�{9}c0˴��`K��g^Z+�b�zە�,s&�ȇ�k�_t�ɕ�p$]��԰��XO*w4�xz-���"� �b.È�(K/�ST����FW6Z&b��@���&@P%���� �5'��9�w{��=
�l���5����Vs��+�?�s,�2��J[w�l�NR::��q����,J��}i�Υ�l]��]"�z��l���J��������b\% �2ίm��U�v�O W	s�G�\���4_���[:�H��э���{��bZ�Z%�R2mts�Ͷ:�����	�������88���vR\l�.6Z ����/|�$��'y+��χ��c�9ﲱ[ׄ������q��;����!��WU����\_�2����O>|Al�_\�<����9t�zB(�����I}='�<���MA�����!�Rc�[��|dȯ�xZ��ًN�T�_���{����v^gn����B-��>�2����ltx���C���5V`P/y��9��ip���1筺;X܅X������j �"�#}�!�A粦TxZ��s�$���R#4���%�~�o��#�I4�<�镟�z&W�\��d�]!��;�o'f�eyL���{��j>������a��Xaar(�>6U'�t�3�l�4�-�G5�E*��T�����oΟ����H�a=x
�}�y")yZ��0�m�y�N����6���m/56a��ޮ�S�;5�ꍷ=��?���H6$@����.>N��&1�F2a�{v</��2�L)��H��{%Z�%��7��ّSz��y�g]���V�\��y��bX#�H��-3�Ϳlt6'͙�6�i��:M6����+H�� �;nk��$:'"Vm�wq	Fe'�dN��� Ɂ��Li�����a�"�û�w����w�֠@^��`@��^�~�؆Xf����%�?k{��h3����W�s�lQ椻5�J�Z���b�=�8�ө6tN��M)N�Ҿ�C��O