��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e����d���f{��@����S��>���4{��ת�AO�Q{����t�FuA��Q%�΁K��T�B�A�J�z
=i�l���SRG�/Ő�������ܔDl�m�W쯲����<^��9��Ç�lf+������Q|b: vջiy��Zxe��v���Hv~�yx����8g{s�FקO���?`�E)�����k�J&ˇ�����	���}w�hP{�A����|�nь�6f�U���` ����"����#���ZL�Y�2�$�A���1\<����C?*��*�G�:�YG����m1�8U�#[�� w���E�U0�Z��|�HL��5�&Ȍ�] �$��oT���?%�8�y��_z�W:��kV�ڛz���1����l��%'1���zN��\<F�CQp:x�=�Hq�!�_����������;�s��k10�NW���h��O:�u���m���;�]�|�Fϗ7y{*������3��%^���j&��r���K���Ahj��E�Wu�|�����q۳,D�D�A�IW]a��>�J�����p֦�J4��:ZK>�+��5'�#�s���"~�zd�Y�m�2��B��ɰ�VՓ�h#��"�(mzY~A�:��r�e&:�A���n� F��#�K4��-�9%k�߈�X~���AH3ď�um���N�  2:z(˖��t{�ڰ�Vi�w��Z��/F�c�(��%���iE���	���@*n�J�"�Tja��X��w��?g�O�'5Qe.�J�h-�%^�}���7p\�y�ʉ�`cI5|y;����ޡ�]�/�QI�i�)��=�+PlQ^&0��醻��G0��'rP�������%W��y@ts؂yg��Ow����$%�Ϧ�A$1_Z�AO
�ٝ�,o�;����i���z��ϭ����J��%�G\F�"�)���>�S���Կ�TO�+gS�Ⲩ�]ɇH����+'���}sM#����\m\V^2 �͎j�V�~�_H�����nq��xj��y�����p��VH��"����ⷓІ�*l^�Sz�pI)'��T�Jl������ե�3�|{}"����v��*�M9�[n�><_Ѿ�O��p���Ql�Sَ�2�)���]���f�jFnj9���[,&a"V�)�2���/G�4���$(RZu�`������v���{�j�4�wZzWh!z��NkrR�Ex�u�V�@G/��d� ����Zƒ��9�����a*�2�?9�׋Y��g�Ajr�!�"+��B]o�on���@�b¿�r \3|PN�����i�ڶ�-����J����#��0�>�p�4���@~}��O��̺�C�%ϱ���-p�| ���kQ��8^]8�N��g�s�g�qU�eSi�4`���a����w��A���=��>]�9��$�<�b��d¤��+{f#�(u�l(_���4�� و���3�����*BN�hT��ߚ�s"����k�!��n\�
5���� ez���#���<��ܺ����P""J�v��R�]\������}�m_U6���q�a	�b%�z�c���坫��1�U ���@�6f�M�_܌��J�L�o���u�|ᜎc>�C�=B��x��h ��[� H�f>OOZ���D�
F�l�TI�8�[��%�&#R����7�V�(8�k W�4fw�۫��Rx�&��<O"=;���l�GF�T�k�1����b(!@y:� �?��Oد1>�5O�0������Z���g��y�>�U��f������g���u �:ǋo�����"G�.J���_�;%��D���,(s�d�|�sd[�������Y��Ć�볛��Y�[�9�>!��>]7���Έ��B��ds8�ً�RF@y��uM��k��C8'j��	-i>�F��V�N��2��M\����ϯ�j�i�u0��`{��XC'��̍�&�cL�9~R��z�5Bbr~Lc��t7� �-�T�d�͎pM�*T����~M݋-2���]R$�"|p�L�Q!�q�R�̮=v�Fm��ɢ���Лkd\�lcLY�
R��Ȼ��7V �X즼�+Uǘ�7�処xy�&Pr��8|��?)F�sʬ���i��k���e���M���B�7Xt�]��@p�I\��ᙴ8��g�-��Ax��1wQ���Kxb/
�b���̷��g;?�Y��1B�ȭ�cf��F�besVnw��n�y���e��$@n[IԔn�F:����\@���$/B��0�,Z�koQ�.4�1�[m��P��6��ע�ST '���+y��ɠ�\��j�XC�GǴu���Lto�����h�֌�S%(�e&Irߊ�#�2w;9���ϧ�����X��4�+�$>/J0ǩ�TP�ޔ� �61f���$��/���C�W��2Z�RG`o�0�Լ�$�ލ)�G�m�����ž�j[G�^o�G�7Ӂ��J#-��2����Ԙ�"�.�~�cb#M�M�Z:5���X�<0��\^%7���4z�V��;��m��)��͔�$�H���Ҩ��+5��T'ƍ�;A�����Ŷcp}���q�)> ��A�XL[�����lX��L,l@��K�{�����$�MH���%�ٙ�w֩��g-��;9�����U��K�N^�e��[���|P?y���s���@��rt�j���ƵA�ʘI�J��b���E���C/�*q��+���|�U�Y���j��z��>�k ������^Xҫ]k��z�О��qt�ZefE�#�E��,�M�L#Y��FR�޶�1�����.���d�P�m+�<�1*)P]_����H�K)�3�W�.��0���8�~�R����Z�:���5l;p�4��9�-�4&�# ��VJwՐ�;�<\���X�2�e�~������=��es
qHb�t�zqҁ�i$[�f����+�<�����!G���t1F=��0�!G�YƖ	�2u��{��W����D�i��ԁl�^y���~׷��	@+�q���k��ȡ��k�_��Cx���J_A�aE�%�U{l�*�a?��!/��BQqQ��
��w��A1��x�_ћ8�y(�3�7�`dkF��	��#�K��%�g��\k�٨i�a��o��JG��	Ix<Q+�ky���;l�����Ŀ�'ρ�����J����1d�.���2HǪ���0�k��5����֯Y���J�-��Y�_f����?f��i�����5p��L��h���V��K�0r���>�:��K��kk�
q";�(�|ּ��g�]m������5_�ȶqw#IIaڎ�!WQ��n��A��;��Y֟�O�=���f?8�)�&HY��!�h����� .�-�Qݵ�u�)<�����M�n���ٲr��5B�oQ��y˂'�Q������Y�6"�s�d�"�0en���ji_�PO8�g u��3�g˳-�m]�݋Td�5gvT�7ʩ?A�Y.
�r���<��k�d��L�:�J[��t�;zĻ��P�[�L�j��^�>hO /Cr|�"�-�VZ�|Wr�\���wZ�$�^�%";,�g��j�B�N��@��\^����[)Ǵ��!���F��_���I?.{O��f�/p.g��$��II3o)�<�"g:֦�*P���B����tѲ8��*^mm�����$WE�������X��8�湈:��8�o�����5�^��sP��
s��z�L偧B�������q�==��͍k��u�#�[8Zn��dBrM�=�3Y���$�Mʵe�!�� ٩m27U�Ѡ{�%�NLs�oa�LI!�N����e���H�,a��fw�����ԓ4�#f	��������KM- 42��4����t.�ƾRa�1\-��C��/��-G�p|ӆ ����pEB�Y�9)�C�84�������{��.�gN�6�|���f���s�F t�t�Ζ��bn�\o�}��Sg��,\]�����{�����Y��	�lЇmt��P;^�ʰGw�BG��V=Ok {��>:�z(�L�ѤP���z�8-�~i� ����w�=5��"g��vݳ��I���Ao���ߤT&���67)�z�e�f����B �����S�����y<Wry��E��4A�~zMT����P��,�;��*坑�����S�#��e��ͽ�o�R˅�l���?/���Q�S����qQie��� %�\��&����ؐ�K�V~��IT� ��/�!ƾHu��M�������m����T3A*���ԱE<Lw���iL:�m�0�bҮR��(C䝄^���Y����'�U�9���V�@���G�vH]�t����XO�~���Moy�l+ώ���M���]|�q�]b�±j�f\�g�Վ�b+� e2�����0���S�r��}�`=.�Κ� �����^���GXC�G���Pr�]2�D@V����s���"��R7!t�S]����D\��0OuX�g��n�XT�@�9ͿO�G�ʑM̆�;�m�^�k���|&ۀ���W���a��#Y0��R��J����֎GW����L񠊞�y�q�O�"�C����[Ίv'���-)�1�Rb//·Km��Ըޣ�
s�����0i�H��]��J=0�D�BQ��?T1��*+�/�5�PZ��v��L�;r���Gi4�$#�f� ,7��k)>�^�G6/Y�����wF�B����̂�� �b�e����9�����C�Y��s�%F ��D�\��tM�2�Oiq�K�$�)eh^ŀ^���1��#aRNY5B�.w���j3�F�����y�7౔�;�.�m����q#�PL��Y
������{a3����TD����Sx��	�ؙu��`��_W� ���ZݥI:�uM^%��z�/��k �/ȡ/|�c!��eJ���c��Ln��v�Ń����`+��gt�?Hlq�R6΍�ŻH;	lb���)<0�]����H~<�:�.���U4o�^>3��p� ���P)��;�PH��k^�.�5���P�������-���R�7|�e�I5�x�/ʓ��Ϭ���q��jBE�` B�i��eK˩�/"�'���ݹ|c��a��6R|5#Pj�p����q�����ࠩ�A!��^3�kY�A� l��9הX}�j�.�VzM�Q�*1�/�3ҭ��z�3#�|�kƤ���m_i0s���ž����>�d2�?0�P�|�k����B�
�.�6�s����͍X~�qP��-��Y�J��퐳��
E� �3��;h�S�<�l�r�[L����`��1 `��T�;{X?�mM����M�Ě�X]��!�;�3�F~4���.+��Ɠ�ՌFς��H¬��6�3$|�y��yz�<c�;����ʺ�s��[����!��V@�xfD��B��zwAG��������j������`z��N�إ$H)���7�9���,Κ=/��՛NprLr��[@�}�vH���CP~��?ß����_.s��݌Z-ϐ����-4�s���o�Cw3.h����=�m��!:�ˢ��O�ф,k�h��y܀�h�\NQ��F�4@ �8��Ab�FI��C�j%+���4w��P�ʁ�z���׋�N ���'��Ap6��.M��r7�Z7D�m4��������W�fQ-߄59��Ϟ��i�68p�`���#�}"aK�eXi�a"e��r�*�]�q��M�K�N��
�DX�{��Q�:Յ�$��T4�*�n:�v�Q�-�-J��$I	`y�uf���^V|]�X�`�6�?�� ��QA��r�X�a��M,���׊/��P�><U8��7.A�pG�)!ǉw�O܈p������m�&�J���]w0���!o�Z��u� hp@��s}O��8���Wjo���O�&y��wo�d9�JRܰ���!=o�D� �}�4���[���<���)wP~��.:��!Ç�Rbo�H
:]%<�p�;hڱ�#ʽ�OQ����9�S�'8*˼r����;c��uRPD"eԿ�ޗ'�O.�*�������!(ĭqv(�!�US/�̱���:�_q��U��;���/����,�*���u�Xtuy�)R�輂e��^�k�b��u�|FI�1}�;ǲ��������m��)���m���mҀ��]4�B�������#�M���R���iS��1�/����5�~���l�By���\'1�^P:�5�H�T��Z.i���ʼ�A��ni��貮p���Tq� �$�h���DeiY�&�Q�8}a=�~w����Qn�^�k���F����5���D\��"���x$7��q�*[�{���r2�1l�� �]R���琘����W� ������
E�h��$��_#�}�^!�XǬ�~���M w�t�ڥ�i-��1\Q��#,zCY�e�2�̝��͐�lv�+J&#̰��\�U�P�V��>_^�`�P)Gu�M?;.ɳɡ��}��WG���aRV�����s^i ���q��b-\~�>�<m�G=$��fP
W2�>'�2�!Y�Em��h�P1��!�b\!�����2i���&;�o��Y��R�YA� *���/�IMB��,	�����(]O&\:�~ZsZ�l���Y�{�{}^��ݲ/�
�	V��F+��qKpU�%^�Ť��w���M��w����CN�N0`�5�M�J]��&��"�Ii^�QV2qb��)�S�s�`����Y\�~�W�i��<@1��	*��$'^>����hS7§�]�����1����]��;�/2ju�aC��Q�� t��{A�ٱBs��}�5h�a?SQ���M���]z-:�d'���6⺙�g�M�,�Mx�?�׌�|V�$
���)�~&��TW<S� �]]'�5`�_Yy�K�D?s:��¼{�p5�sXnF}Gz�%C����=k;�!���߼�mm��R����f�8��0a2��٧j�':G͒�9u`���[�Yqj�|��$�f+ h{�T�!��!���,�3�:����6-���Hn����*�1Pa˕��Ԁ���%��L����/�96�XD����U��m�}��e$�f>?:s8v�� z;Ւ���j���;W�A~��:5�K�e�*��:����3�!Mb
!֥�̥T��V�P�?Fw��ft��c�o��/�F���y��L�3��Q���
v�A����C�zӁk��Ğs�_
��:���z����t��2h��gB��s/�uk@�����>�1m���Ԙl�:�|����1(Y@�Ak�F�-�� �+f�U�B[��>5�C�D��ȡ0��bPЈ�/;i�L��򷛴C*���[���EG��Q�O�c�(���6��W�56�}I��!%1��� �iߤ��x�Q~�-F#�c-�wC�Y��^��p;&�B� ����.S�<����\����g0����_�H�}�_��}�N�K|w���(`�0��}��%�k~`XՅR�{��.�܏�@�n�c��(
������ %��T��>�ϡ�9��8sD^7�
��Yj���CA\!>9D�1��\%��S���%�`������)�^��oX"�'�A�~,��ܲ��@�J�	�`�<�Yl�Va2��h�������f3�6,�x�c)5�@�)2t$.C�����{פ��n���@G/H-G ��U/�ȝ��i��PFmA�s�]QfZ�mp�ΧS���:r�@�m�Yr�"�����O���� �̌���F�l��'�5�,����m9N�F$�vʠ�Sz�r�w�&��2�X�9TE�����?u%�`��s\T��D���0#`;��K9/�z�����������������?��A�Ѓm��^�/\[��h	��!����/pseDѳu��SN8A�2@,�l���-?n�z�O��&�h���t� T���\���9"E�����{����{����9�PlU'�շ �OeA�v	2/k��:��J��<�4�r�!QG������ҝ46G� ���3Q�~x렗�D��%X����������e������p6�����8iT:7��"i��J���Y@@���,_~����:{(��M0s+.'>��/�E|['��4_W�4�������nt)��do�;e�D	�k����H����\b��7�Ob%��7���#��;�u��=S�SmM�Z�9�tݸi�Z��0g�FT:5�{{ۇųW
�{�qu̽\u�3V%�Mmc�V�GG6]�k!�N�@y�v�r��˫k6���[�W��_[��/��j�q�Ӽ~�!��PF�>�I��ϳ#V�f�:H?�Ш�`|�`I�����E�+;Π楟�5U�N3[p�@��!\VU��f��xe�9M�
��p����ڋ���w���E��ͬJ�<���t�SO�:�&EV�Ob�|����D�� �q|�����ٮ=Ȑa���^���f������������Y�! )-p����!���+�\u�����-��*�	6sK�5TV�{:��Z��C�d����JO�3.�[�R{��8���b�fp1ֱ���j�$2�4d���0�F�b��g
J_�5�V�CdR�e�ڨ�S�芘�aH=U��ъ��(haS�#t�w,�Q��+��c��|7Y�4L��l"�t��m0f�9����$����Bu4�#�7!3�N�>��h1�ƫ�����M�W%[X�'�b�!��5��O�e;��=����z+�g",�._A�\5 4�V:���!x!(�����-Ƀ&��O�|��(��zH����E��`sq�aH��i�$���2I�O�MD�1�n����M+[Wڒvo�}Q2���/�z5����J�m�F�=���sE'�Ⱜ;�(��KiMd:h��f=�V7��j�d�6A���K���^Ҕ�2S�� �mo��,���I̊,�
ui؞h�+�c�Ā����z�y��H6ǉ"~�����&�."�Y:lяV�r}�M���f.��=A�c�r�@�A�C��gҫї:�{H�],�xA^�Ti������TD��p����O��o�5���v��ܫ������Vb*�98�u7���_9ۻ��"�h͌���7�6k�gF����b�I�5c�;��%�x�{��,:w�Y�� 
�ʏ�ĘCg����(�?���m:7�v�\���B��ΒXvi�� �D�\
hw�(!L�'~/'��\�2m�}�a��Q"RC�V��Ec�]P�Sm�C��Jx��?9)x�#)Ҋ�&kދ���n�d�S�#��O�1R��K/PՕ4��,����r��)����P�-x��Ϲc�����;ln�:\!7�{��~ b`f��T�r�6R�2�;EKj{�jr��i��;o%8e$<Z^��X�e]�?�ד�BL��D����|<<�_�(�)�-L�, �G���%H�A�|ؐ��H*���ˀ��NЙ�|�8��O����.#.�� �j�(�;�|�-%�=�pU�C�ks�L��·���G���������<�Lš%�i K�5�C�ɯ{��db�NO�mk(���J̶���	C����+�l�� ���p9j��L�0].�9;z]E `�&w��rm� f��U%�_g��$H9�D{|Ц�h�mk=n��3�:�j���!
<7���m2��7��y���6�,�&�)��m���������]u�B�:}��c��Y�I���OB
L[M����՝Z112H�gp��IK{���e�xn[<M0���m�A�,P����}�1w�
}��pY���St3?�<1ߞ��
�$�ɵB�Î�BS¹d�Q��IR��֒aZ ���C��AC�j�G�d��s�
:ք'Z��+�U�܎�a�����s��y��+��UEdEU=a��!1js��C��+V4�A�{P��x#��9c��3%����������#p��^jJ$\>���A1��/�eb��r%T��}k'\�΍Fڲ��)YQ5�ZI�̅!��Tk745+����G�w��R�K���^zď f���F����PDM6Q��[�j>S��3Z�3'���5^0�I�[��ܽ����J�D�e��x]W�Aǂ!g����� ֱ�D�ƒK��-C�fE���Ol��>X�a�&Noi�y��0��<�>aiWi_��E��J7T�X0GR)Ngz�T*O��F?�B�v0}B��$I�`i7a?np`�� �kNe�gZ	�����;�/�ɴ�-��}�O�c �ʄ�I���L3+���٘0��|� Rw�x��
�J�Jc�;�lQѳ�'^��v�$r�� \-]QTY΃7���)>!��EN�a�g�����s���·"P�f�>.�f_���#5GATk���s��퍖t���	�����=�������}�m�T/Ԭ��^�wǢGë|F�핋v�������1��%S,�B[�}���Z[��;xf���F���M<!дyȭ
1�˕z��{����S��naH߂���H�ud�o�Q6��AS%�QA4�Bf(c�ts�&�\h�l��&�s E���fr�X植U�apߚ	�Ԕsٓ�G����#'y*v(�S���ņ%b�.��T�w���<Mg�ĩn��Y#�!pAgI)�5F�$���X�N�糧X�F�v�W-`x+zd��7���rS�/���*�.{-�K��QoG�, ](��A
1g4,�.x7y�K�B��B���*��02�;�Ү²��BS�f�B�j� CZ�y�3e��� �Gl���4Tѡ�={�M�ޠ%��P�J�g{�Ҟ��o�_�!�,}}_�$�d?���O���mn����M/�GAY���|�<ZIC;��m�;ǖ��00M�Gy�5��R��"���\��	G��
�4�	k#�	ܵ�Nh��[\{�1`���|�Ֆ>���R�g�*�ȤIN纑��7�!��)�Ҽ���i���|�5����8��U����z�ӒtÖ#!8�՗zB�H�i���?�5��\��Y��p��	��a�2E��/K~�i� ������r�bM�ol?��N�(֕hqi1)
�՘<p2Ly��ƅ)��|�gX
Jו2]�'�JM�U���[��0�x\'��<Ç!�woC*�q&�;���vP |ңT"ZƓ��~!��u�y�V Y恋��X����jj�(ש��&�/�g�Q����%&�.[/G<�O5)���'���q�H)R~��5�@qfwk�z?�Z�W[�W�a,���`.x̲�yw��d��F׼c�h>{���OQO��O�2 %ԘP�I�� ͢2�����r ���m@�V��]���%��ۥ�ӥ����1C�h��Z���.��`���G^�R-lk$1H�o��zA}������1�D3܄-�-Ũ j��.)-AE�$*�0�~�|eӍ�Yf*!V�'El�_��i�-�\9��+�E	u��5"w�T<f�贈�=h���aQz�O/>����w�7��biU�����3�Z���_w�(�+<�A�W��!�Ճ�֍7 /S&��h��������\$G��Y7S��+Û�-̩;f$��7�����+�diX'���u`�5���`�(�0}�t�H(M������yǷ1��Q���Y�ڃ�OC����v��!�z�h阄v��1b�AktU�%�곦��0� ;�n��>�T�]W���E������8��3᫭�
3?�|R���:�I��\Z�]ܕ�(%F��*$�cD!���:�3m��	܃�Ӂ�j�'�d�W[����L�g�g%��M?��W�^Y`�h]Ǟ-jƒ��/������8�vH<��Y.�OY���^�Q���s�ݶ�f��,/����%�B�g�癫�oGF�M�ڹB��/'J�H�:�tɠ�9�(�v).L�n���&�ch��,�U3ުv+��bL�҆�ɺ�P�1�N��
}G?|���S6���j6�'�QV�)&{���/����C7��Cs�fC�u �3��R|}�#c�w�RۃȨJ��瓀n;�N���%� ��a��ji��ч�����%k�^�nQm���5��l�>!к�)�M�� �X���t�͇�Te	�i42����}���o�'<����6[٠�=�`�������: ��9_6t�(���Cfew3�5����<\������;�0#=�(��:�� ۺ幬�������rk�&�v˳����E,2��w�P�ʅ���H fH�X�7�j?;����+�V��ߐj_��[�����_t�b���]2؝��+�.7�"+B�6bwű��+�}{1\܃/�w��6�kw�p��]Z�X��ĩ�No@ �!�4���.�ᐈb�8�ޡZ��Zy�]�orP�L��Ef�b�?	i	IZ�u@v\7G��\u ��h�I��ㄆ�́�p7��i��8x�&���� ��ƙ����2����ݲ;��v/�6�&��r�"���7����/��ɩ���N�yb� �a��J�D�66�{���m�:������2`��B��Չ�ʅ��&JGm=���'��+y�͌Y &뮳�`��8͒�<�4q-�f�����Id���$��乜�ϐ��?dr(=0�!n�D��f����˧{G��
f7�v:=I��c'ѩ�
q�����v�r�����/}�.��D6-��K��-}��˷I9- O�G��=c�W�G+�2�Rq[ɥ{I����t>�*A@hB��e=ϱv)7	�y�f����ۀ�ͽ�,�ٲ�E �� �hQ&��]_�έ��!�$�1���XxʴV���l��
��kod���Ij2M���Y�yeQ�Cz\qZ�PSEb"�~�m��uk�7�-�����/�,N�u �e�^�d�4�u)܅�Q	�U�
ڀ������Ui�'�N��/�w	����G��{,r%�[���Ψ�3ZhB&1G��4�Hc�؇S�P�F�c\� �AvQ}a��6�z$�N�iv�F�UG��3 ۀ��� r4�jy4/�,�
�^R3T�CuKR����Z91w�&W�ԹF��A�M�ܪ�k��w�)�sD�H���VWoh࿺�Va��qK�I�W���Ƕ���J�1$�őΚ�VV�j,Uƺ���I�f�$^&���:��B$Fo��]{ ��Mũe_��~&p��3����a�k#�]�L������2�|�R�R�����a�b����[Zsە�9�O���*�����Ďb`��cD#N�Z�ਲ਼�x%"������F�N��%sz�����?^I��)�~�;�e���Ս��I�g��=�L",,��Q�q�'h�;�2X����1�7�!�H���.��I��f3)ъ��w�!Y;��5��~F_��}�ucq��4%����u�!�[��퓿�0��W�|�c��z��x6b3W��H�ʓ�V��8���q%.��ڛŰW������=�K|Α����Ae�}I��q���6�|Z�?��dd���Lə�n�@
��Rr����uc�Wj���o#�������l�)ouʦ| �Mo	��t�D�6,#�l��!�l�bDzS��Z����4�-��P�������:���0}�(d�l�+�^�B�t<��M�=�	�֑����yÛΥ<�4zևZ}dЯ[�3��u��ܲ��[��6�-�����᭣9Cʴbh�G_�~ (����>U*���D�r������#��? oF�zHF�����ᩮoP%�V&�˙���\�(�|���-��P��l��I#s-�"n�o~���Uo��/��i��Q4t5R�ў�+��"��z�Y�Nd�E塜�_��z��c&��q���q�>^yo�C���az?G&�SH���#D)ȃ$ep}qV�ЃF���M!S��n� �c�ũ}}����U�	����ݝ����_�؆7j���J��~�10S����(���$�=�!�n��x��wn�R�*�ȡ�
�#b]8���>��|��@8��sg�)E��+Oa�sP�I���}�eY��8�Y�{rn+�������R��6:��.;^Vgo��C����O��p:�2�:M��H/7Ҡ�╸�a%;�����u�@�.� ���B*�l$����	FfwdA�:b�`m��Q���s���%�h�`E��&��'��߆��fh�M7�����q���s%�d��z�	����Fa�1���\B�]O� c,%<�	\�9��wGI�k^�#��X���0����n�$�)�rYs���?�񗬖�V��5�U�7?�
=@����&�8�A+���N�N����R���_,:CY�����Q�k-�y�\�S�bx^��%:���'Ѿ�R�B����&3��=��5!�����V�x)�`�;�ٌ������s\&����K?�m*��/�z��xu�mn�D˯�_�SO��=d�Jp)Squ��*eC�M��¹#6Mf�1d�H�(�U-����"��:��?�X���5/�￭>K�Ie���Nd�$��.���gT��?�2� r�<�3Fs��1Ғ�۩�w��R���<y�(��()!<� AbmG��>�5j&Wu�m����Ų�_{&��	�2#hA�������Z���U��w��E�@8<�^e�T���tp�5=�_II��I�?�{k4u��W򙚰�iCqZ�<u٧"��?�f8���C?KA;�X.���5�oV=���I�*p�Y����6#���x�w6�M�-ǔB�#��8�JO����\܄�MD�C�vv6����ۂ��P�igv2ԥ�s��/c���z�Y����>�sUB�h�o���$*��֞�	��<�8��R�K�9U��/�� `�}\=C��E�y1����]��P���Ґ��i�hxZ��2e�H	.�H� �����%�m��'h`�R�;�)W����֑j�Љڮ�����ܤ'�db�����_��'΄�^�/�Gy�����ӗk;�(��M��/���٣����"^M�E^�)>�{[F��|Ǫ%���	��dD�E�W��{�=��f�F�v�ӊܚ�n9_�M�Ő���?�v�m�q2Ɔ�R�fWV!')#�װ��s_���Y����<'�D�����~���g]�&z��D
����]��2}�]�#��?�[K�(�,ݾ+rg��WߔS� �`<���Z�4����R,F��`�J�٘��*��&v�O�#FJv�5��k�J�]\`Y��b)nr�!=���y�N����ޣ�����y���� �[�OQ#�����`�U�,YL1��Ŋ*��Y�:�,��]�30��$;�M��<*��9JNHyc�����w]z��>U;F(���EkS�������w��4�J���1h�q�t�n���Yj�)�ϲH�(���]�;і��
fv�_I���j��%�6T�x<6X��%�U�M�(���V/c�fOh����f���=7���	�����<�\���v�v��~��E�>�1v�J�0�9@��CX�l,�}��&s ?���A4o����B��<���&���V$vM��̜a!�_+���L�������`�઒�*��S�� �͌�.DE��?��
�����<��"<�#��dh�`��J���eG��c�m >�� H�zg����@�n��3-����F�A�䮏C�4l�y�G9hV�-΅���� �f�?�I��U'N乌4�	N�"8dU�,�J��!��Ҹa"	��I�dv�{j��F�������k��Q����1��ޙ�F�&�zP�dv.N�G��Ą�n�r.���	�6�B`h�J��&l�#F�zG�S����׭
�܀u�x$�%�����Ք�W�����<�������{�Ƥ��p����Sa�r�Sp(�d�i�
��;�9�B��#g��tD���wЎ�ҳ4Jh�P�3���N� ��j��Ւ�Y�f��_����+��z�Z���S�i��<�R��~j��\���`�vݐ	���O;��Z�@��j5�����$d?v�9���Ħ�3/�����d��KW�XYx!gb��=�� ��+3��~	�UW}7��G��#y��
�l��-��� �+�7׭�k�^�AUw#rü�{a ��:!%��ۮO�s��4[���VNSIYMm�"�)��~:���^��w�IL_��k�Zv=�@N�U �B��S���q(�>(��|�{\�	o/��λ��90k���t��ʴ�{�n�5��E�5��JK&�F�����z4p��;%�@�e�dC���#��X��0�|B8���tc�������isXR9�@��חo.=��='��24�y4w�Sl�Q���^���P>ӻFI���6��Дꢊ[f���s�r=��=c�%�lc�,���i4�\�xr4�[7s�L�ZzQ=4�M\H=��{Đ�f�;���U�p-qK=�(�.�ᑝ��@�4��d���1�*x5xG�i�o t=}iH�Q'��~k�$���t��,_A��:y����s�����U��G�QBN�3*O�*�x�CxL�!�=c���Bq��9����Y��J�Ts�� \3b���E�z{\���;�9���i
��g���O.J������g"e����ʪ
����T:��nKY� :���0��"�Ǡ5�)�K K��n*1���GP�H�K��ecQ��#,{��&��HCD�B@�.	�A�;d/��4�����pJ�����Kz��y>.�fc�8`����Sq�)+�v	������&���&�4Ƨ����U�3k��䲽i<�'�%���k������)��蔲��)$�@�{ٴ�Ù�K1�l'6HO��E�k%OD�V^{��8��}��1����R��or��N��#1���S� ��(D��J��=dcedk���)�Š񋄵ӣ�?QȱX���xx��F��Űm�4K���\��Z`
F�ygy Z��8L,��=�i�>���zǣ�OHL��o@'xo�z5@�E	�}'eg����0Y��4����x�r�(=���i=��R����l��р,�:]�}5���W�@T�J��Mh�{
8������.���׃%e w[��ro\"�`/��0�	�V��^?����<wQGM�$ea'��
��W�M}�� MFd5���BP�@:�_V�1Ϳ���2�m�������_tA�XYh��<.�� MK�1E��Z/�c&@�,�i��Zņo		��l�1�V��`�M��� ��~���(�Ce�,�8�����͕n��u�S*�"�F�N�J�,4ٯ�QHA�cʅ�=o V�ci��vϣ�x��~�9�aE%��k*W����<�mJ|��A05��l7�c<�ݴ8�t&�F��~in�+<+�Vt�
����+G��w��!��pMl�Q�;,y4p��V�Y&��d�u�ֲMʼ�?x��w<�jem����D���Ȣ��Ql�M6��ŕ�;�W&>庮���e��GOeu�R�Z���~Dr:�����9�(��yR�i���
W�l�Z���ƭ���X7f��j�\/u�P����5���i���A0���}%�p$Q���_崹t�_�w�
�&.%1��8�8��"9!��z������^w	 ��$U^�Rm�*��·9S
�Ӗ��r[s�|Sy�����N�J�K[}��dL�7M"������8��=W5�YI;}+IY	rJ��έV�#b,�����Ҙlʲ��,���*y�ҰcN;c��銟(���RG��k��7!%�?~X��A&%��:�������N댒��w�{����9����T�] r&��5�Q�.�u<��\,n�X��������ǵ�K��3y����kB�.^=�A���m�+���/T�
��@Yds��n�2�O�}�T��v2��s^�F^]-�j�ǉ�w�+Q��aVm6����m���]�B��-n��V�'G�
`��O��/#�0�2���SP*_�6����~z��Oł�@�*	&Z	H�<c���$�^SĪqǲ,Rv\��kQ�ɥ���`H���=�3fZ�YEs�X&T�t��
�M�(���L�����glΚ��}�>��� �n�k�D�ba��ġK]f�b��A�O��](��˶}c�"�T�R�G��[�F���^�c�xѧ�l�X馴��s��D�C/,�K����=�s�ǡǘƉ#�Olŏ�3�O�`:c��2'][����}B�_�Kr�]ߵg	�\ۚ
��
Sb����)����$ݍ�PGH����L* ��kv>���E�@btuqGV0-��;�Kq�G����&�~ٻ�����c2�	Di�� �7��ƾ$��<���[r��������mi��H�o^o��'=��l9G��@[��&��WǢv=��]�\(K�Q�4I�ک	�?�y#� ���SBij��i�6����az(���a ����8�\�Q�Y��ߎ�a4%�&��L�
�I���b���H4�4�g��[ܐ�i��x��䨸�B:���B��w"+2�f��d����2��G��3q<���WB�_���*
�c!�>Eָ��qCt�����軹x�ke�Ґ.e?�)����Љjs�u�O��\�Z^m�ˢ��&��P��Q	���+�y%j`+h5��=��g�?��`;�u¿����A���Y׌�)�P����zlg�����'���-��c-�}y�E�h_���(�Z��Ņ��� �0z���'j�G~��y���z�EIZ���'ݔjN/�F�}��6c
�y�GK2�S���cQ���'���L�ϦIW��Cp%-�����ù ��Ѫ�35I��,Y�d�}E��6#x�X�8��| a):�=o�Ě�#�����!�f���0�=��iv;TE�=q�����toC��M�nh䮴�%3��W�F���t�Y*(������ӡ��lVD.-ZT��C�j5�lc��B�B���F%���&19��ٵ��
bE�^�$p�Ѿ|O��dc�{�z�2�6�c�3�n�mo�*~8]��%��p����PfQcT�].XVq��'k������}k	f�^	xW= [ZIic
]	oЬ�����V����'�JL$�b�X���AA��BA?yy+(9�sJg_UwA]�ª{�\Ȱ�J��+<���Ɔਮh���OuΟ4�;�]�A��y��2w3
Ȣ�5����[�|�A q�C�s���/�ƤϰƱ���%g*��f@7����݊xfְ�G^��<����������n�Al^�J^cR��`g"5u��A9"Ph�pbkc�A;�Pn�/�x>��.jnؠ{;D[��6?���kM��Ӫ�)@"��2�'�Z�Y�;�{��d.�A�<�Q�AJ�0�:�� �Ł�s�M��wgx�� J�ݙU<��9壂�Gڕ(<e�?j5�́��cO
�@ �;��qx.�郿�oD*xG��i.c] ��W{�q+���ʟN7���w��7�k����zS��W
�*h����3�O5#n^B ��Z�$c�?@�}%w˕uP>�n׽Ux�c�#�Ce��.ή�l�63$Y�ZKk��fl����bq���(� �ǭ���<� �S
LzLGw� ^��W٫�1�N�Ӎ��(Х�/�xyf��g�a�S:|b���N¨�"����G�Ϗؤ_��5(�֣���б���� 5�Os���4ȃD���$�I=�"JJ!����O�[���s9�5D�ϰ�	3��fH��纓F���Fp�����;�=�n��ܮ��(����"����ͽ��ie5j�3{� �+럔'��>-W`���ǽTV���[$�=����]/��<"���t �r�J�H+L�f�B�r���ʆV�M0�Ɉ�� iDS�j��(9W�Z�G�s4�7A�`R�V�H��u%�)����3�6��L��?�u�/U��+�$5[���M"��E�G���?>,Jt�+�'�FT�OuU
=c���~�w�����
p_����JH�ՙ������k~�,ir���3Y�5~ǡ{�`��CW������=%�1l&iY�A��:"~B�I�5
� �A��r�7%�9���U�i��ㅕ�Ps<e�t�_P!�u>�|����<#��V�<�c�w7��W8-�[�Cn��uQ3���<<�|�bo��.R^���)=�����/<�����(�\�|6S�&wְV��BP����Z����:q�.�H'`�oK	[Q�o��(F."��R?ٵU�փm!ƺ��3��62om����0g�x����K�2�������?vH@��f��&���	&̘�Vͥpʏ����+ �dゾ�h��U���$�+�[��e���[Fu��X���9��y��J��V�N�ϥ�tS���/�ƶR?��G�]hYY3f���y���h ,�1�p���//���?��k+��\������%_���-̩�&����b�|�!���p�CJl�"��m8�:�y�44�" �7�r,�ۙe*r�}���R��3�J�C.ӯ�d�bKܮ�:���㳤~��ވ�D4du������(�o��JK�.�WpC�k���\Wi���0�@�o��(���e��gEb�+��M�̓v:���Ne�k�
�;,�|�XK��:��?��nQB�F^s��T%��������w.8�N��99���9���=c�`yhz1$EH���aȣ���~ 1*���K�?uv�U~��?(c���>HYچ�0�(:��d��2NR	���J#��j��;�!��v�$�9-�x�����7��(Xk͓�Z��g�O�N���.�,������'����Ns�+j���>����L���LB�����C����⦓�=��Q<���qE�70��m��U�����Q!5�V#=�=�{� �{�v���Clfd��;��0�����b�H �����d�IW��A��e�Ue��P������5�����G�oMb����	�8��o�5kM�޴�D����PG��XE��C ��)HI�a2�6�IP@�V>�4�����s=�^�{���V7�4�{���3�ZͤB
[*��jF=���Y�a��¸��t��U�jE,��j߀�Ъ�b
贚_4�KSy�ZqC���,9^ĭ?b8$�}��!���RUc4X��<
�̾�����L7���N�&Sd@hHI��	Y����e�ya���aX.�SC9k�F�3�����(Z�<rF	�)�*�?8.H�Miظ�d�~��}&��8˰���{��//� 7,~鋮��ό���ڿ��q#1 1mN
����!P�u��!~\�&
o��K�s63f?T��7Tt�fJ�����a�wC��������N�?rB-�pA��L����+P [	�v㶓��}�ވ�UK4�*�/a��I���-s�mn�3���#s�|��)�OH��5W�C��Ɯ��x��M�9�5l-E��5JV�~�qa�c��}��7|G��K�#����	t0O��-$ib�\"- �T�nImN)�s	����Cjsa蒮�\�$�UPyu�M8C䣛v6��eX�Rx�Tݬ_�]\;����Ɩ<_���8�����4��vN�K��Q?�E��o���f��k�� �7ą���tX����O��l�:tV:ҬS`<���GM�&���p�иP�W�-�ALY�����+�xNzȥ����=�H�Y�Z�V#�������Dk}����������!��^��ͅ��&�J�%�mlP��������:S�m�^��8h�aL R�pZ�q2�$"
-�8�^����	������0c&��Dc��M��鬩RQ.m��<+:��(�D���2�L�NC�UD����x���T��~|䵂�'�t6��.j�����g�)R���FX�r�
r)����YA�cG͚3��8�!�/#��V�&`���c�/��%nv4�:z�.�	|�/���jԅ�q��#�o��by����J%��N�Jm+'v����3�o=�EW�Ja�ߢ"jC?��D?L]>톌��Ȕ�{d��xޥ4��V �N��9!x�
��02I�_by�����?׵���V.A��~�䳟_dc������qw�U+pB��7��
�(P����T"�,¯��L��՜}Y^��)��6������O٣��q���3�Ju�	{�g����3����0�2��O���є����!�/L���)���*�Y�,D�숼�驕v��I��G�$1RU���]��n
|�F1�4+�$NME~�R���U�	[WvΓuF���y�������p�sӬ�BBU �tdw�"ݔ��r��lOm�w(���-���Yi�}�QY,Z�7�p��Ug�߻�N����c��Q> ���B2���7�>��bq�ٶX��(승ƣ�Ze�Sf����1V�\�;����k�a*�Nv|��r�s��|fY��Pf�U!��=lܢ�-c��z���:� �5�[�p���R��W�*±S��],d��Y�C���7U13>�*����/����L�K�c5k��0��s�Y�ő>���mă�Q$G�ĵ=���*N���F��Q���G_��d�9������������.��K���)$oU=��{�����