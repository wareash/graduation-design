��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jåا{�\�u�?߷�dn@6�zf��r������;�&��0�#�8���V��F��(�I~%Y��O4�L�*��u�|��M@�C4����	�EIa���e6�Pq���������'7E6փQ�q�Ȳ ,󎶑�2M��v)���Ή5���Rk3.��/�un]��S���Qk����rs�h���>1��Fe��o������!6 7Ŋ/>����혹�/�\>e�+��x�7�;C�
[8����{��f���"�r��,��ٖ:�@�����|=o�1L��36��2���?<F9��5����E�x��%�����܏%�y��?M5x��7�e��j��H��HBc���\�҂OI���i��L��_J�X�؅(�Ց�z侕߻�I{钜?���E,	K�b�G�d�?V�Ѐ�t�[�Phĝ�A�Q�����RKw��{>8��+:���/�����[V�����;ξ������z���Ha����+Q���ՙ�LF顃T���2�������F<C��I���흦���8�����!qR������#<��M�k�0i;մ�$ʀ���ESk� �[�s��?ȯWv�E�[f%IqKw��n	�}��(@:1�f��!���Y��\'bn�oK�̩vf��"��ߚ �#KY��C�	H��ssױ� #4L:�(���=I��?�Z��ӆ�$�E�@��(�	�q����+���oR�'�psV�˰�t�4^�B��K!�|�V��%~"�? A��y�&�(���rv!���ف��^'���6����s�P~AOr����	���B���&-�O:~%k4�-͍?��J.���F�2W��T�\CR�rRۀ�9t��`'λ���ݎ��4qY4F�w��G��2R�nFr�\�+�_�w>%�H0����u!���$�qE���~]��G��<F���̿�����O}�T�+ ұ�8f�T_�٫�E�
T�Q���7R�.L� j߸�T'���v� �WYҡKy�:�T4�;�g�¦�ԬICyYϏ0"��X�14o�H�TD-��E{�D�O�U�@�3�l�jߍ�o�"�@z�4�9�@Q)��C��b��+�P�&�5�� ��̅�M}�G\e��L�1�xf��|�X��)J���*����w
�6�|�*��7�HY����?�w���c�V��-��
�H]�d��^���ʋ��1�y?"$�&����Y��"����T�.�WIfE��:�#��A�Kn��-�js%�/0�˱�](]c@L��X�t 7�����H���-���|���낿����hI�����w�9���Ty�����vK�|h�@�!�U�J��U��B⤇�e_�7E3bU��ɢ
� ��k$DĘ �o+�����}*JvQa�Ho7.�w�����/f�T�����Pd�(nAL��z�8ŷϋYD�
M�Xˣ�� ���潳!)u>���_x�t��7�3M�8?��h�)�Ņ;����&8�,��|`���$+�\ER�"SaR�������iF�݌�NYc_����k�j?^�A~"�-���(3	.N�Wx߶�f������q7k�$'�Ι�n���\\����+��_�;ztώ��Lٿupk$�c�5�F��
D3Y����_zh���"7��]��Å߈�sq�D������X*�>�Y,I#Xa����_]��񸸰W7�-VϤ�3ed�z��r����M�pϚ(�+�~�	(nFU�p��y����6��tY`k7�)�К�\�s�I�:�|-T��k��ө+/�GW��� x�6Y�� ���%�ب߀T'6ߑ��t���|@v���	���gT_�r�tu��{���"ds�Ͱm)������V�	րF��&�^r��qyqS��ae��t�I�2��)�{�|����'JN�)�o�-z�����,
���}joa�t��{6���d��|:�xT�J�G*�F|�'3y`*0�^4k���R"�-����t����8B4�������o�ʳx���8�� 4�7���n�����ހ�E¼�7�²�o�[��7&g�VݎXz��'�b�9P��7nk����|$}3�r���Q�CА��Dk<�q��]�����
�z'�wJ��߻�ڛ�I��8�&J�e2�G�������j�t�@��*�^@R��g7� ���st���f�Ù����yϞ���9���]8����l��I�X�<t�˗�V˄(�FP.m:ݮN�,_;��6Ea��x����Uc�/kJ���_<�Љ�#��Dh�a$)�#��C�To�����hv*�B�ֆ��,�=�_��4
�(>_p�gI��&��=0�~L��R�l�WW�8�>�����g�\� r�d�0f�H�yi,bմ�6�(q7݁Aa������:	�/��U�}��Ӷ@�Di��	2`����u{��~޲/L�u�n�ؤ>���W�u��S�_l�*yo%�(�*5-�Eq�l��5��ZZ���雂u�``[jך�[��w��������fkg2V��������8���{�[�b
���L
 ������a�ܰ�5����]gE�&�,ԼW>�B�8�֓
�RB�:��&��\�;�(qͩ���e�]�+�Ӕ����̯snL�����X��)����y�	����z
4k`H--��RdL灖�""�o�;�R[
�,$���wȶ����C�+]�;�Vms`UW$:�SN3#���ݦ��Rd��d�p�{��F�G�(�c�*���������O 6���p!���ݡ;��-�!RԴ3g�s���w�T�v�dIMǇ6��w*�3��J?B�m���vqL"�ؽ���� ����z�#p/o�wtE����YO�:$P�؇<qz*��]�9ðW��X4Tx+	eM5����� �O1,�3��<X,����%�?)����=J�]	'�<%�.XP9L1��$�'����{�>-.�����|�� ����|�K��\^X>�]�\�/]5�XEfm���A���n	��VI��"��ԪH�Œ`Rc����"�dm�"a�
J{�������{~��!� �	����
�/�CO�A;w�F+�'
��u/v��Dq9�ay6U�Њ�z��O GLc:������q��������05���Oώ�����O��n~�
�xLU�iv���s���&=�C�|��Ak��T�Kr�
.47�'���/�FA��ӄq	s]a߯��٭"eM��Q�u���.����n3���M��� jp�+�F�C�v����Qڋ#3�T4ԝ#�>��a۾��z����}�1�Q�aΜ6��м���u�Ƌ�D��ݟ�7Y��o������Cp�3�A�Nk�!ן��s4W�E���z�{	v����� <SIV#')~ɧf��CN��wې͓_4���0穸>/h=�V�O��b�΄"F�����]j�{��A���<�R�&��Mg���2np훭�:�:q�N��ʡ:c���g�h�#�+�_)fy�m���2=E^�7�Y�,p�aɔ�6�4�B�Z���8���g~W�(|�����%�.���qsaB��|���0���f7�ʮ�:Y����m5�C�&��!���~�%Y�xՍL�,쑃NB�K�0��+ۆ1J=qWPC�7��-L�R4��P�2�5�y'�c �x��^�Ҁ�2�9Z!�Ee�+���K�A��5����8��,�3�V�`��3V��H}`<]H.$(���T�l��&�L�� '����l'�OvV���ԁ6�-e��Ӂf�����W	{5ɼ�ޙ׆7�5�'
O�ٞ�=-gF̧���)�ډY��M�t$��gW��=J��ԫD��؋u��NU��|Vp
��̆�)��82�&��kC�ݜ+ 几�هFSq���Mb@���Y�Z@�NA��Jr��4W��e�v�@�_ٌ)�Q��.��sR&[f�1I9�K�MB�"�����nP�A����(>_4���@���V��ؐ�9E��?�"��>7�+;�x�Jtu�at������$<��u޼��v���[�0Em��II�J���|�H�30JM�(B��R��R��cݯo������|���[6+�\0@�&�P!�� u�wZ�eT�VH�H��y�w���?j5��),Y"�@���i�.u�/ދ;�0M'Q�'q��۟V�NG�JN���u���h���H
Y��U�/�~o0,�v4	�f���=��2� �L�ٙ�LzF��%��>Nԋ����Q �.�E����ìY�XO�Gq'�.�j���1EއV�/K�:r�������$?��� 1I��N2^&���6�G�ϱ���)��w���#u��d箰X��)4�{f���}�I�R%�20����A� ���d���r�ި��Ys�~��Q#�4��69Е��g�i�:3+/��R���uU�����0�8��^)V�� �:WD)Gը4��	Qݞ�1bڴ�Z}�A�V$�?��T��L�Kw|��A�*v�n� 7ہ�<���Cܗ�G�;��/��;�k����|]:~� �ߧ�wu���@0v��o^��Y�.�*��~FPr������������w����"'��<IP廏�I�."n�Wv�ߍz��K����� ��ř���
�,���ܞ��-uH����M�Uζŋ�H��>T �(Om�-�P�B��9Q@h7��q�.�m����PEg*�ī������!�<��t�_a�%�ۜB=��\�������"M�F��n��ģ+�\-���ա�,=�+к���$2�ټ��PJ6h>�t"�n���c�x��IF"���C�%p�8~�]�}�l�;��&���\e)2͇YI�^5���ZG�-+ń��%I�8���uKO�u�l����ڽL�N�o�~:�o[=ѭ���4�@�X�W�O�=���:)������dÿ������pq�Grv�1���e�*20�@!�� %�sݎ&��Wh��EB�ρ��#�XL}���ag��<0k��(�>�1�T$O�P2���m%\s���]�u,��BOL�io�K[F",�c'��a2�#~.,�w&��O9H��s�F*�Q���v{GJ�M���G���H0��K1��9��5�"����W}�"�RLF��M�^�f�������	�2�Av�Һ�]�fz�f��aA����C���(����$%-���h5���;��9.��� `v���E�YZt@�ZT ��Z�M�$~�)B��۩��W�l օ��C�єb�Q_?��m���5�2$'���EM��dڣ���vC�ul�̍'�S�]ͫ�iԫ�s_P�}eW����?�HW��
0 U|�3=�����+���/S�yu^�J�װb>�1�1G�W�����n���6i5�8V:!@->�^����L���8�+G���
��y:K����՚�_@������vğwU�/����ױ���P֗2�J�K��>פ�[��� �V�r�lm���CE#�~��C��	r
�,m[Q��J��4����7*��;^����ǓI����W??珹EESU�������>)�BO�@�A���/E`����9��)YFi� 	�F��ޢ�e��C2��������Ψ%�K��<�s+E��Kbvg+2�x�N�Q>妣�<��� �rw#ݍ��P���h�D�U�o�����zZ���3���D�q0<Q�E�d[v�s
���=�XL~�\�*H�W�+�����s"}�mX�-Q�� �\�θAgԇ����LY��Q	�#>��??+�v�4i�]�¿�lD��R�k��'g�Q6�"=�w�x�Fѳ�WM�C�~�����;I���B0�.a`�����*��X:�Pq��e@a�������RH��s�V6s�5D����K�c��)VA?`���U�6Y*B|��a{ wq�����6��re��WsC����vN��d
�KM��`:�Aܸ 7���(��~v�敜|���fĐ@i�NCc<M�W�//�G���aG���X&�d��l�ǂ��=N�8�]��f5K�S9KV���Eh	뿷4�zF8�c�o|����{S0�Zn���\�����U9�lu3i��K`�z� ����_���F_Sn6:�ߙ"���rP�PS�"C{��^A;N�6��v9�����	�O?8��L����G+�%$�C��C{'�ڙyo�n(��)s�J��t����k�* ��%�h}*��"]ہ�T<���.PR�K�B��*�>�\���j�zT�8��f�U��gB$�7�շ�
# ��H��L�錛����Җ�-���X���9�N�tr�{���ґ����������w1��h=Ş��$~�=���3�� a�����o�j�a��U=�����O6�357F7񮧷����613<�>7.�⌀ �J5���It�L5ۦ��TNI�n{�z5�"��J$��m�\���l��b��@m]<κ~�d[��ڿ:�Sk�X�T��n=�~"��U5�������A�{�����&�G��!w<���<���W]q����`�W��+�����wG�������u��-��R@�\�	��]u����.ʍ���u0(��V3O�w\�~�L�A%0���e�[�[��k�J�eGu���_�|Uio� �IB3�2
�1n�IF���[|.�cw����l�So�~�UP6q�q:� Ai��o�K��Nys�cİ.�	߽oOt|pG��-�e�R�QL\���+Ѐ��![�pf��VBN0�JZ��'n�_�+IM��o�ѩ�W�&=83�����s��ң4
E��Ϫ�h��G��s`��/�̱p3�C�:zV]�Ý�<b�����'�Tb1?��f�UKހ��S�l�s�^�����9~%}�+-k'];���]�u��7l�kv��K$\�u٧M=��KU0�4w�ܩ��:��2��{�G��(ٗ�XC�Z�5��¡U8ոޅ���9�j�-77��5���`]�Rp�<���H����I,p��v&d��)�J�o'2_۴Mf���^&^�T,�U� �k�
��,�fj��������0���&��d�����`���И�<Wv ���\Z��
�X�����kC �j9��}��{��*�����S���N�&��1����P��I���;�~P��b��N�~cJ}0.o�ԭ�,��(�5��,�o�Vc�ZP��|�m���Sp3_����Bp�:�ȭ���^S&���/���o��[�����~�C�P8��m�)4]wUܷ;Q�hC��~� ���bSe�r���D��E�ǃ���G_	P&���#�����i$���s����S�d#�x�� v���^�H�\��'��������H<[{Yp���$E�n�?E>����F��坣ކ��Ѧ!���g��è�:b]:��L��(]������)@g�8K�����/�t�ա8�QY23j�H M�i��m Ė$��35 v�t�IK�z_��EcKA�[�C�,s�l*�\gDx8YA~(*
�;����v*j�]Qs�=�� =re[?��ɠ���8̴rrP�5�O��P:�QtH6����7S�Ka��k
&�Mӟb�pG���ӽ.`��s�]5b��Y -��H�ֲi��'��H�L/�*��㳟� �9��[|�%"�.��[��Κ=;��s�-�D@���U��d��f�n�W��z�c��uf��YMs#����n�2R�~u�z29�2B:D?b�뫘"I"OMܯ[�"����� ��J���=��Đk<�{Y�Uڿ�j�IBQzv������,&,Ml�Y?�����8���ЯѨ'=�����b �H�Ƭh��̞���#Za\;sC�ۋGV��.�,J%adJ�,