��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e����d���f{��@����S��>���4{��ת�AO�Q{���ָ o=9�}�2�o�V�/,��d��#l���ؚd6x�����şL~Z�]A�j�8bi����q����6�lu�g�կP5Ջ�*��=��,���y�������g����@����CFjkҟ��&���7r�4n���N�w6��`3Q�R�g�˙H�|��+q�%�/i,��I{�Tڇ��'�q��!l�Ǭ"� �F��	�u,����ѫ��)?��ۃ9pl֬/afm U�*��[��� ;+���HO�	�^뿓��Z��q=ӣ��Kѕ�p���d�t�!PJ��dZ��I�/k�� 5Qo���Yt����0��'o�{�_�=�s���e�z�JȱY����6V/��DD�*a;T���ؑ?���G�a.ї����)?���/�q���?��|�VC�p��lɗ�rSm7n���ν�֮�`�����㜦e��1��H�\Ie���B�\}VN�,z�5O��4w��~rQ����D��Ͷgbezh�&��Mp��R�Zg9��׉�A!}{o���k����"��/�xW��NB%������U��`р9C>� ��<g�O��F^�|l��0�զ�W��5�l�i�s�fi�پdk�{�^Ĺ��r�Ϩ0�]�%M�� �Ӿ��k\��ܐ3��~���k�������uNH�MM���ٗK�9,�T��%�ƾ@�7�W=̲�`R���K�w�����В8*y��P�5x��pO�GR��`���(e���cPD� 9�wG�ٸ/����g% _̠tKN��N�}�%TN�a�x��L��t�(����"�".�;��r*բF�g_.�������c-C�{Vq�=��U۝q��
�_Ʒ�R�����?�7N��N*3),%D��*���l#����<ʄ�0������+��%J������$Z^l���!uX��/���]Q&��A�Bo	X�b_�&@��?c�^��)\�Xz�YNҤ�"5Kڜ�lw�,C� fZG�c{�w	�����,�+�g<��`M��f~���=S�.K��|�z� �Ob���cǋ�G���"�!�P��4��n3�Tc	�֒65tE�I�Y(��5�}�Rq�oy�e5�����D.PKK�/��������6[�졔��g2F�^�ꮙmZ��!_��������=��i�X�ŵ�\��k�� ���9�N�v�'��e3�@�2�x4=	������hg!S=v���"h����[.~�c�����O����ÛlFd���dǾq��d��NJc�}�'T�̀�w�yɂ'_N�Y�PI\��ɫ������;TG���r��|����1"�Ũ`B���{�pY�=����<�@�7Lȭ9c���%o�C����5��3Ȱ������4K����k �=��bw��]fA��4!ȌiR�P�M՞�圓``0��p��mcĔ��{�fF�f� ���P��@bP�d��G#�%�b�
[�э!}{@�_C���`�~�P,9�3$�Ӻ�R�HG45|�,�ޛ����d����j�%+8:�Zu�g�n�%os�w�_�Q;�46Q�i�jU%�W|��y=��0R�L��S��.�^.mĦ��l�$�\r�ÃdR���_��B\�S�5�|Z"�v�$ԳH��J`�i�Q&(��)�K �I�6>Rc�𪌬�����ŮǕ����L�$�**�@��W�^�\)�sdĳj��Mid����`�R�� O��H��&���S�1�&R�9�����������7XA��GP�Fu=��\�x��k
��g�]����,��� Brä���ȿ��Ӑ=�VF]���rd��X[7���Q���B�5��.f���^Jj��F~P4U�~��ԀO0��B3���C���,�3G@3]eϦ|;�.٧��R@��$-�cXmY>;�g��P�p���֛~58�2"l��?<����Ԫl�-���ߋ}��A��݀�9��b0�9�M���a������8����]�YM��>]7�$�\U�KX�n*ĩ.�P'|L�3��� ��T�#oe,X���\�R>������[�\y��E���(c会��8��^ P,�]��	�J�@we��{hh�!:�X����7��QB �?�:�Aq^�v�r�F�^�L�^�\��^]c�����
�ٞӘo�纒1'ۏ��c��q�g4း�(�b�ǆWS2���<ܮ�,x����Ҩ�t�4%8$�#�:��R�;ٽ3ıL-oD��k��H���ˍ�|�H�gs�y� "��K��[V�hJ7��OkL}�/*zY ր(^�\?�$e���tw���	خE��9,*R������ȵ;�8���v�vΘx8"XI��ņ�\��F(�]n){=`����x�W^�D.?X8"C!���,��']�N����Cr��s��s���2�M��u���Ī�Ð-ِS�t�C���Z�h�=S�ͼS�\��i4���f�C�Џ,���8���T{��k����[��F�t���?/���<��
��pX�l'�\�� 7�+�n��*z{���݇5��0KF�`���H ����s��t�,�0�ejzy��57D�l�=*H��Dp��Ŧ~!����	|w�1�*��@�N#�R2�$���m`x�X����m�Y�q�R^-F�K���v��>���D��yܨ�Z�����9����P�
A�զ��]���R�Q�b*�|
�j�Ac3�U��Ac=ڽ�r^(���,	�VD`�RĬ�)�kqxk�w���߆�)o���P"���'eV3����/��I�AC�~�#��]o*�CMm�ry����خyvYy�r4�v/�-H�P���!��0��u/дcB��kZ�0%�Z���p?i�G�y^�D��gTL�y�\*{�;Ø~2��ZW-W�~Mjtr��G�Ȱq��a#�O��+
�$��z��i���#DX�	���ŧ,I��b�.#�:U�I�m2fJ����su�P��襛�g�6$�I.��`��!
"�(�o*'2}I�M�j��;_͐���uj�@� ���cЈr§�s|ݳ�C!)�cGo��'Ф�[X��se�A���P9k9_7�ٛn'˼~��$0ߚ(x����H��J"��I��6)}��m�P�W���@ǽ�8�T��(�gg}����}2A�;]���G�I��b���I��-��4l��"��0pY-I�b�Mc_��dd�����}L��ȸ��j�-TI��}]��{��Y���	'�<L�/y"D��^��Y����4�-x�!ǋ�ے}d���N��vmU�ݣ�AO��?�2Z�`i=6 ܬV0�߆Vsؒ'߬0
��Pd�q��i`w��C��)"�p*B*݄��e�3x����Z;��6�Xr�O<T�5�G*	���P�wy�6_,V3�Z=�~^�Y;6����N��~6~I�����o��-��ʡ���k2��줥�UÍm�abL����`��4Ʒ!���pX[�%�B�H	�`�]��/#Cqek�m��-�n\IN�`�]�����ݶqxpq��&|ͨNd gK�EVx���1��g1���NJF��	=T�ڱp��Ӫ��X��?��g�CN�EX��n��X{���5J��ف�*�Y�S		�:g�<��s�k�ڑ�n����+�׶�<�N�#[#A����\����M!��s�khk��t� �v4��?>q�V,`�z�7q}Q3҈���k>%D8=��F�j���y��:���a�Ҏ#�ַ7�в��3��Z`�<����y�U� �賴���eu$��|3D!�A�F��f*���?��E�T����>}Zi��!m��DQy���9Q_(�R��])��O�,�,X��Q���1v?Z-���;J��ٙ�ZBGж�E�!9xIn}$�"u�	� ���q��eJ<x�8��٨��AzW�:x@Jg��^�oA	�fz��R �K�P9���λ��sY��$��V�ڨ��_�գ�,�F14�_�0V\��WB?������@����j �⁉z���Dp���a8���Z�G�\Z�Ɓ�q����m��B�;E�w����Bٲ�Ix�|<Y����p���5�ހ��)N�˩`��OVc2��4�0�%{B#^r���RϬRm��	�y���-�k�b�� �x�x7�ܷ��`�c���[?�0T�K�m�WVe�t�"?3,L�{�o��,��.2�|�X�a��Ȩ��k?f�H�Q��N�<�Z:)����js�}5O�2�UN{[��!�T"�R	�}x��ڝ�2�(T9���r������f1�N�^-���̧|����A��O� 8.]���`���ʟ����r�p�Y�Z	��͸��������#N��g�  ���K�S�6������:\v�9f_��t��p���!ۃ+��ܤ�}ےcV���<|��|�-]ʃ�z4�$��W+-�EK�0�1�?�6X�L��JP���S�|O��OJ&��!�?��k���4M�c��zu�^f�]�Z�y�p�{I�U��K�5G��W�cA#/��6����Z�z�|�\,���'��������G�8 r�y�1m�/H�uY9�����B�
���Y� ZL���)���s[�ֱ�yP;�K��ԆE�)�޾�!�$�\hU��6Ӂ	5��f*�v�-��<p#b4�I��Y3�ի0��P@�;��+ĄNW��`���(4�'������
�y��L��9s"ť���;���̍�ڍt�I�u�2���+I}�|t�lY�k�x=�;%$��5:����*�>0�M�e� �z#�FLQ.UV�7��|��mgr�o�W�ч̦��nn������7�1��x� �9�T�-=R��d�N������w�r�E.g�ɭQܜ^(�MS��kM�{���3��:V�����18MvP��� ڀC;^����Z?�%j q�i��?,��S5������L��߁U՘����N}_��>g0K�{�\��=uFzǪ^���DY��+�$�qp��o����H?�-���N��ڟ��֓`��*�`�mS��R�pϜ���%I���[k�=MD��(ުa�s�{�L�t3gVp8�p��y�$�� ���W�|5{��8�� Wh��N���V�/,�"gj�D�[���8ڊ�7V�k��z��}�����S�K��k�Wg:���ڕ�aĐ��!]k�P-�7�7�]T�DOZ�2��~u���a���D��!"$_E�5H��t�J��{L~�5>Ņ�=�B��^�ʖ��eas��`(/ǋI��LЗߤ�QCw��5���oW�ի�}P1��k�-��ߝe$��e�nM�}��N/��)�<��~i���;_�$�5Z$�6S,��SQ�V'��ʰ�{v=�u��`xH��s��l�P��wK��H��OK|��Nkz��-��48�)�,��2.��ּ�s�6�>P9l���M<a��׭���}I�U���2 :Q���0�G�d�î���Hϻ2f,5�ڎ�D�͏)������a& a�k�:q��ƞhÆ6���*ڕ�e�P"/�"O'�>�\%Ν���i׽O�������FQ�x�/��d����[�D�"S�;�;���${�j�*o��,�7Kf#��׼.';��/�7�Ǒ�m�� z�S�b86�@0z�G㔒M�t����J[\����r7�#��������hrv���Yr�q������:��l�/'��7UJ����ǫ��6��ZX�]�B����b=g�e�f�������w�cu��<(@��5���:�r����tYT��ǋ���*~1z)o�Ι"�F���{�d���޶�^.�YsG�?5cY�a�aE��I����7�w6�7��o0g�x����Gِ���NZהu1j���y��lFӂ@)|��ŅS������a��Y�O���6ɭ/-!�	�*����_t�&� '�*���X�8���1�I�}<|\MRc#)2�iM]@0.WLqd��r��E�PR��^�Nd-�§Z�E<ZYa��ٷHF�IO������.�fĩP���=Y����*�#��1��Qm4b�<���O&������h@�ϗ<5i��Xݸ]�K�Ԝ��F�3^ud#,P��1C[UT$}xsS������7i�s�WI(o���gq��e�RB��_��>���]��7uCd�'��~Oc�p<�T�kq�#�p.�R���ְk$��G�eL	������ň9)A*�@ �,y�tu^��'�S���	�$�^⹔�%c���.= �H�C|���z
��8ْ��x�&{�9|y��ߔNϔ|��%�uO?ܝ�N��5A=o'k�[���1
`����z��>������dZ�Ϯ]}2zz�0Iq�B�p���7!}����w�p��l�3c�>�L��f����G�&�����e���3��.{\1ϐ��8��H�i��.�O��ִK�T�;eң�S�����:��ͼ�:��5YE ��O�+�o�mbm*�2��+f&������N�:X��ӸnE!�d�m�_x���l�D>*�RG��`y{�ר&U���p^�7��tY�D�ye퍌�ĩ#(M��ϕH�?��X�Q���.����[�W�>�$ �(���q�x}�,{�sf���/��T�|�����fy��/�P�=Z��e���p�n�`<�G`��"���pսQnڄ���h]i�����S:Cu�%�T��6������U�Ǭ��$L���;��ޱ 1)0�E���PGt����h�n`�!����T�I95Q|ͨ��L��\�|\�/07��z;F�n|�I*� �2.�1q���kZ~�-eUNk�觷o�OEW�mޅ^�d���r�3�lYq�t֌fZ5򮍟d0���~6��֭ ���Sg�N�n�aP����=� X�=sCKw�9��_��Q�fM�W�e��T��X0��&�)��doG�2�܊&�N�NSR�Ba4t��Cp���q��AZ&�2�����w#��M���g@:��4(+�/=F@n,4\^��-!}@WO��`��ݻ>ɔ�Z��w��F�b�^�F|�r�^;uh(D��� �ՋU���o���e�rUD_��E�Zj�U�#����L1�/E�x��j@�
��le�-2�lT�!���A�l�@�++�b
��0/�u�;́����w
�yXA��R���p"��3ą��15�6�zf�2S�^5։~x��F �z��^vO�×Xw0꛻�h��R%)�?�1��)�#��R��p��\�b=�f��ݲ��;@��J�&��vv�Ld�$��$�c8��~�+6g��P��D%���yIj��SW�~��3Rk@ɭYO��g0U����>��gu)���Ջ�@(�Ŀ�Nm���	��`JM]���P�G��F�m�ǽz���'ô�kX.ξ2���[d�qS-��ɶՍ*{�����K\J�� &���A������[��6���>-��^]'ʧ@0���b���dj������E쌋�r>��T	ΓL�'�%�+�����/�����:^�8��uUҷ��ɶ+Ze�������c(oC|?TfA��7�� �luo� �X�H%������Q�ٖ�Y7h�n��9�h8/NF���{g��3}';���Crׄ������X��ϔn�\3iN�P4��}X�P��G(�N��\����J���c�9]=5����t�t?ާ�O�l���+�ҫ���Z�e�+�q��� �uzm�#��ږ�m���Tռ�@;bԙ�˂��q5���il�|׭/��X�(`����]��B�7�_r��ޫ�vP��}�"���S_�Eou�2j�5gF��
�"�Ğ�1��z@��h�ɘ�&֒�D���\ɳ{PSq�c!��*�o� 7k&�[.����X��XƺQyj�@���v1��L6�0/k�{�,@NՎR� d�ms��L�#�o���D�\�#�=�990�G<.A�J�qa"�5�q��A�,vU)�k�����ޠ����?�q�$U	�)m��������zn>`�S�X�'�e��������ŋ�{�@��t[�g)�Wz�E��MЕ�z����`���jmcj���B���7ӄe���.�[��zUx�M�Ь������O�V��u��:�����JKh~Þ	�j%h/�!��ɾ_A��l�R�X��?���A�x��s�u
�*��K���ѠBjZ�{O�����B��liC�xQ�����,ŤH���(K��, i ��F$'��)�Fn�e�m�qR���#�Qg�� W
E!8ˁ���d��)ZH���Cz�J����_�`p�8��)>0�:��_�L�eP�X~%&^a"EJ�p��ù�3+���C����ؿ�K���w7DӀb��ԃbϏry����ѕ�u�Zց]M>շZp_�SU�z�孂��M��3���A��|��S?|�t����O�0qCC&��"��<�Iͩ�;惧�{�c���/'��<}Z��-^�S20ҲV���T�w�"��ƽx[��J��6N�Z�j�3x�pcV��˷+�P~��n_5 9�k5��,��{!��8*�}�����t}�ı�rD���sP�?�Op�	�`�Tۣ�Z��ȱ�]ٺ���n5�n���i���G(Y�X�\(&����N�P�����j�VA�cΒ�C��b3����������6bNj6�<q �L�%��K�������,��H��n�X(96~"Ί����� ��a�	1����~>7�C���#�,Jq�Ԏ-i}K�f�K���=���F^9�ݣ�T�ι}���2<��;��O)Ư��������2�j�f(�=�������A��߰�j��Nw�'Uu�2���EE�n�.�E�D�0�3��8>��	��j�w�7�O8�z�	eۯ���˻�!���=ZY^S�<:����d�i�!�����w�Cx:���9>|Wn���5vZw�`�����y���v�v�в�[Ď�e	^7lI�jޓ��R@Dx��Jq��B��S7� �f"�3��oer��84ַ�m'�_J*s:��ghe�31��*&%�et���I�(F~���(Y)عjOih��8Mb�pa ���5C�br<���Uk�%ؖ߉��8c�Y}U��G�#�xiUmEgď�����c���A������d-�t*�.'`�I�J���l#�R�!���6�ʺ��S�r�l�ۚ������@='�/�{`H~�GW��%�E|���fC�fndu��Ӱ��e�7��G�(����q*�P<u����~���2��w�E?̶8"uN��W8�?kO�(C@��;,n��/�%kf`8��jǆQ�X�[T"���u�Cl�M����"�� ��y�<n�/Ή�����\g�@��J~�q
�G�I>��Ca�}Y�z�j�����<�[2	e�������f�A�������lٺ6?��D��&�ٞJl��T�][HB7��$�J�nX��ȣ_zt�o�nN�Z"�b�	=���;CPk���P��o^���a7f���0��^hr6�L��W�z�q�1zX`Mb5�<ᵑ�G�~6e|���(��"K:��u��^4@N��؂_ϦXk�OYGCƫ����ŧ6���� X��ӌ��(���꥔�k�ev���W�4{�6���,ڮ�6�u�����|9�C>�]�����խM$��v<xf�,@<��|zqo�i�IF��א7�^��
#�n�
� ��j�"� ��8.:H���~"�ؓ�k6&�Հ<�p"ex\ �@���E���t���~�ߝE8�"�TR�L��=Eȭ �7X�[k� O%�Ĉi��R<��D�8��|9�3�o�L��#���0�NPn���G*H5����4����")�A�NQ|i�X�']3}���pf8Y�߅���ex�b�V��%�X�=#m1�̟�T�tx�c拻�5'ql�g���}9�x�A�F�#i҅����eM��1��;v!�y �Q�2I���#$��`�j�U$���%JXA��H�д�?w�	N^���s���*U�ᣆ@�b��7EK��CvT��+=���@VB�=�Sv�8�]�����u�*5��f/Ӭl���L1���������|Y��.v��e�lQ�%NO��I�v����M�%j�T�OS�n=֌�8R8�Uf��*)!淠��RF���N�z��Ҡ��9n�D���;��}x�K/U�}W�H!��.���V®\B�����k�׏!�]٪��@R���&��HM�I��k60~H�0
q22x�)�AE[�"���CB��P�>��a�����2�M
����b��G��8�@G�r������=�,��Xs@e�X9�`{��5r���5vF���g1�n�	,ڍC��Yb
��Y߅ѡ�Y�=�c'����X@�Bo �1�cn�ʆ! ��n��gY���=8�":h��/����f��?���@YiZ�Q��<AlT<�ź�o�Z@���mi���X���� �Dh"�� �`w�2e��oHN�@tA��w����Vc[�e���	E���C�s�H���;r�Xܦ������[��o��O��w�>EqpK<��B����uJŲ�ȗD�f�,�I���;�tG��ta�Aa�y2ĭ����ė}��3I0R�:��j��[u��t�0Z�S۸����	��M������јo^>H3~��ܚ_��w_�m�����9��z����^��w��7��(��I-~��l��Kq�pB6���fC`�0g��H��j��l�l��Z���|����fe��Ɂ��R��Ol�vr�v���c4o9��G��t���*�M��	�v*�G�nHz{�K�-��ճ�ֲv���#8w ���/^v�w���d����1��c��15���H0�꨽����B�RJ�S����*��I`!|>�[S��S�����K�-QW�ZvXH�b�eˉ��l������Ϝ���2[�P���ކ']x�̢L\g~y>�}��4a��ю4?��,=Q�L�6�$wp��Tz�STG�>����7VM��ŭ,���K?��֖���˵��ؤ`��u>�&�jaK�+�V`������ɺJ$Dx`@��g��7İN���9����ճ���u��F<k�cfM�=�e�a�&+�Ac�I���@��՜��h�T��.��[f���z�}g��G`�{���|���#�a��F���&����El:\������4�v=��{c	�+	 93����4=0���]NG���F�}�W�4�����+RY�f�� ��ۛ�/��<\��R��P��s��L+��O��⦈���O���
��-i d<S͋lM�Q�	$A���rI��v=��w�|j��)v�8���O<u�~D�M�fk��ָ2[�^��U�}R�G-�_�V�ֵ�"�pw�{�-q��
s��6�X�X�.�p��w�3:�8L,uI��GY$%
%1��7j#�;�v�84Lɣ���A��Y Zg�A2����ox��^O��/�+�s�ӻ�\���2��g!@����}'bC_S=O^CPF�=,tJ�+E��Ώ�?y47���?,1%����Xxa:
<r�-/ʹ���U�q�;��_�x�m��E�Jp���G�6y�82��� !O�z�"�fj�*Q��-�������*���������Lѳ�ϛ`D)�T�b��H�Aި2���e�{��f��*0m�Ot�o1 �5
228U���!O��I��%fS�ml��/b�@3ހ^�m}���0��<�+q�h��yD��h����( j�+.&{�H�׳�n������.P��ˁv��b���e��hr�,�-��܆������*G�,�9��0��>ӥK%/vT]x��테A-Ҟ��ױ���k�1&mO��ST-����(�7�Cs㮛����,��߉�X0}^7-��ϑuX�atБQ�@[]���39��u��V�oh���0~�����[�P8Tj��h�l	~o�J�tD��Iv~=�L��Y�[j
����c��N���y�]-(�z�(��;#�&�c@��"ٍ45+Nu8�ML�*���^Om�KCZzLQUMլfj�u�k:��4xSH%[Ґ��
_�&,���!�d��[�D�����B�+<�ˮ�?�_��8+�)�*RQ�!H߄9�7$�H&���n���(�+ϥ'�?��ؖ��H��O���4Q��42���z!�t�o[�&�2m��)�|{�p!PCl�T}/7�&���0a@v���n�-��p�c��d�ܜ��ou	�׺0����9n�n\p����]��e7l��Q�=���.�4O�+u�j�D�^f@ ?�U1����7U�	l���%��6��H>�
���j�-�����[o�W;�X��n��X�%����}�-�u�I�c� ����̡̂�
��Kuoz#h2�&@"�{�Z��Z�V����!���c�T�B0�,��ِ��۟� Ncβ�0��.Z/މ?��<���N��nIg�ɇ��9v�5U�-��ߍׯE���_27s�)D�u/��0�:���ߊB��b��Oj%�񻎙ǗMF��ǟb�7�_5�1*�D�f�����:���?���W0��m!pyx��Z9�����-3�S�δ�`d���F�S�dT�7IWW��a7�Ę���7�S��|�*�;v?�Z���c=�=x�m��\��j+��a�׭�@�<Wy�,gY�b>���.��xs7�̪�e��؀�)����S�R�R&@�Z�)���s�Gs��JN}rO�O$����EX7��O֔��Pw��h��b��Ј�R
��ye��1Ϧ� �Z�j�y�5I�,�TtI1�vQ�Y����Ï���G��,����gaC�x��{�/�����<XF��;x��w;i�t(Oh�-":IH��`nK.�c����M!�F1���W�P�ψ�$��0X�����أ� ��¸�������1�Z�tp�Y���=�1��-gn�Ž�o�{��g`50��F1l��h7ڻ>˘�qy�K܎���Y ���I~[]���T-.:��]YN��b7dk�~<�Q�eXtܝ��B#���CA��3��`vڳ����P��!W��V�8�Q�e166,�3������DsR�<]��i����U�e2��$J��:S���ݱ酋��CG>��N!9�a2p�����z�P\���9��~ҕ�=��Н�O�M!=��i�'x���R&.z���|��sx�ױ�Z�3�'Т�I�ZY,.���ġZ��;~�z^����^��7��/8ZP���-�|�s C��?��JMΨf��˱���=@Za�,X�K��B~1��Z��0xX%�x�T�Go<��DE^g�g�B��JG��p?�P��F�w�s�A�D-
˜�K�:�WL��
�딚%d�����T�mJN�G�o�������>/O�@M����Ɛ�%�F�m��%�H-���U7ц'6�q�99��xy?F��fMb��r,/��Ǖ��0��6ɵ�p�=aK=JL('��'uC�������w,���M���?���4{�{%�H�H��5���x�#�c,�ԶZ��qW<ͳw����E@�c���(��g��'o���YH�d0U2�f�!��c%`�w�� �˫_LN������$�=�,΅�|\G�(3gb�5�){DTo�$����(<I#;p�7�`�p�_����"��#�a�n�z\��l}�xm���\S} ��=M�yk�R=��{���	������*0��˖��G�8�`I����fh�f�:��f�`%~���x�Э�Q�hVUxy�d��#8ݿ_ �Ce�� L-F	��_9d���l��Ġӿ�� �"�`�����Z躂�f^�׿T<�C3���V�Z�/m��*�B��fـ!��iZ �nZm����WԲb�DK�Z1�Xm���y�Ů:�-�s�=���vBR^mPM
�z(Ϯ���]���4��X��?	�r,� ��@���Ya�5c�d�����G�*m3�F�`��^M�<o$ty �:0��C~\2'|��]-�A��J��m;n�~uo$S�[zWm�ń�l}|�q b��x�	}R�%g8�UzL��`���_�4�Zku��*��9k���2?�/�*~��,�5@�uȺe�g�msd��݉3i��Bi`T�(Խ��_H�� �pݘ_�b`�j�4���1���`k@_|��~��H�;����D�j\���֍R� H=��w�u���.����M����Q����T���!��ǳ�D�ޣ������G.�r~�����h�\�+T��5CbG*���eͿ!�U/�Du���,�_�:k�z�����X��|�5��|��ǐ�8���1fD?i���|�m�B�r��n��rI?���%[���f(A��%
?Zn�N�5��YL�$���<*�����K�C�+�[0�fZ�v�6��T��2zQ���P��'qI~�i<�Ч�>�CD{W�6Jh��Y�}�5�7?`Z�q{p�� �4����X3�Dpb�ƶ��� �(m<��_ޜX|r�9�<��e��܇ɚ]�r�\�"&��b�N�^	gi� ��4{��i�τ��M��.�5�޾ъh�j�[)A�����@:�o2�T8hJ�2���ن2N����F8�mm�}1������tg �{!�QI"uE��`I �V�f㴜��ωK<{_k�_����гVij��*���*��.X��	4� �S.W�S�V���"��D	!*M��;Ɠ���I� 8�!��� x�M��QHCSqϊ������Ucvi�A/��d��ꦥ&�|m���؏h�5I8}�0Ɖ�ׯ*S�Vjh9�s:�ơ��J��EE�z�\̷mTT9o���s�M�
�fፏ�&r�x	�	��%yA����;�	�[�\�b)���q�%S�=H_�Zr��gS�p�f�!�iu�0�T�;����]�Tj�0������n�}�G�׉���{��Y��\����}��2y7j�'�H|\�2S�ȿ�3���l;��=�*��-�۞@��JƋ-���������ȥ��#�,!r~8Bd�RWkи�_F��p.�q2�b5��ͪ
?y�`�,gG ��l���i����(��T�>q��9�=��t��ik���nl���D3�fy{ΰ�	�\�:���čTf
v�*��@7hǴ
SsV�h;Z�sP&Y����fJQ�@o�$%�z�̇R�J���`�!�r�;!@��%a��ȵ�4=�r ��E����\9T{�hI��rjЫ����~�c��!�hJ��n�U�#�E�LW���[�0(��Ań�e�5Y)@*{�W�Y�踥R�z=�9n/Pi�8Nѭr=Ȥ��I��"�H2y"*dm���BpI�k�t�F����d�\C9�x�GC�L����{כ����*.F�B&�(4�>��Q�/v�k��ox�*uNoנjc�\�Q�ޥo{+��	���g�r�(d9�e����w���=������׆`=�]��lv����({e V���y��n-�8�&�\^)�o^v�a:�o/��t�r���P�5��$h~n}f2vx�U��l��\�4���m�x�ެ\���0g��z�
xQ��nύ��]�猑c� ��=�`{�qc��,�K��'���z���<��.����Z�Z=���2ǺT�${V�=v��`Nh����N�(1��R�%��3l���	���o��6�N��P�����턩^X���_�3�2;�s�J��-@��вl�&o�������֒��8Xň�0y�.�&+G�4�.4"��*@�{��zD���Izm�O^��)'���#��(3Q�:�'��+�Gtf"���
Ąd�����8�9���Z�C�S
��<5!ՙߞ��S�5�����>)���ߥ��T=��(Yh3�%^Uq8��J'��k�Sa��z���5���C>�ܹo��YfQ^Fyk2��6WR�f$�B��s����W>�2��5��2����ĭ�=i��	6s�=x}���2R5�[F�oU�z��n��<77��LN�!l𡃏�	�]�'*7�[�硴��ǁ��Om�* G~��&�
:�:���Tk��|W.���	1M���9��n��PU ��!�J���O�JtT<0��T��U��t�,w��E]���b���;[̽~��'�j }|�w����3 �X]�����oP[���м4�!�mB@�͘�	�@�]M6��!�6�S�om�fy�B�䍺���4Y��ŗ̖�O43�	���`��<�K�B�߹�
��)o��%T2A��a�w�!S
�ګ��@���;��m1p(�����0�S2���9,:pA�g`e��]���OX�mcНe��Q�K������Qk����.��g�������|xoB�'U�>��`G���8���wQ�cX5�ܻ��B�<p-ꊷl��FH��gm��ʥ�o�����4�q�i��e���
���!BP085p��'uZ&x!/o݇`d�5��c�9*���:���}'w�DE��x�@:tsb����������6a�gm���Y3�l�9�'�[eS����EᣑA�����_�:��G?��UO$�r3�.A,�#�w�z����s�2��P8O�r�}�us�T��n��l=<���ђ�/>�sJe���o1��mTЂ��h��}vei�q'ꈢ��V���Hb&
�
|5?�=PBl�v���%���Vh��UXJ�[���Ǡ(k�9��|X{�ȱ�i�;j�cs������Pk��q2�ᚡ�/ahȰ@L��mSU���(��Z�UGo�ؤ��|�)?8�f���u�$��3����f���1���ź#�3�? �C�@]`��7I��h�g�4!1/{���y�#�n��b�B��:�!�Q�J�6fM�����AP��~v�UA�w���
z���B}֜��A�g�p$��.p�>x�S��uf҂������U�,n���� ��K��ye�;ހ���{�l�������0�b������R�▏��\>դ��
x�[�㭥�0n�?,PLS�sZ�tο��ya�לy ������&U[�Jry �q"o2�Y��?�y0 &�vCb��\ާ�*É�T���[gvh�~���%d㢼�T1ƶ����u��n�Q�w~V��EgPR�W���2^�'�(�CI�d�b�s��}i|zz�"�G>�y�C� M��0�b_6�N��d�s<]�%U�����o���G�X�o�k^���������?�\)<څY��~���YD����*������gVT�@7Hm9�Eq��.�G��d��q���A�ؓX� "N��Sڴ�[�������A,bұHX�L�.dz��ݲ��!>$�ϳîC��Kܒ���- 2/����ȱ3#Vc�.��v����Z�5�����O�v�ղy���~��W���g���#� WIFA�X"\D.��#F- =;;I^�^-��M���V��WR��N�U�6���v���|D����ei�hW�1/��P�Y�Jp{��=-��xbV�kyD6�9�B��d���]&�A��~�ʍ۲�!�������.�Kޡ�x�"jV��cM��@a�����������Q��"A���=��Έ��2Do_�z�GG�bF��|@f��������߄-;.���Q���t����q��n����X�jn��Ȁq����0a��!J�R��<��oxDe��V���{�bo���`��j"ؤ
�]?��`kl���ٚ�<S�,mG~Ds�K���#�c�Q��O�"0
S��y�g����y��ʹ(���heĚ�Pu�u�7u�Kc�$��n���*�B��$3�����H�? v�W���=��e���5fE�f�k�H�U���}���̊�ƻ��0��ߨ#ua��@�S%��r?��%i�%8]��PZN�Yb?O�5��C��ˊ�d�T9:fV"�c7��
�kBQ~��"�N�V��
*��)m$���/����[�_�7Sh~{�䱪���h��r)�SL#_7�)V\:�_	x��f�G�rk�i�:b� ?<�����sug�

��s��B8�ҀV��K?ŋ�/vX�.�'�m���]h�h�".t�*�S��#0%µ)��O������oa�FF��!�{������%M����S	�v�'���{���e���D#�Lܚ�$/�r�jev�N"�
s�3Y��l�ӹؗ���ȘR趸g�F۹����E��K����`�C���) �`[���:Ky��j?��>��ױ?�S��e�1���@�ѶiQ.]9m��&�@$�\�!e�M?!��Wg��Pm4$%Y�w��I"�"�ǔ� ��<�t_�t�;��o4OB�-�� �+��Mi�bW'ҝ&?١Ur�l,�6"S�2r]ke&ɍ�k=�ǹ��K8{�,�{}�qs���&v�w80e�� �_ӟ����"6Gƛ����l��nt���^1���+3�����k|���	;%���V����H�fO-�+�	0;�<���>���~W'Z�%nz�J$�3��#��a!���әI�r�|���C!�w�$I ��ꔸ����cC8���}�:�-�E��0 M+ԥ6�-�'p}!�@�Cd��
y^ކ�2tn�ўY��*>Y<�q]5 �K&E�/x��D� #Xb�Z��|`�q���a����Oˈ�v:��܃ϛ�����\<v�`brb��F
-@A��9q��vA�N2{��p��g��u�W�tH�6�]l	r�_.���'����چ�P�x0(��<�O�_/q�*��8H���)���:?��̫�B���&�O����,~�����^����N	1[��\Z�\t�cLk��/����>���`T	Do��������r:�Ĺ�(���q	SI�d�
��Zdx:�`;:���Rt_ݸ{�^����q��q��y6!x��#{�g�IP���Y��NV����YQ��7:X�T`�He�v��
��������L�r�Ѭœ�v���P�����<��C~��Xqn���E��!<��S�W�~i 7�hn��*�ņK9���_�ަ����:S�"��;�ې��Pm�����:j;�	Q̬g�dޫ�>m�N�Ge�����4Zi7�Ӟx�KB�j!lR����?󳰠�
���'O �4�m޴s�`��K�$�;���b\���� ڏ�.�5�h��!��Yն�������fj�� �s\GpQ�����H��&���I�+V���x�e�s�9�;{��S��Z�C {�*���8�^��ɢ��@ٺ���k�|bks0��Į�e�k#�0c8���`S2�"�+�W �������1���W����_�"�4|�4�W���f�hK'���X��f�҇����B�3����L N%�j�@� ��Y�<���cεRߨ��W��F�W���M/) ��Z�5Jh��o��B 5'��@؃6�)SQ6����-�����00U}6	4�D�9����f?{gB��6M`��l����P��%B�i�Q�s�;Dv�[;�HI<.Z������瓪j�rU� ���_��l��%�L�d����OYxz?��R�4ȧ.?���bʱ���U��>��Sz�H���pQ�e-?t蔩�MJ�x�G������Y�,����i��
B4ר��!�l͒ �"�6� ���Pꤒ�K�1E�Hmy{�D���h���***˺IRn����S���7��H��uu��~`�����;<�x�)Oy�W�-���,��'���RJ��I�g��?'���E�ā�������B$���(�p6.{��<=���g��M���,a��!��S���۟:�*� �G^-?Gȝ��F5ۑ�*��&oZ|b���5Zm$�[�'�
W�&�L6�z�:΅0A��v� �%J�q�yC��BZ��|'@~Obt	�	�&A<�1&�S�fB�m��_�����u<���i2��I�}�tdתKI���@j�Ї%��b�h����(�3��Ef^�М���Ι��*���96�&87r��?0-�VO���L�)D'�q�8����{rY�c1��ڍ�IA�6'�9�,���K����w�N���Kk��4B��i��$���{Bb�$�e���| �mH[������tf�ȁ��a4]��W�{�d������%��{��+4O�<�
zc��2��'�M�^L��v?��/�A����oMyj��*�I��aZ+t	�re�u����8	���Pt���>�r�&��H��.JP�}�}��)K��);���v�8"�9��c�>|`�؆x�e�q���Κ�P�ˍ�=�|��IE�NL`YCG����C�3�R���Mb\́�Gx��F�#����=���v"��m�B�۰S�ԭQ�TLH}�3���\u,9���Q��|�6�i��!�a�]-F��/�!�=�V��]OU ��v���݇��`ݪ�[σ\�x�ob�x��}�cb�|-^O9���W�.�#^o$8(���df�7ǅ`������xwu��	��#�#!s���QI���-�:��Y��c�ό,�͞�u֡�p�?H��殸3�*�0*�˛�=Č\C<�8Vю/\�:�´�����^w�s��>�N�
$/�֑�}В��;�:��J[������d��9↉��ӎr΄���c��v|��+gxf�X역(G����*W$��X��2�w��Yr��m^�q�����).� ��s�v�ra���ߣA�{�¸�i>�u��E�,}���'��T�� c6h�+�K�L�˦+�v��I��YӖ�`C�k���K�oX��:�=���������I�Ʊ��Ύ�)��d�;�d�������CyTZ���c���/u�e$����!P�9��:������hMKr�f���1����nWGJ/����"h��wy	�2u���n��W&����P-`ȭH�6���U*����ёNU�mK!��C��\�h��60�ĢD2�i˪r�D]��?�+��I]����$>@��b��z���L�e9��Ib��ŞMaˇ��W�I̜XO_���,�,�:��鉙9������Ń�D1{t�+��M,��1&�íQ�.ˮ�T1Ϣ�"u��D6�b���e�8y�%i��gn�UȧL��L�2�#Ii��j�/l�I!�Ic�Ș|���A�G/ِ7��~����~�#��v����O�h ��*N�0�.zxR���A;��D��Xy� �����b-ί��D�b���vjG��!��-D�l���=Cğ�o׾e�.�x�c��"6�6j#��h�k�P��=�)�峅�:<ﺝ{h$���4���2�+�Kn����c�B�gRq��3/������R�+@O�@�ϙZV��l�j@�(6,Q�Ͱ4[y��>���Z�ӵ�S��$��[f�4�>�K���Px�(A�L�;4/��ܹ�����a"��  ���be�к�J������4��%��L�ƈ�d����.�P�V'w}�Ov?�Y���
�&L˖�d{�V�z&Ku��vp�b� Q�|�c�Zi�Lq2eX�i:|�)�} A�٨!G؉����h�_+��Y�|5���rgs��>��er��px wZ����v/y�T���HS1�;�k^{bJ��HJQ�$3��<K��3���.��I<&�R�S�㋃#/M��X��U�3�&���n�/�,�iw���cp���E��@��������&���C�諒Prjgg~�tt/�<�e�pg��5BM����7�B2�6S]h�n[p�����n�t�d4�����2��N�W��p�P��I�w��1P���c{�Ca��ī�[0��T�+-��Y>9��"/	ɕ'<�eN��-^��=��Z��3�#�	��箘�M �S@�KM~���zjO���a��?�᳐���P�UHa���kUpwye�k����6<FƯ�i���$��ñ{4	'�<�-uz*���h��!%��}�-a>h��6EH���m+�y�^YE�(�� �#l,�ʄZ��?~+]R5Z�u��4�����=L;O"������:΄,�����Sͪ�%	b�gzb��H��X�7H��[ѼA�`aiͷ�����./#H�U�C�I��0��9W@j	�?]w�3wġ�����Y3���p�ѡO=HD��I��*������>���2��w���E#�Xڵ�!s�2n���[���8�{�pjz���������׷HZƏW���e��wL��=�"װ�F�Q���m|�X� ���ԋG� �_��[2i�<%uU ���Oege�y,�� ڰU��J����9�>��H�y���3$���Sn�3����8�l�4V0ǒd�+|�Cʮ�{�oÀ~gsW��'��h���=��;���ew(��e�^�Sd{�Ðp5�y6)&�w>��S�{ٝq7G�B*(�k��h�\șq��S����/�~�n���R?�o$�P��[-ѽ��(4�rUʬR"�I� j�^#�%:u���}l>���t���z��گ�7t���z���k�y���A`�h������>Bq�-�Efi���H�y<G��
>9��R���S���~�*��˧y�&}����45�/R�Xq���.����4ؖGԱk��Y���6�2������tHV\��A��=}�uC�B}��G)Gu��B�"%*-��C̖�D.V)p`u�m4]���ZJS���@��m�kDＰHѥiK�1i!����Mj�`9p���S�.���b�Կ����T	՗ν1y	�|�x�q��q[�������:u�U��Ag!�����N9:�=��dr�]���3��/q(�e�����<������� �f1X�>���F�u,L�|初�7�o���h�!���D� @��$t�bʖ(t��T��k�%5,<x�S����'����O�x���(�θȌ��k1_L� ��An��Tε!)0���%<��D�>`�].\^�2\���\y`�|oϥ!PP�`"�%����$j��}�`ϻW�.1[B�����n�Q�"��F�e���+(��D�ζ# 29)=$	����ӿMm�j����]m��D�G<��%���Z,32P���j��5�۲L���A)�ԉ�V��|��m$�e�zUh����z>]�n���+�`f*䫡|�Mq�6݇X���K�.�}b�_����w�M���B�-'}嵫k�Ҩ�1�A�W��'%�G�Ȉ����|)���נ8�l��pl�����v�L3��Ƌ���3�~�c�r�W�d�`U��1.5@���G��D��N�n@1Ҍ\})@�5�"���c�ղ_��U"f'��0.*� ��򉠰k=~e�3����I����D"�p�b�����Z�-�d��K�戰�X�D��AP_�
t�g�`���
Ά
;W��s�W�˸��=`�+Z���+;��U��ְoH������0K#��$/7�_Z��J`�C��ĵ��F���q[i#�D�'��mwJl8�j�0e��jc����mUU���:�U�b8�sCy�s���L#�x�����d;<�P)��e�F�	��:u�u����D
�NJ4��-~�'�f�|m�>7�C���ً���)��*?�c��X�*����=�l0�YvrXf$8������6�,f�Xր���)TK���fpGi���?"_��4�Ogz�h���z�fN�s9h�F,������y�����L�^�㢅�聼�f0]���t2�~���e�ڧ�z9�c#È� ���:AKN��[���Pxec!wd�}Ge��/�@��pc$�-�� E,�j��%�A����H��L!�~�-1;��fUr����x%U���ն�� �%�[�k�06Cn")��iOTKu��r�U�	�t�t�����Q�%���r6;��z�!CxL,�R?�).�?;�P�`$��G�L��>�S5U�J��(��Z���c 	�@R�_~��Mv"��W�ܭ������7\��՟�C$�aZۑ�E��C�jC~����&�c�P�����y��&�/'>���Ӧ��VQ�44�+x�=_΁��W�~�N�@�5F��+S��9�>��2t�1t����)G6�f��$�J�T���7оJ��E;Ft�H�%�/�	�|�p-0$�_ >R�T����%��������3�\���B��2��:���gH �4]kxCJ�]��A���;�F��(){���%kb�R�n�l,�Dq&���&��q����gx�,̊\�����lU�{�g��o���3��h��)��4�a�R�<�G=y�q��J��ѬAW�r7M�g�$֥�2�`�P��a��U���:����tn,߾JD���U�9� ̽C3w|�z�3��鴆[\d��bG,g&��ED*d_�T��[���G�·����q��Vz��I�K�c�߷�TL'H�jU����ei��]Y8�_�Y8l���G��C.W����-w[�s�AaR���U��(�7��ʇR��a�3T.��ɚ��4-�,^����Y��/�x�ݝAG���}�)�����+h�/��B
���� �J���]4��'�%K�w7E0�}L��Z�8B�6|�uA�[�+��̗rA
 P{��ĝ!!4�9�K����-���\3�y��@)�Zd��i%�R+�����|t�-cw��u]p��܅d�uz�d�~�����]�=?>�γ?��Yp��x�j ""�n��%�0��Ь�H7���F���x<ֽ�d'L]_�T��pc׉�a7y�~ ��%��h�fW����Ҥq��\��}4C�;�R*��L��Y�R�d�f��K�	�Ֆr����6���T���Y�����*�����Ԧ{��F�e����[C0%�˾T�>I��|
�(�pPU͜Z�>�*rb$rs�A%hOL��1���Y`J�q\����h��&��$�0
Ij0��cLR�����5Mp)EI�G~To��,^�,!jb+��y߰^��m��:��2�U�=�4����3���Ռ��n��3j��/���\9��Il�GU�!=�ը�Dc`��z��w����q�ORw�aQ8����k��?ƷT��W��]?���^y+7,������g�'�����N�(a�|-[R���#�+	�-��w�����D�h��Y�ȅ~j�~U~��Unt�.�A-b��z�a�T�_+/{9�w�z�W1���\i��9  (C�ԣ�,�����̺W)cg�����9��r����>E���FͶ�翚�e���U���?��]W�wc���&�?��*����� xX���">Fɟ�mt���Ix��@Z�X8��묏��w7&I��s��%�|�����GZ�h~"�c�`
�{�o�]猑�`�,�ߪ��9��߇J���)꯺{	p8{R�GH�!%��f:��)��Z��;�Q�ǹoFV�g���0���*0D��[�x�d�͒c���	��ة��.?�k3 ����C�R�K�UGE-"v����9�x #���a���3�<&��@AQ:8U��௷Lߘ���ī��+j�Ui�Qj�<U�Ezu�ǲ9���ግ�'���E�w����Es�P��H�嘸����r�_�Q\�=x� �f�<C9\�Z�s:�
v�~�V3uKz�����u��<OĚ�=�}��h�|OE�/vFI�
X�6f�tY�qŻ�����H��'(o�p�L|V!V;�_�Ŧ_��}���7����0N�ˢ	��o��:�
;}3�؃��&r�ܸ��,���/�����*c۾�_͖���腱v��_T���Q�|��?�`�F��K�A}�fa���QW���?��N�UInX��s��
K�nn��?Ǖfص�B9e���|�Ԡ�Kp���.��5VI�~Љ�U C�<S�B�s�5�gl�b�F-�[`G�i"d���U���A��E]�vQ�Q_-Z~�~v�eU��q.~�*��.�䇥1���b,��R�������f����dt��$-Q|�@q�Jf=;jq79��gZ�qm��ۦ�,��Q�8\�y�q�EQ�?�e��@�hW�	j�V�,_'�YP��M�?��~��wg�m���`�e��?��2��#�4�A���[��7�w�]��:X�M� ~O�}���`���m�*����t, ��?��̻��	:�@H^�iv��S��]T�V��F?�=�t_	Y��"؍d�)��n*��}��#�������B�6bi�NE�t�7^�̆��򵑞0�(��Zt�m�C�ѼT����|ޣ�<����2��ݫ�ThjIH�Q��6�t���t�7�T������������@��.̑K�5�Q�9�Å���!��/�������������9k�������\E|�M~~�{h�0@����F�#��TRp�>��i���<��,�Z�o�(��y��!�ˊH�5%k�ε�8�t)�G.�Թ:s�P��W��l� ��w�}l9A�rg�����B��ӆa�����)iT��Ƿ�h�[ߠ'�v(���7�`efT�H.1�a���2šx�����pkD���>u����tRwȷ��]:yo�w�/�
�Fn�6���G2\eP��i���L�\r����7��������$��7�P�Ӛ���PdN����2��z��;�"����?q
��wL] z*���T2p�.K��Xͤlƀ���8霉=�g������d;!�\y%�&#����e���*q� ��#c��;��r�+�֥��>�#�Y���H�������[^����F����;0Uy�0/�/��c'|QK�"+�'�E����_(��:� _t����E�ˠ�P���<(��l�ξ��u����V��}���r �AG'�s��#Ê�/�6�A�9���^�F������ʚ�>����ڑ�|���Ba�����w�2E�^Խ��%2�?�,s�g�DYP�Bx,s��.)�e�G\�$�r釮7��?���"�i��9h�D��>D�F�O�iU-�c]� �X���ݸ���#�/�����F�.fD�"��:̙txC�����6=�FF5��\�KC&ֱ'b�b;��������w쒊��Pl�(c�4��K�xgd(�Z�����*�c�^p/H����2B7/���9�U����`�~����lS�i�VW�h��&�����f$ւ�,����5��N��8lM!�t/��L(as,���v�2��mp@�SC�s�6.m�Y������ҡD�a�T��ڿ�ha��7�-�����E���ta,�Λ+Q/O[�G���	j��#l�2a�ic�m�HM���Ը�CZ�~����¶�k?TLwR#ٵ�~��HeDY��O�/*Yo�ù:̌R��&�[W�w�)��t�7��d% '�o#�k#:�u�Y9u����xlo��Z%ah7Y_x�2L��޷�8��&HAw�޿V��

��_0I�sR l�� �ICB��ӄi1+�ʒ�y8�F)�p��H�.?��/�FC#���и?ﱓK�`��J�X�y�^kB��nۅ(Ot�3o%9C��*A�g�A�ޝ��� ��R${'O�d&�k��ԥ���M�g��<��b� �ԹG�g������(�_������rc+���웏�6͎j��"�e/z��ǌ��m*iS�PWNÝ�))`��m���?z�$k�^C%=�g�|	�Dj}��$=z=�<|� �L�I9?�P�aT�L^v���Q�djʋI�j��La��ԁsy��_�m��O�~�x�H�����wυd{�*�r�d!4S��� v������+�O ���&4��,i>[�����N����&�T\��r��Qa��7��m��0���-�a�L����fs-~��aӟ<d!ϗDnVsxN���!2��as��$�ܱ'�@|q���a�m�E�䆞�`�GZ#N��̑p��r�0��|�����z��J,� �w)fx)�m����w�~ז�Ū�������7�P'�h��5(���"��-� ���'��n$>
��G��7Zf��ע�u߰���K�ɛ7a���Җ�ξ`��)g( o��(~#�����*���ɨ粂rV��kҮ���:�E�Y��ߴ�.�`q�0�W�ӄ�]�X�@�~d�/��Rie�s����>J���Q��2�SH�J̻����+v�4�c7	;��gy�2��_�t���A~\	8������P)~���De�x2��t4�\2>4��˖G�(����e�O� L�'�x�s�h��
��!�z�Ʉ>}���8�$�\�i�ӕ"z����,$)-�����C�drU
��Ƌ��C�������Ă+�+�0���#(��� �W.�D�r�D+
��Z����N.��J��u�#11�s�@D{��֔R��)�	�e�A�� \/w����r�֍$ͳ�Ж`� 	F�OC(,Ø}���8aFw� D
�|]�@>k���l��}�'Q���(+��vѴ�K�f�Y��8��l�L"%��gٛ��:��x�)G9�r/K��="�\��i�D�P[E� �8��5�ݓЋ3�uҟ�����[�E�Qqo0����z_4=G�zJ+܃�U���I�.�9-�c�ɓ1�^)�e6[أ�n� �������d��U`�d�b��H2���$A��1KFP�,�	P�����/����w�vv��T�C
en�R�	��^$�1��h�_�R���O��5� ��dF��H,��}Gc+&$k&��O57���bp7��%�R4���ub�#�"{SOV$�N�V~PA�M���v���bK��<���&V���ҿ�?�J[�����9�M�2|�JϿ��i�3v��61�MT�5�Q��d"�\N�-"nP�K㓠h���؋�?�d�B+zq9�$�B�8���f�=��d3]���'^��>Zf���-;x�@�8W$Z�>�-X�s��<hh���{��Ɉg�+�iw������"n�
�V=��ͬR��� ��zH�r\S��ˍ׈9��w**&ݸ#|��x�7��2��)|�4k��{	�x��L�Г�ǇQ�k��na��>9E8E�9���n5�%�W��}�`Os��W՟�~X�̂�H��aQQ��C�/t�'�^X�ȑf��{�>����a���8;��Ʃm1�a��ѣnw)�A�^��>�{�zҵ&%��|�qi��+Qۂ���66���H��D$���6�1]�+�߂�px�R��0�QH�ii���S;Ȅ��2؂�ʕgc��2��n�K%���t���92CDG��>58�Or����-�
��1�x ���|F�u�lh�wĲ�Mg ݶ�@^�s�S���T�+�ȤIO��!��Th��U�L�-�����f�"M{	�.�x�ÄW�G"�$,�O�ty�KI72��;��"3�c9��|���"�mL$v�]K�b���N:�����D�4��q�&Gw�l��/�<�÷����
�6JdP�>6���	2��ǌ�R9B�|���Q�];x��n1I��9�@3G\�Β=���γ��Ǌ�d���䳭3fkJ�kk���{�{tI����0������Uy1�<��~9=R<�%�X�뺥�)�Gf ��H�!�O�C%�`@��Ĵ�V�`�U�[��2�Y�ؤH���V��i��	D�Ae���r��a��X��v���SucA�k�+JF3�:���}������/X�%}C���&K�`'�_q�'�!��J@ ���Hy$
� 6�ls��3��Ta��0��IeRhm�yNu~>�B��yࢰ��y%}��,5��z缛���Ma�}ǚ߭�{O��xS��6y2 bG�|җ��*�9F���$oU���q�Wpk��~�;j����bs�ղm�w3�#���K(���^9�+u�=��h��w] s`VO�UOis�tW��^+��H���
�����>���?�7a���N�$Z����в*�]EA�Ȯ
��8���&+Y��cnx��-d>�vFd��Mx����'_�O2k/�sE)�G�(�f�+���l�Qt�h�X����f��,��:6�nM����>W��4h�r���l�|���r�j�}MW�%�y�A:���	BF��>: Z?�DI=R���o�x��L<�#8�m��a�8�s�0�}��0���O�;�)���^����+���,+q�f=�-��,5IǕ-E�`=l�m�ok)6hx��/�M۹�k���H�jx��1��uQ��8T	�'�l�M)�6O2�����,�yiB	50��;���ܳ!����bz�4VIu�r�\�&�ы5�ު���cZ3�4�G���Y�RƆ���W��D���7}Vu)G)����+&H&mq�,��V�B �\�ZZm�U,+�n��=	 �>���{�Ԯ����"���밶���^73%���Q��Kt�H�Q�H!j�Rc�H�fm2V�מƣ���E
_���#�9�l:�4'�k��CaKb�kd�,���/�)e���/~[�|x�p*a�,slFK`.���P� S%�8~z]�]�pDTp[��ە[��V�>
����//����'}��	b		H�:��S�M�|���r.б�^_�ۙ�W�Z�1���F����'��E��qe"}�Y؆��݋R� (R�;����,l�ih�O��8rv��Y����ЕI��c�&1�O�Y�_a+bH��#${,�5�{}hͫ�����\����SB��Ju)a�ͅ,x�jt�fNҊ�0��(T�����"�na����.;kf�K6����¬�*��m�mf��gbl��ͮ�oJ��X�$<6��`-F�q����'�'_�i���mtI��[��JJ�]�Bm|@����+
]�)�?�%5��	�\��b\���(��+�?��*�@�-��4\��7ꀏ;��� ��[�w@":&.>�-ߟ�|��T����2N�w�Ҿ�Ѿ���t�Y���ސ�f?�D�cb�HbV�Ŀ�{$�h��ϛ�,&1#��H嫗*�[k�x�ì�6��!�����l�+K���{����F�4g��E-��F�p(��zܐ��Vb2��zy��R��O����\a���ӂ�V^�v>��|�y����t�$Az!�
�΂}}+�0
tkJtr������wsTҙ�Q��	�Jr�}6Z�E�7��ؘ��v&v���ڸ�D��^X=��[9S�#�CH���)�y�+���}���������G��6�6�y�R���S=����ϠQi��,��Af��y",_>���� ���;g���C�����|U�T����l�x [�@�Ґ��)�3OrZN(�o�-�x�D��x��W���V�S�}��6�����% �VB[��xQE׏���Rl�'��+aS�T�o��6L�\7���H!��2�7��!"�2����L�mzـ�l���߫v����(TE7	s)DB���@K1��IQ�*sĵ{��볨�Б*��ՀZ�#��6P.����EM
չ}���
Cb��t����yc���$��$��K��1�f¬�}�[G��p�%��� � ˋ�J6���VӔ*�kmP!�ǆ^MLF�ޜ3���τ��R��&=U־�-HE���w
oy��s���N�R��7�dO;x�|�H.�"A|:��z��=cL>���|�,�/:�RE�����\�pP��+Y1tO�#���1ܮ�j�L��5�Fr�^"8;NpI��]mv�k��P�
AP���Y�r�e��"eWR�l�p0����_>�&g���5��'���o��V�����zb6��4�������tW�T�p�4g�{W/�~�#!p꽉�3Y�-�0R͉�VR3�Y��yr`jZ��
�O] ��cR�t�^Y�Pي��B~2;vi+eT.��|1�!ǻ�@ �J����xF��p��dQ9x��W�=�8�g�Ӂ$$���m��^u�DF$�oL8�GU+�i�BD��Bom�J	�N"�Z���
�����ב��\�~�U8���r����i\\hV^z�>�[rŊL�Lt�����?̹Qw��	&7����w����:�w�M����!�H�Dv�a;�I-��/]�T�\A[�'&�o�إx{�I�.`�u��������%W��:o.�����Ո��U�4�Ǐ�i&bt)*��6�ZW�*@�j-}�8�Sk#�\�`����!痢�m��j��UǶ_�&�W$"]-ә ����X��":�.+	�� G%�!$*�G���ȍ�<�(A/��u�n�M�#>��xr�s΀���@ ����g����
�甕#Q���P���}�6��Ft�QB�R���oP��
pr���ϳ�@�;g+j�
-s�+���8���c�WSL5co������	��j�6� ?D���&���HP|Y1E'Cgg,�Pӯ�(hoLs/���2�x0=�|A�n��Ҍ��	�B�*�-�x,��Y�a��,��
wtG���V���=2I����4��ۭ��Νu��x^�D5�K�r�>�t�D�0���_��d���p��n���n��I��\�y�ǒv��l"�_��4r����a���w˹��TBP�h���L����o�u� Z�4�%�qZ�[<��"Zep<�Z'���������X���pܥnB� �4����&X���/�h��N�&��+ʫo�.T&i��J�Hhe�ň�\>�ގ����?�5DTͯ��H2���\�$ċ.���d����#uT|��!=��7�O\���� ��2V��O�x9qLԦ#2qUPeT���j�����Y��QkU0Й�b�34���|��/8b;�����Q*U�O��~<�TE�\�R��r�m�������E��r��I���р��!�;�H�x5���ݻ�ڝ��Ȓ�7�z	�+Mi�� 'դ�(�������H b8�F5��܋�3
�9�l��G�1����Oe^I���.���
:+\h��8�,k�b��@��YB�o0"%�)-*�"uH�(��\���T|��-&��D4���"D��l��B�B��e �O���9#�Ot³m�2����.)#I����"([��YpY�]�K������ �m
���	�<�����9�R%.�ګϣ���i3PS�O"~|!�Us��/��,����K ҍ���1���f�[� }� �|�&l1���`��L�a�b)�QR I���k�2��0�I�0�*[h�d�OR3^]�� 7/r�ɋ���r�}B~�ThS�Zn�aky��w���m��W`��H�N�V�)���c�Rp��̰E�]�y،�䍼��� �d����bq��,dÍJ������Ds��V����C+�zzܕl�����_��Y�H&(hؒ���L��N�k}�����zF:�&%�aq �8�A�!�~�J�K��yJ@�zc�cR���/RI��M<��G�ODa���{A�!��5��l��z��N2c/ B��<%�Y<��>�0x`��|F&Sh#Z�������v0<���7wk��TBsc�eKH���C	nM�A0�l�&�F��B�y)��'��Pl���{�L+�|���*�+3���^�l=*�Uc�~#�v��3��Sg��b�{�>�{���@#�����5�����c���^uK;N�3"�*5h":�H$���2;�w����s�a����fs�>�X�1���`ᯀ����̘���(����������5��?�:;������h󬉲�{���o�� �'��FK����W8?٬55��w%�44)���hm����@&-P��g�|:~�
�:&'�be�%km'ߔi>B1чD�Y��d�$�;��^����xD������u<�)�r�g�C�8A��wy�*zA���m�ӂ�$��$'s���A,;��
�+'I����?����`�e�P�4u`����Mt�L Ҳo�.]l�J�(Vɝ*#)��
$�ԺC����mk�9��T�i<�}+�O�K��(7�Z�S��R�7L�k�"�Ñ��Ez����<\9��u��S4�n���/f.�zb�9�A�h��`�Ə?l���� ��0C���P��z9�P~���V����p�XDC��y�]���0���-�U���m�@|WJڳ��/��ky���/[��z�7��/x��J��Y��K�[������$��z�._X�pA�������MMU{%m_
��+�����b�(\B�&X��&шkL�XD�h��x�}d��Jx�	�Jt��yAσ����'P���4r�)r��!tU�HFtز���@x�����}�R����߲cwv�2���IX"�]��A�*��0���u8w�m��~F]4�IC��)�댒���u���)?*u���y��Ho��ˇ�c:��`�,۔;�94����>�ƴs��鱃R��;����/��^���>�̖;e.����n���~���<�6���X��
}��c��Oa	/���s�^�١
�J��s�&��-u�*�J���Ǥ}�9�8�+�PYE��mG�1&Ƽ'���mA�+c�%=n���z���3 ���7]G̦�߬���{�S�His�GCo�m��zy�&�� ٰ�+8'���j��G�B�#����b���X�ze�d����!�k����]ɛ���q�pw{d��U٤5G:���}h����RcF�vm/�	�V��D'9wk��2���;%�Tz���s�"X��{��"�$�V܆��x!�c���F-�l�%庖ɵG�Q�d��%�U �_������ˉ��CQS�wॕ��7[�Y�4 s� ���uFcZ>��{��Hn���L���`�8�xH#0d��,d���f�Ru(�XwWJ1-1rF}h�\�V�N�Y�ȡ`B��vɎ���g.��eN4d�Eq��c��x�����B�̔��S�+����e]�n	N�e@���w���.���_C��i;{4�B�kl�7�m�.`,�*�A#�4�9��#l��rE�s�/��a<�vo���L���I��[t�ƌ&�O�WN�q'����ޥ���$;h��Z,djFI�%艸2ݫ�Y}�:,��jt��
�m��-���u�^5�x䘜B�?K��֕��)g�����6M��	`� ��r-6�Lf�6R*�uv�$�k�]�����e�	E2.>+��`��q�C"�Ѷu$'y4jL���(��Ϛe��dg4��g����4�v��7�q��ʕ:1ftu�m�o�����C]�0u���q���:��
ib��r�,�g����[�0�%��V{/�fg{!�O�]ʂz��Ni_\촸B���8�<5���f�Ԋ�ɿ}U��w\̤pt0����=;�$y6��|?�4�w��1ޓ7~P����_��@ƒ�����r>�^�oa����Dk�1V3 ��]����u�恣�����0�����8׏b��xl;=�X�!�<�k�N�d3Y�5]�1j9��`h��;^��s��{��?L���~؆�T��z�>�)�} �r�ϒ]y��/����p�I�<��l	�k�aH��lP�p6�q���$~��V a��sh���s�.�2A���BnJ�b�a��*���E�Nv��ο������s���V�8|m��Ҍ���r��Ȁ�ڱ���*�ҋ9��M����n�Vg}�Ǧ��sQ^Hdm�<8P�O~�_fY�b~j����N!A��E�G/�>�4�L%��2��Y
��Qz*Ki� C59(��R_�m��������s��"�<��%Zu���S��b�t-���ņ+^�����9NM�w6V��L�����]��:v1��޶����8�-��{�l#��g~@�4�gl+�N�ώ�y�{�UL�Ǩ>����Q�j���	~��q<��r������Q�*�2P̑%�<h%�54��:9���[�����F1��Tݎ"J�n��߹���{P��u�r���k��_ 邖����{V�%�M(��������l�4[�x�4Jm#�Ò�� �b�6kh��eV]���p�L��lY�ãs��|��b=���>�gҖ����ܝ%��a��F�q�K�i~�	�?���L2�a�Q �d�{�r���$����݈sI�����
k,��߃��>�ǳ��:Ue��x	�N���Vp��1�S�i�F�W�!ȅ�ɡ0�p�mۖ@DY�uh����}�e��n]��G6�ȎkKmOS����(��9�6@�M�]4I���(Q��4k��*��S�Y\����*o}Lh��+��I�j�L*��?�T���]M�� \#�{�������p��/3V;�	,!����#�;r�k���Y��N��$Yo[��5w�s��#����V�w��?��D?��<���f��[�q�lm���:#p�>��)��I��)v�X�F�{���nR�?�i~7~�)�k����@xK沍����Jq{5q�����\�}t�G���!]:�@W��ܤ[s(�+�$�PФD�� ������U˻Ӧ��y�1{��E��̓5-4}�`��N�
�����oY+f��Q�*̉�9��S�c ��N� ZO��`��������0?\�;0�Ek+۷���.-�u�rkw���-��f�`��A�&�{���U���|#u�Jns�0�m#t�u�'�3�;�f�h��m��O�8����tA0�R��+2��A����Z�@m��LC1��$�����?oB���� �
9IB��ꠜxv�(�v$3R=�OԧBh��Rԍ��4��ib���$���%Y\,�\�;l��K�:�~!N����v���-�r�ՙ��Eo�,��I�,@�&a)|5O�����>���̀�/�V��<]w�#G�N:����bX��9f!S��T:�s }�ܘSf���l`�K
�̖�k �$eG�H�Mx	c����ld�ё,���*�#I��)�C�6HO�,Y����"�٪{�c=��s���\�A�ƃ�f�vx-�~�و��$���o3V���|l6#<Zٰ�O#������x��������0Ƞе�׭/�]�S�d��$���k�P��̬�ޅ��Z�=~96P��݇hΊ�-�~X���+���nei�z��$�a�!��~��B���b�ơ<4��@�5�РdL*iJ
L5�_Q�lW?}YR!!(Ն�,v-i�Ow��O��༙x@~q�ܖP��	��BP�I�g�U"� �0��ymȿ���
Rc#�O�on �d����ᛎ�c�Jc��i�/�HF='U�����8��1�A���P�wC}umL�1?#�h�[IX	��7<]�:�\��P��^���f�(�×@�1<��$ Ugn|�YF��>��z�DGXSR��IĥU��IA��!
��h1��_@����#�ְ��I�~��Z��iQzy}���$
���WuT[�&�3+�g1��2x�E�-�q��rvH?Ǒ���Bo��9A��S�'��'�eo,?|������Ú���`�q�1�}��EěG�m2~w�z��`�jݻJ����O4�׿Ww)4 *S8d�+{;�g����i�����%��vy�J��Y'R5���*Bq��V��\ƒ1�!n���t��>a�g)�k�@X|4(⨃S�W��V�?}�.b��!/�u�R��@;[X�Q�j��a��V���C�v"�c�2}m^���tK�_�y����jNeE�iI�%a/f���Y�+=}��6Re��O5�K�
�p�L�+L<5Y�����!gF��ȴ�	m~�� �����L�pM�lu���N��m��BpA��)�"џh�?D�0!�]q�U1��U�:��ኡ����av��>�N�|s�+(D_�s�AƑE�F��?�=������_:ಈbX��p�כt��5o��0!9ڨ���FT\�\�.�i�J�r����H������WsT�pt�N�^M=E˙V<}�a��;a��T ���iO���t�p����+��J?�� �D�����c]C�t�!��hf��@u��v=/���T���}�lo�<�A����D�*��Ԧ-���<pw����;>(S�
ia�o���seU��VA�c�,�Yq�!��=D+5�h�dͅ���8����:��3h7et8~H�TT�\�֘��%]Cg����d]��DuGA��
#-��[�跆@x�D!�CF�MU�U��:��_��G�G�2m�o-��?h�`��n�{���%+� -���$��1ٔ���iV��J�)	��$xl��\X���,�d�w��&%�!^�<��>��Ã(7�h$&n��6�TM�{ݲ��=��3������8n۾`u�<��N�W�EN��-�NU��D�r���P��kOM��}�Z,z�T���L?�Z9Q�@́������?�����<��4~ �3�Ъ-rt-R�Q�TxJ_f�Ua�%FJ�Q�%Za�n[���`U����&@^�]c��\=!��;�������+&��eiS:E�$�+ix��e~c�A�r &��N��7Ψ�S����g<2.���%�CF3�K<zܻr�ჲ�7��V�a\�ʾ���3��w���EK��c�#�D*tͤ4�]�~]���|ܘw`�8��lT�}�3^�&��s֋��O�)�����a�����
�Ϟ�:Z޸bJ�&�����Z[�<4�E����7�nNN���(����!�DЬr912��#�	C<+9�
�J�0�9������%K ��M��q��$8�(��6D5��_��)�;� �,�C���d�aҲ�|-��pv���b�_܆���wr�h>WK�tgX��Sh��"��w�#��,�t�w_h*�R���'XFNg?�b�L)	�r��o��,K�Nuo/);-��u����)�s}ρ����v�$U�Bq���*�<�'Q/��XY���$�΢�t$�Άcܩn���S1��������RG��� ��&�{[�}bB�L\���o����<��㊣iD�4�{�i�vP�"�Wf�}��{�<^LK���h�ڥ3���� {���&��$��?�=��kQP����$�!a���3��q�3i3�[tz�%���
���5͵�,$��0n��̰7�XL��f�zS��!b�B¹V�x�T�P�wvԘ�/� �>z�'��V�2��Q�$�,�װ��� D�o�̶�RHW؇�z���� -eg��J$�#|�cm>c[��J�w�F�������� �����:8� �*�#j�-��Ȟ��B(��?����� >%  �O����PU���|��g:�Q7��h�w�����8���Wtx���l��i�$�^�aQ��A�,�(�O]0"��s�0�6ϭ*�7��c�!AA{
�����I��&_6�1���Ϩ��

���v6��XjV#��r������9� �����A�@�1��j{�1�B�mE��2�WT�o��{�������,ׁ�N��$���C�����3��Cz�C�X �iw���n�#-�(�c]~q�	��'��A�G~1��mʩ�3���I"YH��"�l���@���O��oJi$��^4�`�:�4�"�$n��=����HH\]�)�ن�p�#Y3��E�(�;�A�tB/�s���'�6�Y+(P�Lu :
��c�`y�u(�`%�B�u�Ѱ[E��]%�ɜvf��Ⱛ��
Է��~_�Ev�'�`�ȵ��;)h~e�����j�f�������Zr�̈m�����X	eQE�_;CÍ�r�|~V�A;�r$Y�����H�;�.��0�L\n[xlPD�K��Ǿ�y8>���'������hD���^��b�;=pR��4��˒��Z��J����ʊ6��$��E�rAFWZB���~�i��q��
����|��?��|�&�N�E���Ͻ<�JzL޽r�p���҂|7�����X�X���dC�ȫ{XM����J@�����:Y�`����={�>p�!!#U��)�h�;�������u���y�^�,��{§�����=>8.�?\|��45Q��2`p0�φ5��v�.���~Yu�R�(��� 0N�*��x�8�??�[��l���a���t�g��(j�
z~r:ܱݛ3�6���u�_��[QK��l�*&"(�0s�����1�zWn|�f3��nl�H^v;4݃�z�a^�3s��:3��$�CIa߶|^�v�ޣ����wD�C��.(}I@�#��D��a�F��SĨp�����w� �N��\����/�&�Z5��/ȢGԮe���`.f����W����]�?ǽ�h�ԭ��?V�`�W_����]��2S��h9W�������9�B�*#���,Q?\޷m~5��JA�����ٿ�d�=n�˪�x#	�����+s<�!�oާ�z6�?��iڻ��l!�Jm�؇�����N�=���0Gϒ���%�;��֫oe^ԀIeYkl��0���gwGs8��)���a3tT�@θj�Ag~|��#��(lP�l���\��VOSVm,��rĶUѳ)�N!�U�z�xY�,�w�]~��>M[]E:5ԧt���\�F���WMKw䖰� ÑJL�øa(�N���GMb�*h��}�0oQ��|���"{{B�7!t�⻭I��׸��҅��w��7l_��Ҁ����1�׊fQ/���o5`PYp�!Ҝ�?�eۚM�:,W�X�{,
���O����L��-i����a:�.ۊV��ѱOk�<t)7�����Zg���TH�J��g�����O�jc����'��&f����2x"��"�����ӟ/�f�C��]�ZqT�P��_uU?��դ�*�3����wvO��`̅sw�����n�Ĵ��i:��}�Izw���5ժ�f-&*۷ �#+��Z�f�>e�D�L!7|x�h�����.���D��,��l�mp� �1V�JvU)yL��*�x�I�ve��D��ew�r����X�kL!c��v�C�5y�#@�i9��ƂC����{���U��Q ����;����|9���/5J����H�~���Е�7K�Z)"�CFM��־wV��W<��E�9��J+�^%���bS��O�H�6�"!��yW���cʯ`��U�y�Q+������D��(C��9%�����js�֒�^v���C��*yq�=��,�;j�k�Vd���#�2�]&���>o4"[�'�n��?B�o͑��wQvq0$�f�Q�Gj^w��Z)����j��5�*z=���H�֣aٴ[N�,Ӝ���|+�bG�GB��;Դ�5^ʥ������zW{����Z+)�8����s��d��ֵ����!gfe����?�ԕ�� ��h��;
����sV�Ӭ[25�*v̰���3�ʳU�����#6�Rk����n�V��f���w�dc#�Tw���|v������G.2�Y���;ya�F��Bt3LI�Zd��f!#LQi���uw�g��1���&ӎ���ň�Y���11S=�u��k� �nA;��0�?6�2�v�:��^	�{���|��!�|K-c��w[@�8kLK�)Gv��%$@��+Vln��s�Z�u��IW��^����я?�_�X���t��/>��TQZA�S�������Lc�NV��$�\�lR v.1J�?Vk�=�H�{���t���/�o=O�l`����}kt��:�ߋ��\��\"ѥ[��1}��E+Ͱ�j�-��wB[�]�0���D^�MS�O*>^��������+9Aw�eC��>ar:m��D>��WGr�7�f�*�+.�Ť�6��P���k�8�W�ZV8�[�#8����2����_}a�"�z8�f+֋>��r��,�Ģ&+��#���3ܫ	���l��:r_u�N�K�b���S(�!@蝰�3�����؄���WV
H��3e�f��w>�ސc[�Zܢ���{� ���>�77��E,�9�VF̚����Π��܃9'�D��pT��*ů.)�0yǳ�7#�S��X8�d����wD�U��a���	��[5��R�a	1j�Ef���ۚ�� ��`y�Nq�D ��7��̼v��/M���N�ŗ'���`e��'eI�MT�e��T�@�lpj��}p���+OwB����:��F��Bi�r�][�wm��V㿕���&o�d➛�'ꙍ� 3ˢ�i��� ��ͩ�5����]��[��S�қ���]���ο\N�U5r�����N�[���HO�/@��G$����v����^B�MM�8�ۅ���)�I�rC{�5Տ8p���qQr�Z1�Q�1ؘ�ׁ.^s࿰�L�,4���rPF���ɹ�MPҁ�3��F��`�"�^N:$7��3���{�Yϫ���w�f��5U���}p�#D_O	:_܅���E�2sBN鱊"�yd'���!�)or��;5�FC"����\S�vj�����{���v�A�T197��
������s(�9���pO|T���6��2�%O��,�~�A�qI�p�ׅ�y�ωq:�����m�q`�kQΩ�p��Ә�s�H�1�|ڇ8��{�ZF����D؍��HpȲ-�@1
+6��� F�x�Z���_~R����N�a�Q{���l���+:O,V�YC&�����׻�[�(~��އlH�F��G>{�_������Y)b	�(����Z8^b�u�\�+ò4wK�g� �A���_K���+�x����!��f��d�.*f෫o�pkm��.�Hrt�NÖ	.P��uu�>2��D���r\ArH��<Zʹ|��(��P�>��X�E
��vE��[�B�e���R�
���5��8�'{ܣ�9��]�Y�5��$#q��%J_�6Pr󜊋�bX刘��}�Qf����)�ϐ !�H_f�#$��Bqre㪁㒗1F��"��[�Q�� 
k��s�t�C��^�����M�I�e�GH~PI�?���F�#}�m�9�r��4E�PV~��seA�I�MZď�u��U5�R��R1/+���O����P��P�MDi�}���啻Y}�|�K�۬����D�xOT�A��V�/b��xJ�B�0,�#�#Ƹ�W��
��V{�aVSy�õ-����7�8��ύ(��˭y�5%�������G"��_���`;s!pSz�7L��G�)�_4��v�`��U�ⱂ�5�m��I�<��$I��b���_vWE����E?C*�R�{��0���Ӂ
�,�c׵�#7/ڇ���h$a^�چ�lpJ3��/���`SaԤ���O��Z�Q
�t���͞���������Oh��x���/b]���A��"�ے�Ɂh��iw�dBH^f��a�C6C$��fmx+xx��%:^3�^8�,���y���(K"-�Co J�/�B�^�*(�K��h)<}w��g�<lq+�&�����*G�ħ���Q��3�	������Z�t΋5��ׇ�!��T�-,DF	�d��ܼ��*�u�@��d��}^���U�Z��'.$Ѕ�h��r�����Ϝ�װ8Ō�5>��]Gk��y0Wm`o9�g�vP̚�L�V�5ێ1[������V'�Zː�{[`Y�)��RSĞ��p_�opf�R|�74Y���w�Y˯�䇣w�=H	�>'�?�:�� 9b��Z�o���a+mS*���v�J����?NV���]H���f�:O9y�[󰲆M|؏k?���\Ja����{�L����܉�ηX����F��1Ɵ3 I���@��y���a�~����K�d�ˇ����w�7���\(�"�I�_@��G��+��D�\�ULe�,K�a�������A�!��\A��*�C��s��WX��`Σn��}��1���'Z�:��6~d�{�$g��)�pB��'݋�^��,�--jh���
�A4�b�a^!���u ...A�d��_���:X��Ԥ���� �;�$���w�3s
f""�t�`K���o2�w��G*	J�Mhs Ik�L �U��y�,���n�M3�I㰨�M!PZ�B��x������^UQ+&P�}\#٭?�'��B���w���_la�m$��E,��M��6DoMbp��ɋ����fV��z��3N�`.̫B�A�`�BVƖ��%V'^�=���>�����Fp[�)f�q�y�$�Ӄ��~�$��?�n��MH{��K�~"�殽m�؆,�O�s��Ȧ�!XK�O�p������	�@�
�V��*	���0�C{��`6���y���)��4J���Φ�����%�k|�|P�=��#d�_ecG"�ƣ�
�1Qi[�!��A�,�/ܿ�{߱�G�00�����6�t�~��M%"��+�x��a�����g�o�u��}Nn2�4�}��ԓ�7�1w_����N�G}/�k���������?���6�������^zny�t�*�>�W�9I5B��#�,��o��9bs.#�����V���;$dפ�^����	8q^vϒ'&��	v��^<=�yn��#;:ۗ���B�W�R�_F�*����C��Lp�sX`ڪMS�`D���$r�:�K����0� �'B�Z&�UpJ�C�U> �Aq��i8��=Y�I���^'�Ōx,hi����N�a�V�����CR� N���$`܍���a���#=��$��x��ހ+�xU%0�,[U`]��Fjô����vY�e��'�l����y|L
n|OI\�dK-�ZtM,�ʂ�w�~}$�z�-��Lw�����@�lҌ��}�7���=��g(����FZ�a1���7��sUa�cT� dﹳV�C��@�|QJ��X�s�3���%��?�W����𿂫���oh=��4uC/��������DB\��d��ų|���	zם��<�X}X%�ۢVj"U:�mg�L�hA��S�;2l«,ѷb�߳���N$�U���HSU�<uWk�4Y�p�,�\:�B��s��e��:�+�&�!��2]1Gf#���*,K���Q8]3#��r�Q,�E�Z2����Ǔw0�%�}���N�Pt��f��޽ȕ\�A�e�%� ���;$rZ� �N���e�������n"wϡ�ѡ�ƬQ��j"��՟��F�eс=G|B���R��'���}��m���|�G�
���y�;`u���W ;��)�xhK���C��-�zM��4��N�Ē�+i�`�N��:Z�J�tOoa`�=$0���6<z�$��є2��ke�#�GW��$$n/vX�N��O#����\�A B��4CI�: �'�9D�k˿7���R:��C��>��Q�=n��{]�l�,9�~���1��Ut�ao�����%筽�D:�'�z>n��b�-s)�c҄x�-lt�t�ּ�j�	nTZ��O�| �u{���f�;���]x3�ei�tl����{�e���g�fc�b,��|e�(�R�Iz�>�䤂���h̢�	��=3ǰ�+�����;�V����0��T�.F�����`��.���/���r�IV�![-�x8a�i0�m���r����,���v��k�:U �G���%���c���H�3Q_���R�tf�w��@sP���"��Vʞ+īJu��.�3��&4�{���]��)!�cC6Pq��N߿��8I�y��.� ���O�Iq�r��I�J$���e�I���V�-��7h ��J2ķ�硴�B�К5v3����?�ο�WCL��p�}��|S�:0�": �H���(p���R��$�a����y�I�A]!� �z��(,|� �������p��?$�Í Ռt܊�����"J���(A���6�d�V���sڏ��1��!����;@iR_�ד�\�n� �Od~�;��g$���$�B%����k+F�g�$�<��bi����L��ܯU���t{��s���NOA}_���R��=���)~[ �9��$r�{�=�ٖM���ԟ~�vB7�M�#�r���9ͦ������#C��}�m�j�]���d�SF�_j�v�I��&%x��(�kxE��s��������ͺƼȝBv�C9�kL����"��%�"��*��6 ���%S+C.�KA��p�ۤ�&���+����"�u�����oɛT��������-�mI?y�(�5�"�C)�'�.L��N�~
yB?�cl�1>�k5<�zb����1�sOғF���y��ⓔ�G��o*��d`2�y���K7��=c�⬇p�O1��mv��Q:��Z�<\o�E �Ԟ*EX�I0<~�q��B��dJ>,�v���G�6|*��o
��;��J$��$�BK�D��>K��a*E�T���z�ޟLg��f�k�&J��'G�'&�9��Q�WGʟ�~\�A;1ӣ���B���s�D�[`�Oy��EP'�+G/�S�ëhi5-d�QL�7��u�E.F&:וŋ�ۅ�k�ڋX����X���I�
ⲃ���v�p�)y��yt�m�A�P�db&p<i��)�ypZe��$�������y�RV�Ɋ�XAN�*<Ck��7Y+��Q��d���g%ޥl:��0�z��M[�83�t���;&�Y�v.����te|�د�����5���+�W�
B�pv����j���M�N�4L����2�bߓ�� �����%��^S3wG|�`-\u��he�m=N"� ���Dq.&�ٴ��l��J��Q�#��2��	%�ag���b	�V���ݱ&W��\aEnMO� %�Z6A�j�=� "X��-P�P�:5�.��������Q� �E0a����BP�,����׺��u}�G43�ݜ�03�=�^�9����'�3�(XC(��|��8�W�?z��Ħ�#D�P���	�)�$���S��hhq^���'�[4�2�O�,j�(Z��ٴ3�z��О�#f��+��	�&F:V@�����}adY^�}l*^C��[���/����rC��H���.����M]
�XT��Taw��ab��"�#��02��&�q	��]\Ѭ@�)~���wl��A���B���:��caC�5V�$)U�!*J~�B6ix7�vpwY�8�l&�\ٛ`j���kI�9�@vE�ܟ�X�><�E��jh4\��/5�I�CU�$*�KE������	�;7�oN]�4��/����n��h.��ͺ���Z[�o(�G�\R���Aa&�k͆��RKO��.ǟRsA�����i�W8h>��\��t����Ujy�ʒ+���+��ӊ�:$�"R�>����D�o��׃<}s|N��]L����¬�u9j���$� ׾�h�93p���!�l�JI�'7������S�^��"�fD`FG)��_p���w��
��v�7�Pn6���
H����(�=|,�a��'����
�\���i7���b"�����@,���-��X�{}�1fAtz�,Y�����<�ۨ��>�|�6��e*���`̤�뷜�H}c�tv�Rps��K�v4�Z:N�m���O�*�����3�}�6Gbw<r-�[Cy�u"�(?���L(`�jc |��H����o6��y}$ܿ�s�\b,�,�f��md!`;���zA�I��4c3���⚷���J�N�?�G�������	����@�v��<<g�yS�Gnx<��I,"�)"�M�����E q�9���*U�a�*�;9]LȂi8�����K���.���}�+H.�q�1z/�+�K.�13�|���O1~,R���W`@�5���K?V���@�Քn�r�y�|-���J�ya�;=5�C�_�@�Ak0e*���2,a���N���N�������O������jD��&�X��b�ƻ�����%������g�$2�Q��ʹ��n1$}�i53���,iȃ���&0�M���އ���t�F�t��U����U���q���7}���5�ةUhE^qq��aU�+�aa7W�c�G��§���ی1��Ky��P��dB�������t1������� E�q'��P�_6<`^������^0n���C
N��k�0�H�Py�ϑ��ط<������9���yZ��+�x�N�}?�&�:���������9,�im�*�,)�S ��g�o�X�{#�ë~��9W����arDФ�bb��i�k���i뽵T����4D��3�MD큦^}�h���C��0��%)��u��hw�W9Q�L[a7�;����`	۴�+���j�^<��$^�c�_}8��GZ�;U ?���j���H�� �WyYز�R��Y���U5����~&���q�W{�>56�����TԊ�&�P�59�w@Q��,]_���^}d�)�U�:�)�w^�ܻ`���K�����ӱ+R��T쓉oƑ��u�C���v���'碛_�M��	⟩C��U�P�r����t�<���˅��(I�R|Q��g��"�P�Մh�aDc	��D�]p	۲Zm�� g�K/�.�j�Ӗ k��m %�m�H㚤��C3�O���� �T�߁�n]Ɋ�_��-Tf�I�2��tg��P�=K-RmyA�[#]d^��j�n~3���R>U ���<N�v]no%�j-�w�[��:D�\,�����_�XE�(8v/A��l�\X���(WCD�[J+�cL͙�%�����8rB�L �敳���Z�8QSr7	� �im[p�����7���6�-<�@e�&���Դ�����>6ڔ��F�/�ל4��<��ۏ=�n��[��IWbKMt�QE��r�i��,t:�vs��/�/r�"_�QV0{���9����{7��O�G�_?04��E�Δf�M�Ǥ9�bk�_���w�_e� bG�u�p:����D(W�h�����)zW�I�3�lk�� ��)R/u��;؃W[��
^>����ה��{_��cR�_�N��u��f����6̳ {$�g
TŇ�|AЭS�k=��zU=��rC���	fJ�笁R{�x��"s7�����n=A�Ѿ�ϖ�@�|,�g[l��#��*0g��D��p;_h��u0�����c��`�����6�E}Y|�
�ӻ��18�vv�(�ŀy������-Ј�[+P���6ɲV1�+����_�M�1/&ƏN���Y���>��ꕆ���C�}s���[��q��n?Y��[B���	=�H���6�-�5��P>�����z��&���J� �%2ͥ��kN2���a�*G�	�{~�
�ϩ���J�K��g�8�?hC��Ž��/��/��3�ޮx���[�V�Oeķ%{��Y�-�V�S�iS�~ ߩw'}�2#��������:K���7br�Y�n����́�Ǘ'$|֑��=5�V�-�#[��(|0��v�3K_s����Hx��H���b�,
E�f�����"y�S��ƾ��X�"�u��������Ȟ��<a��@��u��e���$S���ڋc��P������`rn~)
�y�lgn+�nke�V���sӚ'Y�縺<�%���;P�9 �����:d������f���̍ZU w�j�"Rk��z"3�2�q����f�It����>ne�y3U�=^w���'g��1��7���JE�6x]�q��ujN�����)�$��)��VT8NÐn��+����U9����Bb̎�,���4�t��{���_Q[0�}U�`[�6P+�Ip�=�0��j��V��%�9�����&�!��*@��^ܭ�]o�+�v������qc#� �{��̿o �Þ['��S�@�����yxm��Q>�w�\ºU�{ �A��z�1��:���~�������
����B�w�� �����K���Q�l�K��dD�ڡ8.=mdhy0�9L�(3�捈M��D����Y<+hdl,`X��f��v8�`�w�g�9��Hpdۍ�S�*BT���6>G�a�5Ĺ�t\�џ��!:��4�>��]��F�GY��aI����J�H�����&��aVL�r����J�4��MI�����P�a^VQ�)����[�&]h�F���Q��z��'�&�jfI�U&Z�@�UIV?�$���!�`�ZN����0M��l�}]�I�|���,vW�Ά���4k��}�f�����������Fv �=n{鲾jhd���n@6���i.O�0t=)K˼,�*<'ҿ,/9{\]�w���	HE���L�6��v���ӋɄ<�(�~(r�E�:Ve��s��A܌Q5i�Q;��_���Qڗ�{7C��W��"��c�4�uK-;`�m�љ\nlWCq\�#�.?hI�6��W�&ǣ>a�=��N�O}��3ݛ�U��֗,��T(ߢ׸��GQ���_O8ޟ�ѳ��؅?�ZD�M`T�D������ݪ ^�J�+���"����iG�,�F��i� ��j��� 1�>�����S���n��WO��EY��,�Н�C���e|
a�>It����+��g�.I�l��&��?�W�=Ta��H�; ��ھ�#�9���z�aL�+�&�5��o��Z������=���Cc���A|�q��Ԇ��7q��		c>���XP=�����Mk�i*�m�����#!� 8*-.0�q��JD�����,�pͻJ��d�|�iU�h �Y�����&�7��SR��|2�m(.ڭ�3C0�/�����;3���1C_b�pԠq���K(P-=%�:���"�T�h5,�֦(L���$aN�J�u��!�#?��;C����ڥ�ˊ�g��|�c�u��dW�NT�2G����G��Uރ��`Zb�(������o���%�&�����{eV�u��~l��W (�}�i�X[2���9��o1��|��'���Tm\mD��ݵ E$F������J�@�s���Z������8JN�6�S$r��צ��h�RL�ۿ7H�Ʉ%�
��y�ٽ����
N�6V��Ċ����^��;"���
L!Ъ9��gW3�E��J��I���i֕�+�ڴj�8�2'��^����F�0�cS�@�xk�6�`@x#*u�!�G���l0Kez�%��V���i%J�<o�5c�AM�c����\moI*�����������S
E�(h̤M��o��Ѕʪ�n���A�?|9�3/���bsP+��ΓC��X�=�厢�_������&:i����p���aF|2͇ۥqq�j5�,^��������ݪQ��딊3_�t����^,*XD%7W�cA5�۳5���<�R׷ۦ��Y�`C�'uN�$��u��&rx݁&j�o�m���M0�Mw��f�ur:��>(l�`6C]�RJ��0<W^�t�k�
��~��ɫ#u� �p�S���`����nBb�����a����(;�1��Z���B/�N�s1pSb�\%Uv��
3״�\�yV71	aQ�?�<�L���g� #v��!��m�Ұ�6���l���ԕ�����Ƨ}�7�3�6���~�*��$
q�C�+�)9?�W���q�o�!�~/X���c���>��+��.q�h�H1i*��[V�:�u�9WeR5{Xh�����*ٻƂA��
����˨����U�s%89Eq������s��fd�����Zf�1��N΁a��Y���Q��㕎���E<��ǭ�7PM�'S�ɘ# �|�ZM��=6�F��G�%�y{D^gD�|���y�ݏ��s�^���o�fgXXL72]��>G�u �5{�I9W*�cx��[:>S��$+��]�wBb�,�QB��/�?524 �Q��g\ѺF�����1KP�&	d�T���܍�J�d�wR=�NZ'��N@c�8
ꤛ�v,a0I7Z��vH��l����B�G�gv��S2~$����P�6S��è������ǫ�蝦��l�=ꁖɤ��{�UP�]?y���pr���`�83�?�l�����wgg̀Y�X�t�Z���0n%��/��<�v6���K�2����!|`�a ��ғ=nh\�T*��s^�{���e@ΖΟ���ǧ�{���2���g��c�4K����'�6����`�X�Jk<"4��3�����Ћ���modQ+-�PX	��]S����}@��TC�xɧ�_���Lۮ�L?�
�%<,�ƅ�Z`",�xf�\@.B�HR��zx���.�9vXz&��u�W�<����MH&>�O$�g�y�L��,+�G}�*�d.L���	�ܔ�'Ng�c\/�V���O�J��'�+f�&�
�[9�x�Yo%�*k� ��X>��1��;���q����6IH��������U�'�_��'��1�` zl��a>�0�ts�p�.�TcX��Þ�?��F�1�)���:z�F�D�m�Eڧ�0%g��rќ`ccw$�̄������x�.M72���]��^b+`]��O+v&] G�a���
�W��LN�[�u���~���b�������:�0�)��;�_l�|�
��5a�6
�f�mvp{��v�����z� ��=p��O ��C���2��:W>�g#��l�����M옛{+i�q!�������u�+T?�!Sa}�q���P׫�(T�/ �Qe��~�8�҇���'.)�;@E�f�A>��NY�?�Mgc*v\�SԽv�sC��*.c7z�𣎘��{�Ο3t�Λ�ə��#~n��j������R)��d�dSn����WL���ڋ1p�Xb-���`��U�*T�腑���'v��<���n	�݀A��g�`6��a%�m����� ([�ke߉��g�1�.�<B���'l�mp��>��K���rb���*�f��೻�=UZ{�ᖄ����q`я6Kolki�d3�dj
��AT�i�c7B���ӥ�)0cSd��z+����Zv���K�i9$i�d?o��%У/�@J�Ƃ���m�"��JR��ǡ6��A�]��)Ւ�'�|'�g;o�*E��0E| ��9���~K{�u �>��F��GD�Pn79���]�HAP�]8fnk�!��vI,������
�o [,NBl+_��C��g.��ݗ�'N!?�e0
t�Z�#Zx�
��k�%�w����>�`\(x�RD�qR���㇐i�J��;[)y�z+�s��7G��y95��*��`%����>!�Pb5�w��V=/��<�	�+�������j��İ���������};6hQ��J.�UFƃ5$b�;��Jߊ���>R<#�r�a��^�y��v��f4�ib�-�(C4C��n���D��|�tM�V��f��2���ì�D��F1�\�`��U�lE�EV�,e�c�ɘ�W�q���~d	���=�@���k#��h)ۆ�{��>��+/7�jXF�����1X��-S�t@��������={Oo]/�Ga�az��x�]���s���ag|V򉕛�}+�!��SZe ������A3�k4C���7�>*3w�L�ĥ�g�0��ؓ��t�ɾ'|��fT��^�v\���/#��9]H���f&D^5�F>C_9|��9�b��V�&1�oj�b0R�d�qV b�hA뿣>50�x�s|����6%��BªeY`�7ǰ���>%�_6z��4�j�h:���/�9w���mz|N�˗��<&�l�h��-Dh�/߽E���_�V젥"l�KD���;3�-0�n���!'�|}3g�����_(��縴�V:�겯�f����3Pghn$��s��&S
��7��ld�K݆����9KHt%G�k�AơO>#eY��@s'k{��M�TۢC�v���� ��,7��/��0�f�٪~�q��>��+nVhM@����4ԒVh��`��g˼�LĽ�$f�� 3��=椲_$(���}|�/^a���cտ-�鈧N����BV�|�/�&�!y_�
�
��(˹F,�Ȟ��évc��;��V�q��S���T�WUv���wPO��^�[�/j_����=�
�8;�@b%�I�wցӶ;������~�B�/#�O�F q�R���XIF59n��)������v�x�D5u���E�k3j�=�n���H��*�4QdtU��^����2G�(/���Ie5^��{�᷆� K�u&A�V2i(�s�=���,K�T���oos�S�����P�I�;���~rd�o`��I�X���`�q�u1��v����Ù	ɖ�;n��$�A���;��;�;YF2�U�t<]��E�p�5{QZ�!Z�+�Q�_A���.״Fp̓Q:w�\�̺�~��;4_n�-E��O���V_��@	5��[�33�C��,�k�p����{&s����!�N�o�r2���	��~0]0�Lg��K�'�8����g��E�"i��kp�����A\Wó@Фu��*�2�������%D"��؇�����#/�^	��"�A�@���k�F_�<@�||��l΀��?�z�*�0��Њ��f��ٻ'H��7����x�l�]�	(z����Ó�c��^ߞXػ/��u�-���e>�; M\	��$2{�m`����A�O8Z��x-��U��2�����i�a�v\á�&��E����rzо���U*,If����k����^v1{C}K1a�1�P3~x�_���ݧ�a0k�:� �\N?�Nyrdn�&@"�7l�,�P�U.v��Z��`��6$��	�;�A��+��xFf0?�@\7���i�ok���p�aa��|�E�]R���D`�'y'�\�Rz�^�Ǚ8S�fd���_��U�!�h&����I�fѐd�b�N�W<�e��;�M�pH��I��U��g���� z�c�u{~mMIA����3�Ąh��Zb~�Hy+~�\��`A�n�^�S��t�e�	�7G�;�q���m���孬r��԰J�rv�.�͜����G|��]ۈ�����$����U�fm�c,�q5�I�}ȇ�=< %��F��K�w���p��?#ND1�8TSC4��8�����ĪI.8¿j�Q�HVl�)qM8R��I�w6]G�_�'�\r�u�Cʿ��I��������jذa�g`���U(?���"e�@�� �|^$N��AmP#f�t�m�� Q��g�Ɍ��z�K�u(��{�Z,�:	�8x��B. v�}PdlF�մb���J�bk;1B�3 �+h��ͭ(�v�c>M#Kf�맽�;��^\��#�{��jRo-�nF=
�D��o��2{��s�ǝ��bm7;߃����Ԛ�$�%�n���I��'�����WcU�u�t3o��U�{OȮY\B�_�������C�*��g����F˫�k�0��7����ҽ���g C��w�Ev8��6������l�u�7o��1��eU��P6�^��V�Ih�zG�'�x�b�z�Ӥ@�a�n�q�#������+�+T ���j x l���K~7��(zB:�{�9���KfNz��d��|�Vi��<��[�V�E���rS���������=�N�W�I��D���n��
��pX���������������N�ٮA�4��My>�/�y7:�"�VZH�6<��ojZ|��n	�(����ĥ�W�I����O��r�^�sm��p���'�A<��5>����]Q
*1:�`��	�����2<�0��Sp�D1V��?�R	�v.d��ts���Ls`�ey0�����=���Q�em뷪i�(_E���q�ų��#N�����M�a�h��e�9��t^�ﻹ	#3���&���K��!l"r��c��#! }�к�⥂R�� e�W5�,L '��/Űܔ�Z���,��%�Ko-����CH5�4�O��C��H�W�����������~]^^/dh� �FC�o��Ρh��j��~mH�6CV[B�Ҟj��Bռ���7�}��F��5Z/��g�6���e[�*�:ք�3�o<Gߟ{R�To-9�L�4��6"?c��t��p� x
.�cNO�a8�F�=��%���)���ԃ���L�o��U��G���Y#�U�x�|��uft�D�;AL
q��4մ]���,,xfo��<��r�:�!��}9ԯ�r�Ё��m+�PV*�jl$�������e�T���sK�s�ln�[ILxUP�ӽY
h�M�=;^��������j��&9����(:'�Kf��f�lM�$'��"��o9>�6�����U������)��;�j�e��V��;���s�2�H��Zcg����>�J����ֵ�biB1Y�W���{���-�h���$
z.l��c�!�-(v��5f�P���Y�0E�H��5,��%Vc�'��C��p�[�i��`�� ���i�=9)S��3�}}��w�x��k�L"v:�T,>�Xq�_��4`a)z��Q��x����j�^���K @��_���e�Ѳ�l��4K�gp�E��E���IP�"xN��P%��R/�A���>��E�w$��0s��VR�P��C�$�j�H~��a�eڤ�׵���t1��3 �$ԉW���h8o�^ǔ8����́v�X��.{��/r�oOE�L�=Pg{�L諄o�����ܺ�� �ha�j�T���!l,����`����o�K��{�Nc�E���C��_mu�������?B�y�i0
�9m�����Uy�K�|�Ė�5�ˀZ:��R�Ы�t{���b	O��#�����n0�z��yC���&�*4��l�Ʌ�����]{p�zl�"�H4�' ��ɢ��FZ�u�ƥ����+X�u��7���p�[�|/��X��4����{�d+��W����Z��r��.��eHD�P9f�2J5�P�DK�9�,md�_˪%���4��Hs������
�PN}��|�O��C�{�q�:�X��T��/����kv�\���t�2�1�r�=i��������JB �GM𡝰*v(��K��̩Ծ����C���7�F�Ro&����a�X�hW�NA�"�-�����S74��I��]>���y��L5���ۣ3�
�?w"F�c��S����"�L��y���r�,��1i����9ϸ��z��u�.��`5��	3�����=�U����L$��a��V�x9@���
�����e%zj�� ���:?hY�Yoo��Xw�Ʈ�(�i���S_�&Rp�)r�Aa�_&
1�����R�_�#�S�f2
i7O��XMeT� �0�>�@�@�e�J���<&1�J����G�0�ze�V3N\T����X��ݤ���e#xA�ٖR�'���e�����݋�&��D�� ��7Sa�m�g���N%e��S������k���d���1���#�9<�XSMZsU�����?�"Z]��mݫ71ʭ�R�|��J��c�iGk'�Ѯ��t�J�3������LQ�Rۖ)��y�VU)��c?T0"	�����TY=t���\@�ѱ?,\��ӠE�ܑɐVX�`�ȰS�I�ULJ*w:��i�6��m2B�m���j�w�J���2	�c�4�aq4?��Ċ��ȿu���)��63�OGT��//o����$/i-��b���^�buaT�sP��$��ً��E�*��\��<�2��mn{Up;>���:���:�;W��v��#�^;�B�՘�������������}�����M�'�!�0+/+��c37���Zj�h�<GHp5�m���u,[�}�Y>P׵?.�N��Z������;��������)ʆk��w�t���A�*��dc?�
Y�2���^ܸ7��,�k�{*�ԝ.�+��ŘH���n4��)a��$�4ꏷ�+U���'*<�����9�����M����ȿ��@���s'%\��8B+ �-	V�X��w�Y�p;dE%���ى�v�˥ͦ�.��R�f�T����m�x0���o�Dݯm���{ �.���t!��N:xp>�W�,�����#;�@vB�\sUĵ㴬�n٣���(��<�T����Zh�P�P��'[��!j����?�SO����P��&y�Q}�� �p߀�� %�~�9J�4��%�}�2J����̖nK�@ռbp��v�<�%+�w8�p�D�z��J��b(��-�a]��<���`/����t���*}ο�<*H'���԰j
�Ry�.�2y%��@���ױ~`h�C$H�z���Jv��_�j�dZ�tc%�����ɝ=�H�D�z�ﴡ��G��(?l�YW !��3R�y�Y�����d�ۧP��e]9I�rk�a!���p:Ag�a�&��W�� D�����6>�����8B����b2��:�XJ��StZ���fi�i"�e���Z�,��7�B�����O��4Q;�,���MSV�i���$2	�	��Prٰ��R��`��;�8�m��h8�S]3����"�8I����|t@�z�2B���еj�U����n�'����7�}�"c�M���{E�쎐��妫��VERd�m.�{���\D��4u���n���WVxF�,`�8�d�u
GX�c�6k?o�V�Z�:� �9������l���4�3��!_�[p��܏���R�B���x�.�r�+RN��@�Q�����csob@����|���0��vI�յ �8��i�K2�� 2w�=ڒ�.���L����V�~bع���Պݨ��asBC�U��i&7���L���V��Ж�W:A���}�Ԓm6c�m��׎�����:�<�d	�j��q�'�ҡ�#�DS�U�05��Z���^�;>�QQ&�#�[��'QR��CH��]��,:�"����*R.%r���e�q._	�~n�J��w�6�� �����m��w�9�>R��4����D	t�U�<5t��I�����ش��Ĳ���FZ�1�q��ZR��Ά���	�s��H���	uy7#�P'�ҁ;lHW�������|�2����f�ɡ���ݎׁ%�;X�$d�F�0i��$[E��O��I>�J�A��28F�8����q�(��6
[w�THn0����#-����jaj0FY#+IX�������<�����	4S�VAi.���A���>������v;=�cժ%k�ϷTmͪ����D��i:�u�� {�#��W��z&5�N{6����@��y3�ZE.^�1��!��L��!KK;aYˑ0��/�nu=�b5w���4�#S@:�)o��,1�j�)�JYWftR����0���;��!ksZ�E�woa�con'��UX>�vv&��ˑ1� ��?��g�3S3�П2��������/e1�Q$p��)BZ���`�M��@p�T\d@r"X�!�eF��;����2�}ߏ��qR������_T�Se�&�y��,�r��I�㠣��8	�3r{�At��{��+�J��qM�W>�eÛ�|UA�-LEk�X6rՍ-�m�>��wx+>gV���	[O��W�ZjS]|X��s�`�Y�J6)+m�����E]�q��~�w�j�;|4�;�I�1�L��Z�]������37�M;؛k�^�W��Jc[J�נ���El����&1D��ޠG��<��`����,������
�S����PZ��.E�D��gH��s�RS�U1�\.h�T���E��:7n[O�*G��(Mke}#4�Ï��fJ�Pm溺������3=�TV�
����n�gm�U��7-ţX�H�׭
��SAU��~#,b�N�hL�b�] �n��oo��g���a�[]oD���������Пϼ �4��<������|�ivOj?���:Y/�B�N�z�E0Q�E`�3g�؞M�:��G>.#E
1��f�¯�v:�}m �l|%$m� ���	'�h��s?��Z��@��G�g��>���V�YB��g;�N飇ĸ��y7mr�Ny  �C�V�X������#����l��GhQ٣�s�-�w��9�3M�s�<��6�(-'��#���]�|��Ɠ�d!�_і�D.�yvҏ���$0u���Q�e�ɠ�l��lH�o�ʦ��w :���M�qF��+�g>����zq�Hs���cr!2τ�ʭ=��Kַ�՚�tȥ��7P�y ܥi��j����� ����w�3BM1tC���X;�[S�ߢ}U���ʐ��m��qV��(���껒�����p�c�2[�6�0ʸɉף�u4ӂ&�.�4����;Z0����C�%��W�����zφܫy�hH�Zg�����ȯ� ���Iυ_����7t��iA�^��x\"�4_rr���dG��S�~ƧLB��fv0�5	���'�*X����hc+)�_Dʗ*�p��D.i�M��ef��W�c��l6�{�'�ݾv��Bݸ�x9-���>�$��-�W�һ�Ԃ�f�[̝� �E�q,�ê�"�=r���eT�)}��:Ay3�Q����k'��Xh�	�B1=�{跃�F<-�}1ᣟ���n��`��.;�W�%�du��;L1؍:-���_�L��{{�ko���t�8�Af�*K�D�14o����=Ү?��e�HX���������:��{�2�Y1s�Jyuɘ^jd5�G����ο�hn�ꝃ�;���t����ba���M�oCJ�e��F^k6�ƹ�if�u12�~�"�̈́?'�R��%�͛��/���*I"�H<�E]ifByB����]�����V����ɣ&�#�%+�&w$��V8?������+�0.��x���}Jk�$�b����Ɔ�.tqG�
�W�Of����]���\[y�of,�Ӊ�wM��I�P�ż�C�X~�M�U���G[��t=���@� 0�t}�_k�
ei�H�s��dv��q�ܢ%R<R�	������~�&�Q�:d�~^4��.}��6�����&7��;�j�`�����2�A�$#M��򚡏�F�WK��`�~̑?2�k��{Ƒ ��࢏h�G�`�M��"��[,24<!�|�刨����`f�7GyNy�l�)��/t˖����b��u�=
"�����|r�K
Z����-/[c�,C~����N4u9��P�@���o�w'Oլ��:U�rZ5�@�3�b�}0!�ל��C
�X*G/J�1�PQ��Q	q�h�,yC_�`XV��S�V���j��x��t�|%��k��=��8�Br�h}��p��[5�&�"G�Ԛ�'
�t��(ϩ��w��0s�f��`��7M_6� ��6筬���4��o�Bu6�������,~�����ݤ�(�5Y��J�t2�	:e?��+��z�T�{���q�%�������0L�lPKp}�����˜]�o��CI�&��;� [�5V��6�Mb�V�d�OɴQ���Ml�$E@���(��I���ۂ�LE!
�(�II��	�N��hr�S^����T
Uh_��֩j�qvc\��K�1���eG�GAB]��aavw���t��O���Qb4ŉGZJ��CH�ީ�RY�h�0#��&J�l�Y�y�8"Ұ`�c9���{��eT>��?Z���$C���'��իb-�T�@\���t�ø�ڃ�>�:��,5�Slo��K�@?jx�jW31��7�����Y��r�嫦�3c�n��Y��}v��>{�5,+��z @%�隬ih�8���f���oD�������h7n��
��w��=lw c����of��bn�����	��ǅ�KD�>�4P[�5�:-a:{i�zV��1on�Z�:A�J��`r�ŵ��I ����7�#�U����:F�0���W���X���N�E��������J�u�k�:0�k�.H-����𦁱��_(¹���)(�7�������|�cY�h�9c��/����1i~$�w�b�o�%xq��I��mZ,�8���Y�=�!���L�Qܖ��%-E�u	��,俺���21�4����&Bӵ2��`Rx��h��-</:bx-�X�T��}�6�{����+�Z1D�F�7�{��I�k�iGQ��.���k�#��j�T��L�$���I����ө&�PF����1� �v�����4"��Q&�`�!N(�
@ ��_��d�w�F�_*k��+Y"!G��!L�ZPf뗾��sϘ��3��a���M&�t�O;�5���fV���|G���>(���~oI ����9ɞ������B$|��m[�b�XP#���S(Q#}�.ǟ#�^�3�5bZݙ-?�O��k�ˆnz�^C�^�Ό�.W�p�᱗W F�G�o�b�_b���0�I��Qe<%K+�^�[�8a&�����t��10ʅ]�������溌�9�{�L|zi,�֛d���1j����	���(\T����c]���iz�HT�'e;0)���T!�'B�T>��L�i�
�t7���>JIл��چ�#{Jd9k嚖 =ZF�묛j+9�P��.�{�$P�C��EF��Nh�a�?=i)R���9!q��N,}��\8Xq:B=�Y��䷔��+�U�Hm�]>ͤ�b������6�8.�D��-S)16e�QG���b�r�����A.�� �$��q0�&!P)_�M�Bt��E�9�]�;�7ω�nJ�l�~���H�;j�)�[�`yQ�ƒ�RV�-����(Rj���;��<�-=rߏ�8t�
�r(����M��p��X�u_@�X}4�e�P���:�]U^r���*����?����')�l��,�	d�K�3D�)��q�cq��o4���ٮ������є'<��Ő|�aN��/�n�H�����(	����!���zz�R�ǿ�,]�p �\a*�'����n�'��Ѱ��#�C��B緊��q��Z5��a�[����k�%3,��-2�_�0Ec�!Z��2R�ns�A�����NЪ�v1�Z����7�@��1�>���;s��l��~��$]qL�h{1I�(����fyd�<���5�r�9��E�g3_؝z�.Y{�{�ʾb���J5�!��A�������<�F~lqL@1#�az����c�
"�+�2I�!��!3����|�G�< ����k�����5�3U¥�w��Lvn_ё,�s��;�~������@�2J1^���9AƥT�����XJ�*V��8?����f�з�+�P� �bt]@&Mײ���-����v�e�;b{@J&j�� 8ȋ	�=o�1(#
fZu��Lގ���+r�R#�`x"�{�h�ذWfF��>��<;WAq��s\�qh��v+�C)1�f��Q�_���<>�L�l/H.���g��||S�Ft�+��$m�e�.�{׷���`�jx1��O�����Kp!���K�<e���{�b���� >Y�|8Np�����ݬ�J* 5������!�����^F�nܽ�\���gy����ev�]#��;�}�"{:\�f<�ٿ*�bL�\l�8{N�ɺ����\ܰ�H�l���E]���^`���i����6�g�qx3���W6dm�">�\`
��
R�3��I ;�U%r�E`���?�;3#��ھ+G`t�λ[],,��oȷ�#}�����V�<�4�ˏ�8�BX.�;n��^��"tuһ+�N���,�$��z�Hk��Drh[�n�ꈭH�Ps7%���50˱:�Õ��m��1Ó�Hb�kX�[�Cc$,D�+��̮O�`t�1T��>B��9��;��jb_��G�x�b��`E��[��%�������hE}�����a�ͣ�O������J��s<�&r��`��HS`�_�6��ɯ�%AP�ʻ�`uz����8��1���*�4	՜Y���d;��CCX2��N��z�xF������uW�s4�K%'�[���K�k@:��,Ƙ��0�q�o�����5���� �B`�V�������Q^?ݺ<�8-��EOE�7�_�?�83�7�HQ}��8?�T���������]�ZU�7V����k��2�)wyVJ���2
�Q���Lhꭽ�Ծ	b�N`�ͪ� qL�����>U;X�u�XO^�	�!KR//C�ӫd�WN�$3���Ty�T#�4���>�F�-�7քDg-��`O���6@�. -�ִ��ys�ss.��+ ��uyvX2��*ca2��dTn�����0'PU�ho1�KP��F.�D��'<�CyD�`�3|L���g�����$޺%�֜�r<-��
�o-���:]��U]m��$� b�9�D�4:E̼}U�6t�3�ڏ� �K��[e��JKz�R�N��+VdR���[�{!�&_|��w�\�ۄ�J��{H�����*��(��ʙ�"h&��(�Ͽ����U~)=܌�0x�M�:F6�Ӌ���KF��Q��fp���`F��`����p1DW^����/,�d/��d!�MjA�0M�wK��#�OF(L�Sk3W1�!ձ4
�+�H�z�kZ_M�"�`m!w��:��-��=�>o���u(H3�\1Q��0��9nt��ߋg�  �f�l� �S�@uE��?�d������쫲ɧ����w6�|߮����g'y��a�8@���+6�D:��c��Pk�Ao�-b���I��u��_V���m-z�c"o��=�)�N!�=<{�����o��6�G.��P��8��I}�jhJ�,��zd���Ɍ��(	>�34�&�T��h�4寙����I�O��2����c�x!�[�++0��+��H�l�9c� �ދXū~�S�qic:0}7$�N2��0� v�m�ؽ�?2��Ѷz��w&ts�)�%dcqj�W�7�N��ۨC�����W�e-pl�7dǣ0����Xr�"kk�3���1��O�<���b	�-�1�u�a��W.���7N�_(,��U�N}5�9�ڏΊ�Y�韰��8��E��Q"&�Ϝkܨ�p��t�V�A�-H�Q(�O^?".�m�|K2ZRp�ZmJf}�z<�D������_�f ����A��Ц�QR?�k����K	v����G_k�j����n��a�C`����l���<�����2n�cl�����qH�7gĀ.���^_I�F� |Q���\.X�h.B36K��������6�+�&����ز��6e}���]�)��K@g���S�m�&�����y�m-K�V��T՘Ƒ�y7g��m�_�q�J�<#t�$a�򐡅5�m�B��@8y��(���\e�O-�����.�5�XF8�"��I6�b:̇Ϳ��3�/���O��B�Cj���-�I��wĢ́�V��惠5Q�N��{<Z�b�-I�s�yv?�{�3��f$C
��!	��d`��v��.j���=�t�����4�^ݳ�^>��}I4r�јr1��-+��IK�H�U=j[��c�1T2���_� Do�;4���`��b6�ݮ�^�|�!_7����T�y6���7�9W&g�) ����g��;��Un4�����`�2��ј�h&m����Ӓc�{X#��y[�
��s�m^�����BKÖq����¿b�ڰ��|�����X��Ӝ�3,�3ݨ�b�����E�2z0���N��U!�� ������-� z����f�B{��}sno��5���_,��J[�n��9���-��s�g�ߓ6�趁���MF5��3K����!��h"O��$������9�eW�M��hCվ�/��s%�9���#%ܵ��_��Κ�pN�Ei�
�n!��8߷z�.��ǻ�)}���*�v����䲳 ��x����?N,�)�^8h)ϕ%�T�t�Gs��41!�FbYlA������x(q�ya�t��'�t�����Z����Db��kg��.8l),*E_�
EUo�hЈ5
zH��1�0Jx�uɨ`-E�sq�����akc��}{��sf AnVF"�6FS'�~���l��E�k�������q� z琠��'����c��'-9*��r���Z�I} d��	�/4��_u<u.B
�@bڬ�Ͳ���m�ꮭo�L���\/U��<� `��C4ب�/�'b�!F~�o)B��H�W��=��I��fv��b���1���F�8߉
�n-��ٶ&��M!�٣P)أھy�3������\��UM�f�F�o�b�
��T�^����*�ɗ%�Z^3�Ø�Q�|I�Xӥ�~�����} �V>lK�{����wGZ�<�m�Dm%��!s���0��a�5�0���4�;�,�YZ �8alC�����-]�yIÔx
<���-)��
ř\���(|ւ��HH8d���n;�1��/A�b�&�4���Z�X��xW�^ǋ#�˙~�I���Ϲ���Cށ`P�;Uݑ��%�Ԭ~^����W�!���L1��ۮ0Q���t-^΄��X͔)������^='V���]b��c�)*��?�M#�i��y����<L�="d�ķy;ȋ���n�$IV.��2?�Z` 4y���ñ����
������6�[8�����K����k?A��5���s�jЍ�>���4y��գ����uF^4zN;+֖���5���F�@�^tį�)Π,<r@h!	|� ��?=4�sNÆ���M�B!�L
+�b��îo뙫�>(�i`7n��Bz<(����S]��O�N��c���\iLqB@J�E�f>��Q�ld��{Ȧ���i"u]�c�O��R.9c#�c���D�'}��(3�:Ŀd4(���9�F��|I�#�ܫv��
�\����`_�y_��Ne�-�l5�v_�Iƣ�G�uW�E�>�/&s,j^�8_���������FA�� ��
!���\V��F�;Jm#`^_7��d��-�Hk"ڄ���f��^�����"�����P+NI�^�ϒ�j����,H��O�ќ���b�1q��/��%sO�0E�R�Ɛ�]����T{���g
����?rE�E������|E넟M�l��?��|s��Gԓ/ũU��9S�B:�&c��V[v,�(�F�?�&�1ʄk	Vϫ[N���.�l�}�_�˟��%�`����DǑ���#s��Z��e	���+���5�<����%�T~�D�b�-���uj���-q{ μ���d�t��L�p>�9T.Z�� ,�n���o���?����́E؂>	�`������~��/O��ؕ��]f����`�ǈ� E~d~	�}����P7�����h�����Wq���F�$?�Μ�ˢc״z���S�0[ 
�1@���JGWF�e��08�G���~h6��3�Y�ӄ��=d�.��+�9�.��T�L���xT(�_kb�]�K3Ւ��n�i�u���	(�1�	��sg�4����T�e�"jS��j_��j�2��C�۔tW��� �C�j<<O�m;/��rо��Ğ�;�F�7��#ǂ9��%i?����}Eh�>�&h[���� � 犓i�3�Y2��>U�U|B�����E1���?ʨw�,ڜ`�o�sȼ��Yn����7�7�Z�K]��ѷb&b���Oұ��ۃ�����4(������3���[��
|�J�j#~'���dK�B=�Cw��#o�)��th޹�	�C#��%��U���z����,���7"뙅Q�4�C���E7;�!U�F�dFt�B�]FՂ�U��>5�5�^T�GA�X�~wcQ������[?^2�)�@��H-�	*<���vY��������[��x���7ݴ�N��f�0�{��Y��aٔ̔&��$*TGe��I�g�/���Y<O�Oз���<%�H��ߩE�<b�G��g
Oc�qu�6a-��eb�ذ��E�qʨ���Š�\��T�%[�t�zGR��
�4���=B�D=���#}��_4m�^㰅�R�IC���jg����{�� ���!��~����������D��|
<���#,�-%yx����7b4��c\<�?��[��8���(��VH�!�< p�����T?�c�w�0�vC�ʌ5l��sz����� ��e�ݮڕ*�x����QՁo�9��`���*�C����F�@���QՇ�_��L��)Wa�� OhJ3dUPER���*K�C��%�8_���ʮlC�A�ë��Ɯ�B�� 
�����f��,��<��ȲAL� ������1y�t�!Ѯy�_��	cp���%�$ᤇɣ����k�y��m1����5��Lq���˅��2I�k�F��j5��Eg�#@�'6R�@�2PN"�9wUa9P�kG+2�w��i?������2�f3]!���ZT�+��	�%�N��HsD	�\���$���Ð�����<t3��({�4�y�e� PN��� ����3}�@ƱK7�5�Ac�
��Ci�ʫR��)�eT4���M>��:�@�H�MnlXGYIbm�����\H� BF0	"�@�KK��)�!�i��{;�7���3����ʗ��0t1����@�2����{4u56O5yi�6��<a�+��<��3��i��rY}�2�:��a�nʇ��޺�Y����Q����7��Ɂ&~�t�}e��_��W�7�Y�?洍�}�	@�����zH���	Z�7n%l(���_~i���q�;���|��v~��5
�ga�u`4da�1�G��D�l��<����W�kW��c`��F7��ő�8��凰�����SQ�#��u���J���H��g�?��7}M��H� 1;k��c���Q<LŒx���K���Jz٢p�eZ^K��P1��h�|�o���D}�58�dRi7�R�6۝�3K���O
o���~"��&=�6?)����?/\"5,�k��)&�#!r)V0�͡�I�UEh�:��Ò\C�3��	`OA�S]�}�0���8D�aB	S���)�rv��ލ���l)�HL�6R1�-���`i�ݴ�{��Ȓ��@�`!��(I�9$�rR^��(�A�9"Q2S���o�L�n���?'��l�cy��=�S�����YY�gެV	�N"�&f�
�׺(�PN7$y_�w;��i�ϱ�)���9�h�B��3%�����ʁ"��S�$P��Zdqs:�X��o�U�H����c�d�*0���¯�w} i���!���j��g���S?��r�] ��?I�W6����ۏ�1Z��߳����pbdp�e�M��8�Fϲ%�O7ܽ*#,r��u:ܮv��ɝ+�FWr�Ǡ=����m;�k�7�0��A[�w��-v1t�o��Օc��+/Q�ٮ`� ���e쟼���h+M�=�ڶd��C�j�٢� �<����ͮ���� �9'���֣PUζFF��I�A�����ݢ���]#���Ri�8�e����ޭ�}Q�����I T��l�-G\��@$T�:r��f�sb�A��ީ_����\��Գ�w���p�p4Qa�U��^5��S>]�4b�:���J�����]aW8���t�	m�c�ug��9��y��:�y)XJR�{��&�����K^�jdx���w�
��`��3���r_Ԝ_
�#|h$��l֟_�꓍�e
�g	�_ȏ��P?���E�Ƨ1xj.8�t0&�`�GY 6_t�Q��F��O��S�>�(Op�B^]w�L���5���@\�wq�3��[[�M��}[�Iz'YbSwD����W:r9`��:-m6�8[~��-9V�ϫ�j����o$��س���!�����ѭaT1��6nAf�7;��7y��y� ܤ�H���,|.o<��H5N�DOg����/��T��&ֱ����L�AX�(=ٔk>���C�=���![������A N��n_�� ;!7�����>t�Gr:����u=��LF��7���w/=Ţs_�i�m!�X��N��J����FnvF�~�s�[~��`o	:�&(ݥKM�9����|֦�@�'��ޅ��,m���~���hZZu�!�{�oX ��нE�I.�5=x{���=R�=ٜj�0�G��sf��O]~�?n{�aU�X�ӑ�	ʈ:��
���j@Pj ʇ�v����M>U�)	����4r�h������['�$���#N�xb�`�pqӡ�p��S��|��j��1���HFQ��Ae(�^�㘿�H�Vo��i��8y��ji�����kRu�{�d�@\�����+��X�6e�Z"0h�0S�eʐ����h�	�OZ�l�RCR����ߙv�#B�/t|`}�KŞ��9c�%9|<��%2~�pm�iG��/:�;���|>��Qm�hRE�W��@\�5�_�h:hS�W$�)�$���h��we��à�.����!�!��B�~����$4�D/�a, -����f��%�:a$ZK��y�p?�7A�ٙ�뭎���EϜv~��_ʻ�	b��������ڙ<ޮ�f�B�
����O=�����-r�ГV[�}���ey�%S�f?V����h��9���ן� �S'��V��͛ovzq�tV�[V��������5��bfO�H�h 4s�����0�to�IR���r�<�b(eF����/q��tx}������iO����K�NՓ 3NĂu�e���FD��]��f�˒�F�m�^7:���BTj�4�im}��򫂃�C���`O}�E���M �y�&֨U�}ToȈ�qP�J�!#���[��j�4�Cc��/<8�~�]˚c_�����N$_4�-9������伺ڌw�z��`�
u+N����Yv��۾���O,&�a9q��)�"��Q�����-EYP%�����B�
X���5�}��D��VF��F��AT�� �d��E�<�K��*�e�OQӼ�v�㢝6Zaξ\��h�+��b)J�'�o�^*�?/ٿ(>Њ�e����).>��¨���˺�HOs�u���0����b������>��
F2��&��b��"��b�|��h�ކ$)zV-�H�y�ջ�n��"�*ot^�|5r����3�8<M��c-O���H �]ʉ@�$?����l� ��In��u-�����⛲l��o�.�v��*~�쯣L�)KE<��V8
_���E��
 ͊wVP�&�}�ci74�t{�Q Zܔ;��~��-��tUt�<��<�C_dE�i}�z+l��l�sS�f���kA�u�J���s���� #E	]g��X��)�,7��9��vv���b�7u��킫ɺƞ?�l~z.��>���/dE�*�l�E8��� ��i��`���98�,��}v�!���G��9Y�L!{�ʼQڀ���e����b9�%���
��Ed���B�D;��&'�)�s R�����_��1Ԫ#�'e�� �\��sz�9r%�R���j2�+�,nf ���S����<���OV��`ag�)խ�v�m`"�H#(NdW�V)2�2�(>P�B��J���:�|���'������W�E(1����l��%0�[�4#f|���f�[�rQ���X��[��R�.��C��Td*QD#�@��bm�M��|��Jg���$N�X֫t�j�U�� �tE/p����$l�RJ���bX�9k�lp`wǌP���غ�|��Bz�/ħ ����ѱW��:���݃�p�}KT��tS,�	��$�}2d8�����s$���IwR����~��i(��r���cV ��c����a<Ϛ�e��ȓ���=�FOP��7���2;�v�
#�G�v��~�^q�vE��?�B����e;�_}n�z��Z��3|�r��\L�0����T���ތ������pf3p�O�����9!��1Jq�JX�Rd�,���t9�^)j�Ft|y�c��;��x�E9	�����(��A[V�fO(%PC�w�̪b&u�2R��-SF{�!�s����/ӽ�3��}0�b�j��CQ�vu����PB�Y����(Wm����m����~�|��$您el����K��?)ΛI
�7�$-zu�:'f���3	��\�znjo�	�:�JO" �?���8(mK��s��N�O�wu����ivL�Q�O)�Z
 ����M����'u"�l�.-8:��>?6�t5�7��k��]���j`<�7ϖ��:sFi\����X�kZ�tk��l��E���s�j$tq�o��kz���i�σ��|��Z��>8�"J��)�G������0�n�A���	�G
�LܿAF��y���`&t���ok�(ҕM	M;>d�x!���4F>��Ĺkߵ�~�
C!�ٖג�-툣d��E:��h�Ó)�Ջ�b�|� m�(�`��:�E�_�|g���{�a�
�� �]�4׿��y�e�<u�}l����En��Ig�/t�'���\�U�sQ�n̘eG�,�?L��0��+ʂ��I<�#��[�̬[��_.��G�2�����FԘ�f� 8.��:߸ؼ�QBk�/�ya��������9�(���Mb'�N��]�؈L*Z�]TS,�fV�EmL��fO{�^Jciư�f���c̘���69C?��`����!>��"	j>Ǧ��!NL�o������=,u.
�pF��	~�Pc[i`�eqxКI���b�Y�;{5�MV���GU��IO#�Ja0���Hk���Ws�$����*�x_aa+�xE��xw"h�;2?{���i�4�e��B����C�i���o����|��7#f�L����U�\����n�K�G?VtSYg��tX^4������Bg���w�=��;���V�L�m9�b�%�*&��%v��I��ڎ1V����kn�T2�Ii�{��]�	m���UU)��c'~ ��������5K)6�E��[z��K�CZ^���pv�U�g�׿&v�e� �5c����kgB����d���u�D��G�O@ <�kEH1HT.�kR�~T�-�,|`��0��E���d�k.�h�?�	�C�%�  F��}9��3Ņnp�!���\y��EyA��7/�d�sx��z��)KE�W��Z��@+��bmS���/��Li����yqP��4l T��{�3�Uu�KZ�m�N��S�dל�@���|���{w�ۣ��+e��$�ڎգo<��Z�SȰ�[�:3�����:D)Ƹ<��Ea0�!3�;�Jb!�c2����"�!%2C����^�����!��.�zMc<�հ���)�NPӘ5�S�3�͐|´������S�V���e���λ���]|[�ށ�6O=�gh`�a$ ���Y�&o
"�\Q���+�����qQS���U�хh�LE~\�}}S�����h�xv��. �>ͻ���d��Jb�m&�˭��s�C۴-L�$�t�l|b�!v�L.�
7U��U���6��J�f7�N<�mzda��<4b���q��QQ��, �2��j Ƅ^)|� ��F����qg�Ϭ*YWpK��m1��.����� vʪ��]�8?c�E��`�� �٩˂�����O�XN�����~��?�0C.#��c�	.��Xou�/�ೊ����p�VxZ�,��ja�C� p}By������w���Х��C�p`��M���M>�5���u*�-p�)�����V�=^8��A�����=��m��(���7t���S�t]��Js��#��w
�)R�Ͻu�m����X�J�CZI�������1�Z������\ue��$����tty�7��k�X��C���"�����to��͍�	��6^e��6NG�V��B}<]y+�mz%5�^?��sx�ϕ�e�IA�Xd�{d��E�q���ì��F�9���H$�e���%�.�S��i�I��3��Z6�UU�9ZD��1�l��Ti��w�СFR�!�W����e�T�#������ �q�)~q���	J����'%pP�}�xn��J����J �!}PPy<b_)���~�t��U�����m�����~�����U�Ť��-�Oa/�J&G?��,�/�F��6�+��"&Y�ri�ٴ�F��l?��S���R4�O��Fo/��`Vc��8Y[J>�<�_0��S[Wxe�ZYR����������� $�v�ܓ�R�5�@�F�2"���r��������"�E|��b&�N��:%i�@bA`�Ot�@>�0NMyc���-���6ʸ�oܳ@�'N��/$�i�o��_�P���hv�id�0�J�(��vՠT�k����ڌC�I2�$`�ŐEQ�@@Mb1Z=�,�kpX'�⚞���"��<��b�}B���bt��$��W���_%�ÆLU�d�{}aF��a�ܖ��}�0+�H���x�xR��ھ���<�|͢�B��H«���5|q1dz��H�}��!�	�1g���O�?ʹ��Π�.��>�S��ɨ\��,�肸��S8���Ql%�,r����2�X�@�!/;��(%i(�ôf��ܦ�qJ
	x9���dl�����v���NLg�!���w\��g]�A�s��<�ӎw����SN+3���O�B�L��5;�@B�S�kz��St��{�p���u�"�G
�qԂ�ho��4�6��h�r*	��?��"��[(G��JR�f�%��D,_�����T�:�5��(����M�|D)h�)2w��R5($��n��Od)za���N[���T�yh$k�g�x�-��$�oL�ZQ�m�5G���(��i�⾘�cl�Fn��z�=�#I�24��߁]��PAG���}$�<4�I�����([�������N��*D�=�_��y�߄���d~dI�^�m��۞��2��E� u�������CL�C�i.:��3%�[�Lf���7+��?8S�\��"�w�s�k��FkT0�2����=������ϙ��1\I5ijU����u�,�6O�˧�b6��%�w�����T �(��x�r`�X�*�[�)����M�3�4�ߙ%ס���_��'�H�H�ޗމ�5�.���B�q���&�z}](���	+^�Y�%z~_8�ެ9i6��(s��˻d�h��'ֱ�c���
`��r�S��R&;��!#SO����qHW�Z7~����=p��Y�[��e��7X�1#��pn�Ѕ5N��j�[���<`��id)d8�
z�P��%��Z�(,Kɕ�I5���
T���/WueP�,!jH �>W�"����}��A��s�� ̟Ծu�N�ȱ�F0dL.=���C��;NH��:��FS 6���%x�#��$�\����ͷ��2f�m���FBVA���n�Su.��݁E�ε���j�.�2WiU��g% TCN@��a�`Cܚ��۪�&%� �����S{����E�s�uF�!� \��?4S�����\|9�������@������5�q(¡$��{���.
d���ȁ��H[S+����z�<�ө0�߾�U@n�`����k��d��:|�]E�b�
�}8W��z@!�=��n���� �["ap��\`�fKZ_O\��˯�+���?����ɐ@֑)���@��>��Q	es�mXU;�^2m�8�Ѫ{���;R'�U��՚nj�>OQ'a���{�7�Cni��v��@���VA�ڲm�J���~*�hJc9�q޶��A�SL�H�vĩa8.�����maE�Qy�Tr�'�aY2���c�/a5�j,�k���whs�<G�^I�@(|&.��'�nM_R떦��/pq��*zF��"��(�ԈƦ��� 8��Fp�[�'���s9��Do�d�6����*7�-4�g)Uo�:r���{:�O0
0�
&!�0�x�t��_ ���I�0W�9�L��/RL�v�����!?X��evU!�Ǉ�pWlOu3��+�񉻥��vas���\�a��X�0�L���Ż�u4Ԡ�΢S��<�yk�1_+��즌7?�hm�֥�[�A(���5b�Gb�%yYl.�
�4 ݜ/��걚[i� �S�|�,ܕ�4����9I|Ph�ĺ!�#�j�;��c�Q����su�<�r�t.k�;ۚ����Wwjc�;�)6%����7���UH��B}�(��^��'B˷�#�O���z����[��� F���0��Y�8Y�@�&Z�}�n�[Ba�R�P�&[tS�#����Jp$���c�)����	�dx��BV�R�
�w9W.����a�0�R���T�Z�?;�p֗��M����ڒ"S�T4��C=P}�` !XZ�k#��(�J�$b&�5P�m[�;G+6�\�� 6K�IK�����LSz�5s���;���j���_YM��(�Kd>�ۭ'�G�fU�!*g2ҹ��Z�����@�b��C2�4&ɌjD��'2e� 2ߦ��5 	��*U���J��X^\n�3����NC��q��B��V=%�yw/��v��؇�#��8B���<v��6}4�����#.|���aد7��|���z�N�ZYgA[���=�1��u<���G������[�+��=ѭP=�u	ȍp�����G�:��5\l������Cu��9S�@rkΦ� �8�\"G�z�o��`S��\���|g&�pg�g�OA����2F7���evp(Lw�3�=�Yn��&灀�t4��G�Qou��w_g�_j'�Y$����cxq��Кǲe���i��O��z���
o�h1�ҾL~���IQ;b�r:�UF_�4)jO{T��`�f*Ip*o�E� 5�� Κ��[������#�N�*vy�h�	:�G����>)�{�Л�'[�F	�S�DHaҨ����-VFۤ�y�:M���t��g�Ͳ����+�%�K���'xʨ�VN]���N�ɢ��i�n�VeOnB��`��W�J�0��\��W���#��Je��{-�l���x��@�\P�:;dO�fQ��Hͮ�>J��Fw/��9\�J�}����3�n��j�'"Z�x�m�m��NV6�~�p��æx=3�"r��]m�71G(A��|��������ѝS�o�
}W��f�MC_qڭG	���坻�ѕ��H(R��<�����U�qW�5V���Mا���+�ɱ��F�f����ɸ��_>�9�F���b1刺��8]I�+y�I�z�Ƞ���()�'*�-k;!�4?Q4ڀ!��,��L:\���0�{	j�)�Y!s��-9�x�|� a��8R~%I�Jdk�9 ��C`p[��~��I�����3gȐ�����	Ϥ�f�8C[��>�彟n'.� ��a�>����|�}/�*�Ί$~n/�]T*�N�<W�zYnԊyg:<�t���{���qn��^H�ӗ�*Ie���
�����_��`R�?'e^�:���cA!,2��|�K�v���e�x,���.VvVM����=`K�{���jC
,(�*�x�bL.�bidn�j{T(�(i����׋�K�Y;���t�!_X�o=�3���Һyޫ�@�k��Xӷ�]J>˧H-���<8�.�4�T�U$UA&
�XbW�m*��F�|���Vk@�3��N��� �T�#�����F�a{"��iV5�(}^��#��s��0R�X,��\�_q,+�w�=�cFe��L%i�3�X��i��T��O�%]l��`]�s�2=��ak��� ���(�|�A���ٗ�$�Ef�iɤ*���c�ˣ"�/�tI��#�@��!re�⨻��A=p(�vZ�iO|RW�+�l��ʥj9I�'�c��|�ơE=��6X��+'W�����pk�O��[�w��R�P�ߜ�G/Sj��D\IA��I"TJ������� �xJuk�3|%�X�
���a�\�v96���$�`��y��g�!U1�Mm��%�ڎCS/d�cK�I�.�����ׁ�K��`B 	���t��0񓧐Í�M�p!�&LSS+�ǨN��� ���uC�Eg�]>�e5<�5py����*lû >s������a-���B$��Ǭ�� .#�@.Z�n�(�)A�\�v���Ob���D"Ÿ#�SB�ls
�h.
�Nѱ��DL<t��ǉvV�2l��N$~ˁl�}bK���	�f�VhV8��C�]}��8���j���T�$��1F�@-�zzm�����ٛ�����!���u���sƵ�����ô%|�e�r/��ܮ�l`��������k��d�Y�=��e�*Z�e����	 �gr���QTzy=7J�k�a�p�dÐ����U��r'��{���lȜ��F�\ݾ�vCc�V�|FS����j�Yn7f�����Ź�9WI{���@Z�ܒ��c�#�lƙ$�/p��1�5�ߦ�YH
���=zk��@�ω���U�{�fI�E%l|���E�G(еQ:!��3�?�c]_F��aJ����4�Q.����ZĆ���"n��d�*�o�q�:j���������-y�V{sӅB���Ǫ�:������zI���%Z��!�@���-�ת�κ}U��8��y6��co�mD�L�`)���)B��b ȝ�Vx�c��^z����xf����Oʩ�z�m��jb:��M�*������]����oB"�g8�HЧƞ`����֊�g�[ʜE�n��d���-��39�Ĩ񜎋>s����1~�eBk�%��RefP���)��<�]����z��c�Y����������4�o���h�Z$��郡�)'�5݋��/�^W.	���� ���s<Jd-�[g�Wj��^R�C5Z�+�P�Xɇ>'�PJR��:��yz�烈��FrU�m�6�rN���xaGB>��K�0�`˚t�XYi��������#=]��&��w���M ��ct��b��-�l���gy����\�l��'��6�e���"wf�k�΍.Ӫ��b��"�ܯ|����0�Y�>��|��H�*YX��<����j���-Gq��􄷑��z�|�~n+C.ա���&b�f']�4<���b=3���O���l��n�\Έ�<ODʺ�	 �C��Yyt���̥��^�ɥ x�o��.Գ�=���
\���`�K	��1���7VJ�zI���q���S��ב��<���`C��J�УƜ���ꏛi<9�δ�3X��Vi��0������U_�~�G���u����9����28��/��~Zkʭ�p������q恒C�Z0�vD��!���`��T����D������D�<?�������܃:��R�9}NK�QY~̈́���G>��Yʮ������x��g.�$c�������p/�h��8�إo;�ë�5MP��o�0T�j8�L���%֝��Q����E�.�vp��s�0�?��Gi��B!������&�(�i�&��́�᪎�W6%|��Px�Q��%F>��0��R��
<�����-M&�ß��~HX�T/Ǹ !9������h�[��{#�N�����c��� NwM�s���X.Jy��%��ߗ�t�r��ַ��5cL��!Y�=�q�u�%j�$v���ӻ�T�h�\�ü9F�B� ]��ġR�	�	yP�Wޕ;y�g��HC�r���
4�L&�mKj��?��-V��H]���Jc������- VR�8i1*X����aKA�)����o'@z]3�(�.�'�v�znv��:����?֓:
��E�K /������1q�FHX���b�U���>?�+�:�:*���Pf�U<����f9)�e�p�٩Y7�K(ҟ���^^/�ϼa��h�v�h��R|�e���'�J#�c�,��c+pG� aӷ��ڦ�4U�`!�Wgփ{0UR����6��@kn�����Z!���a*%M,�.��͚@s�l�g����ů-�2��y�dIv�X�D��_�.�����>�|~ū6g�_��_"��=�ɧ���G��h����K����A����n�<#��} �n�q��┊���etl�zikt/��3�	��=M.���Pf{�Ep��f��,���镠��I���&pR�vd^�r7��d�������bR�\к��9�V���cE���oƫ��w���gm�h}^��+/���O #WSrW�~�?を�-���Vz<�W�W#��C�q�No�E���=mW?LA?ߞ_7Dʏ���� �"<�^�U������O�e����q�^�x�-�ߢ2Y�U�A���V�Br��oib��g@�Y��c;s8�؟�٧
�5j�
��G����є�CmI�%��.�!�z�Ro,�7I�w����o8J�Z�5����$�E}-~�>.����9�B�pG�V�󝽏�E�`�`�QO�ME��B�T���{ƒ�+l�#?���2������|�r��`�8%�|��i�I3��c�C�
�z7^m{M�_�z@f�҂�H�$7_��5�k7� Z�u6�/e�@k�ٱ\���b�]>���+� �.a���ܫPޣ2�@����U�F����5Z57R��$5�.mъC=�G����(�2��Vm��"z��]���F�J�V�� ���K�2R���uÑh!г6�^�}P��	4�,e7�Y�5���_!�Mu;�����͜�T,���2E���/�+YQ �n&c5����
<Q����GZ�8��n`3�93�Y�L�$���"��[y�8�JQ^O����F�_�%��aEv�*]t[������A:�ti'���h����Q�dz��u.�&��-[L:��0p��Vj�2�P���ma���=��ˬ�;ʆ��L������W��I+��w������ʮn��MV#��}L)�3��h���pBu�l�?�f�OF�7v�6�����\�
jZ�ޅs`3)CV���T�~�*��re;P9b�q���ߠ���l0���YQZ屆�q����GT>GZP��=3������lq�X����W�&�xSj��{�\釱׉sŇ��U�������gg�_�u�]����`~,>V���P�+������)B�!e��Y����Q �ѓ�g��?:Ev� �a`O�i��B�n��m haz��[��\d$|@�͟�#?�o1g�2�\��3��uޘ7��YU���&��Ȁ��`��EYptS!�y��r�s��Xu��L��E�?�{���df�����pԦiVEPa�����5
-b���>�[�0PD��ă�|S�#���z�mnׅ���q���5��$�[
e/�������@�Gȅ�&��[�aM(JC��W�������-��_�9�:����"h�\AU��i�D[�p�K�}ju��(Ck���o� �^�x/��V��Bf��4�)g�SF�Hw"��U��qhfɨ�mmM�~պn��x��/�H4�Qqɀ��Y�goɟB�5j�1�B(`)xb�H��� �a�\:��F%
�'��^%�j5��ܨ�A�����)����D��F�����>!Ο���q:�ZG1�^z�$ca]}�ض͸O�=|��Z�=���̔ݞb����.�4�b���6S��F�Lz�f�F���(�K�1#��DކQ���!h��@�:��{ET�ZS�ٵs�Ze)Z��SI�^���N��+����`����=%A���D36���g*��3���u���)�d�D���\��;�b�]eEHFʎ������*�-�x� h��4�t��������fp�K<���Q�h���'7N���@uꇂ�������ʠ��eҗZ�p�M�U�~bړ�RVZ�/u� 6�&��G��h�C�*�I�Ht(+���u�x���T�s��#�&j��K�[4Ԃ藈7�o��a���fł�T'޿z�F�W �^�Gv�]j�1�p:�j�k�Î�
��e���aZ&'��%A��k�\s���Oi�Q#6dO	刬������P��v�m�(�"����G�<�jI֊���1es��4 ��=Μ������v��I�qz���y܁�۔䮆���M>�[)͘�RH���ۖ��	�W�bHQ���M0��n���YB�*�b�X�������L	(lK+�Qn��0�M� ��b:�2n-� !	�j�eG�@G�\��v�p��-7����=�?J�E�C�s�:?ˢhe��h/��bk�a�a��" � �&,O������V�`�6N?�ߙZ��^?k
]�
�!��s���G
w�hW;�(A3k��i{Q���ַ�)@��k��b~�R�}\� ����x���:y�����
��f��(����~`���Fl6�jHf[�w�Pu'ԭ�������C��B� Ű�oIo2�'�5�K(�,:�}��-�ww���F3-�-����>��=K���7��Z �Ҍo8M��hfh�\>Ŝ�
l��ٹ�^0@t��ԑb�ѡ;���9�ݍ$�׃��mCX3�Mu�'E����"��m9��׋�{�<>Xg�XK	~�e��,m��[�Ob�M��MǕ-�#�����]f�&�������>�M���<:X�uE���R�Q!�(���'C��l�IC� E@T�{���M��RD$�yip��FY/����E|�j= �̵V�lvr�cÓsF>���h�����s9E&.vd��~�Dfo!4d'�}����@?�yD����`��'�16+,7(8��"�,��<����ꞹY�I��N{���Ί�O�]"Co<�Z�޷CG��o�� :9�Ja�9�P�^���{o�~�����1)�9/�c����ޏI��{�����/#��z�S��ò�~�-��� I	E��&�đ3�����(,���U�}�.��!(*�wF�Ϟ�S�ǂ9`�Z�o����T���ש.�m� @��w@��{���!0��r���g<�{�׋��vdN}��<+˛�s�.�mr-��~4���C�����ٖ1��u{�B*|��Q���p��v���y������熂 ΁�7�(��TrF��j|��ɯ�EX	�Ψ��tf��%99�Jh4@����/x!�TI����3����5:\h�0@�l.�~R�I�M������@��k*,/���亖[�4vQ�&[�|��mJ�<1�W�;� ����"��%'{�5mg� B��`��qv���խZ\r?�H�͡+M�NǬ��RE�6�j"Т*S1��}�'��ޮ:7�g��6g�딲5zUC�8����k��wx ��dI����:`�<6��'sˀ(/AB��� ����)��Dd �
 @TXX9�>�Dwd�V��X�]r���Z0��#�Ep�/N�A�=b ��(Vl .�E�_��_��D딊l[��ď$�x����H]57�W>J��||�� �F6�V��8c1�
q)R3�@	�E"r����f��Zm
]��=�9W9}��S�SX/���a��
)���(�;ZnRz9������sz�� PW�� �����Z��MKVf��Ǹ�'F`�9:A��7u�4L-|��kԈ�d�g���E�~�<AS�����E��"kk�ˇР�������dU�z9�˴�YMΌ�	e c]Q�9�GNS�KFn�ڪ�i��lf�A�a>���BE��)g�˼EL/���8�����_6��=.J�O �v�Q!�Ie�&���&G?~�:m�JԶ$wоUm������x�X�V��ʦ@BѸV5T���7+���ǰ���G��tC���u�_lb�m�+u[�Ao`��)8���P%�nz��\�T2����$K���k�i�= |��B��r,HGZ� W��KP[�վ��@��m�:v~�Ѽgxe:#^�X�	��f:��bbR�3k:5���2!;�! ��^�]��۵�w4B%yr%<�|(x�xF�Ho��C�w�$j�۵/� ��dx��5
�ѫ�`�~7>�m7C���uϰˇl�Kj��f�<�(����p�'3H�>m��㴁���H&k%���I|fE���X��������!��0=f�5��`�-�WOm���o"z��� V}����5��q�>��G�QD�4����W�:���,�'��"���������'�dT�������p+\�����YQ�b&��J�{���:5����O{@��(;��LM~'0�gd=��j�=�:����CnE�
��+�6B�b������##%HFD�HT����@�S5�a��|��*κY;[� ���ի�c�)��_@ZCt����
��mY:3��ŗ���q`�'c��ܭ��xL�o �z8�� "��a��:�S���<�d��cS��K�6�q�&�����=Ut睥��!z� �v���gW�/R���]~ڳ�^w.�":T�Rw��U��3gQ����\� ]�I�?H�
U�##�����	J��W�_d��N� 1?�j�f����x��1��I���ޝ��2��w08�*Q8x��R��AbP��幯do��7�����%�Ü���HO��YWƣ7��p�M����מ���
,=�ˬ��n ����Ro3�
֬͢g�r�exh�u����Hayn��
��Y��s8�ۍ\�؈X(����L�S��&��-�n"�"t�--�'�jr_� z}j@8!31�_�%	�9�zR�+��qY{���J��O�t�Y��Ϯ =н��B��aFc��78UD����U���E|F��i����E�g:{ѝ�Z���o����4��t�
v�J���XmQJ���*҉�Cm���`��˱_5�z�Π��L�Sj�G���+Sc�Z��@7nE�3���^k�V4�:{^�arͬ(J��~�A�I����G�~�ϙ4���a��DA���*��C�M����q��{^�>��b��QQ�PQ�i�����ί*@+۩K{�(+2AB|�:����TnF� �n^��g &�R��h�9Һ~Ŭ\�?˟g�i��k�{��L>�b�0)@@� ��	qnO��y���,{����ɮ��B��S�Ȱ����}������x�6��]��yh{�(ר\/kU�Q��+�����dPg�w��a0��A#>�,�Ʈͯ�N!jJRb��%2��ڊk����p]�pud9�)Õ��z�V�=��<0DJuqV�	�ˌ��,,�W���&��Z*�q�����21QH!	��^xQ�B�O�A�b�.��%F�_��麶��O↨WxM���ݷ�bݽ�Jȱ�_��Zs��K�� �J�zݰV�JK
�|����~hc�bTK?bBLB��#2>Hϩ�ܹP]B��U��q��A��fO	ä@�� �Ɛ�sw�|��C���TՀs�S�'>l��j=ZU��}��@�� ���?Z�*�Y:�w[G����E;�Q4B�j�08f%cg��tg��U`>��*�{�ɞ.���)��}�!����:��x�G�F�?��=A;&6�fk=�e�$���Z��gב�ad%�W�'���N�F���|�B5�q�|���eyaip���x;}@f_�SLᨍe���G�MK9*W ��nG�ᵘ�^l�*�7I,��&���ܦ�j$ժ| 1�t��}C�WS���L�׵�@�hqQƛSт*ˎϑm9�ۊ�ב��?��x����8&����+��n��)��S��H��f1�u�
PL	ư^�P���
+�-��>���	�W�*�Y�>(��q�=a1qR�#�P��S~�b�	i��!	�ɻ�0�)�z��2'O{U�|m�tއ��>���J�p���v�>��'�L�WT�����tx��?�vQ}�,U!��V�������hL"�([��������QS����qp����<��*.���RF^��9�*0LSN�K�=���W�ł��1%#�3���͋����A@�+���l^�&��"̢�s��Ŝ3�C�D-ա���O�2B��R�m ۦR^�E���*��1�EG�A�����W�O�;�Ȳ��:�ws{m�&5���mP1��B�
p�%P��h�A��f)��DaH���m��Ž��F��P��v�L�XkmxeS��niD�ُԣ��q/� �ň���r�6OU�R���[�N^,/�D�j�Y4+�ϴ3�l���-�!{2��/��\����^|Y��6q�	��u �\Cl��>�$�QF#gv5�F��]>M��N���R�_t�?ɢ���]���NV�7�H�'K�&\a^�ڴ�������_)�HB�"c'�xNPc.�٩�R_��y�br�泴��2#~ֳץ]�8,m���v;gR�~��b�):@��U�W�E��Q٢��'}����o��4M]�[��*��XB7�ӍI[�!�.^�8�zk5��T�8��įW�����Sᚔ;��q�B\�FL�G�n�{�_�.�=@��������i�P�݅{�,0�k
u6	����֕	GI�w������+怟�j�����j�N"߭�eH��w�_���
6�V�3�:�ԟ��֌�0����B\KP&�^vݙ��ݒ��dpز���wh ��w��`������d0�?L��;�B�F
fVXՠ�Ưטμ��#�IZA4�ቡo���=�4^��
h{�D��dQv�� A�n?RE�m?�[tײU�o届m��H�z�Y���n-!��_�'�J��	���tK��\�b/w�f��D�K@5�;t;,�[��^N4a�R�tU�e�¢���M��ׅ�����\If�����FK�����)w.�1�5�M���.LE)09Di2��=F|�D��l��{y�t:71��j׍�$r�_0�eu�A���Fv$��<�nU|���1��))fU�Hs���)�7\�n�޹7���(Q��l�H#N�3�Y�:���mr5�	�r��=�1�U��n�,��Z����N�J���KGve. U��T����a6���������'��o���n7}���ʨg��=�@)#7��9{+��"�m���0h"~nw�s�ywI��T��%C����Z����#;2U�����,hr��J��r����]n�p��iͧ �:Rh�r����j���IGa�/b!�o3�n�,�m�ݖ.h"�"���uH�6�#F�ɰ��tT��.���^br�W-+���8���cbKl��.��9� \��w�u��P.��H���F���IwF�q��_��kx���*$yKi�����mA0߸re���m�m~v�=s(A�sj���iX���i�9�hr�HNvݧ�&��3�K&@t�2���Д��5���2[�wr�J�]�>��+�9]f�UUT*��2�C[ϡ}S���&G`R���R����_��*�O���/�eCx��aO4d �)�	�%.Q���okD��"�T�]�|�bإ_v��sJ�<.ˎ�/�C�a]o�Ů�#�@[�G���c��b���t1�VsfJ��L�1,w��YmXTk�n��!;Ndw�H0�˃�1�3Xi�HU{�5�a���`��<�_���P��jygF��
�f�;��Yn1b���_�SK����A�&��9m�Yn���.#:��/�ov�CJz�e��W��:�ĝ�)��a����F��a��9 �z�.Ote��e�!���'��;u���&���okR��6;�*,P( H �jA�n�E'��>��MQ�R>6�E�].K|,z��k�LFKMs�{x�ѵZOx���ԯ�Zd�HuϺ�G��~��C�������::�q��}�?�슉���,u�;$���k������s�a9������9��{��4ˢǭW3\��U^�x� !T�;�E��� .̗�����gW��r� FW�(��n���۹Q�1���RE�B���n'��."嫉�xGW��`.-���B¥��?�ÿ�U�I
�7�[<b1�hf��D�}pN�2??=-?�^�tdk�B-�E.�t��J�l�
��Y��<��!�����Y�6�h�?	���Tn@�t�V2�g2�#����h�ʌ��3m�G�����t�T\p��s�э˱vx��p�dI�7�)F;�Ke�7��U\$(��	bYla������$X�_���{�8"jƐc%��� ���g�� ��?V��d,+�i�!ن.�(u�#���
�����p���I�l^��w0��|�-\O�I&����4	��s��Mi��9�є=�3�?w?`L�	#��m JAK�}D����i+#v����h�ؿ����r�Ce�Z;��^�N��������!E����Z� �?��DU��W$�,Pᡖc8���h�رX��.&e8*�A������;M���L��	��̷�I�Ƀ^�p�;�����̹pUB%�?�m�ڛ�,�B˶�aaBp.�+{Ph��C���v3(Z>n[\���3P-8�,���6�ޥ�MxS�n��T��Tq>x��d������l$w;XX��e�%��qq7c��&��$���{���G�ퟔV���/��`���~��)[y���J�3�-�<�Uf'��ҭ+�l��7+���aZh�NS��is�H�/�E�P��g��q�� ��N-�����G4�Y޹��]|�`�!n���
Ǻݫ��6�͛J-_�l)��{cA��X�댉A\�`�����ÌNJj�{%}��$"����&RE�&�,հ�{�]�14X�wI���j�8��~��j̭q|�O����vm���M������7��D����-8�����7�l_]g���/;x�{B���B�0�=/3�(���'�N\�(�!C�uy�7��U��0`���f��V��qI�
�(�������b\��ֈ��<�;KAD�zS��.`�hCѲo�!-���D��9��ۃ�l��2`�&Zڼ�w�-����=�����L�7ֆ�
��!��T�l��YK$鑴3�?�|�_�O�P�ԏXG�K2g>�]��,Fr.Ŗ岃�mu�кB��]���ی��Հ�, br�}W�B��9����X�Ri)�+���d�d�c*L��A<JG�oq�ۺ�U'o?G6��BA�ׇ�B�������1}������&w�f�~���`ږ���a9��6�@9�?���Y@f�o��HڴL�n�s>+3]7Gݣ���~��Ò�L`p�T�`hS{ۑP��� �z�a�Ky�,�C��lm'j-0r�Ҁo������y�+F�@��ڥp{���N��7�����B����o��6I�o����G��g[�ĥQ��Y��pU�p�)z9���3[��4�K�KZ��4���L�h��6�{t��|[s�a=Hq�!ó,mKȲ��\�Nb�$
�'��uX��8��e��U7�(4�w�����f�@�}%Pͨ�ɛ
�]����$��RUt�_^؄'���m��2p�_Ax������+~gT �#��u��q��8����f�&�KE@�D���f�E�����������u-�*��������U7���0�����Z���`2�h&��T
���^�p77� )�/����VŎX���f`6�C�Q�T�mZ� Ns�Z����p����P�Y��������Խ�M}�G��!��w���Xb
D��O��n�U��|	���mU��a
t��ͤ5�߽�.�()���fY��H����&k���$|�jϿ|��H-�#�P��4M�$��� n�a0-��KP�G�H���-9���	���+�Ly*=KLWAP�sG�w;����7�\�~wbo��#u �� � �D�����b�Ƞ^�-�:�7�@��5ϖ�Z3� K�]ppq.(�>H~[��Ea�+�a��lˡƑ�[>��,����pwJ�/���z�p�#��l�a��nG�U�"o�
�I/���_���T�p�1�/��/1��#�F	�%e�1�&���fOח��������pG�G8���o}`�����I��þ�r$?�� ՙ��������7�
�y���+^&@��.=;���-1�O����AŸ�ȷ��⃂ }W���d��ɁA�{���S�|������@�ļ�\�a�6Ѕ��`��Dr4��έ�M��*�0�����f��p���do�e�飖�${غ�|'��@ܗ�U��8(Y�$X��c<Q�Wǈqa4�iҠ�..���p����1L����i���k~T���+���e�+�	8~�凁0��coXSZ�� �5"�����B��/w�~��r��.I��ok&k�Ŀ�j6�����T��.��$F�.�	 =�g�҄WH�J!�+bB%�#ar���])Kp�vZ����Tl�ְ�L�n(�Nt�ؔT&��>3���sw�0���jD#�Pk׵��I�|G�5J9�=�P���5��:�}7����^��u����2�L�����h�_e�+�\��h͇�{#�`��$|���y�S�Y�#�+�J���8N��P�]F�6�RzDv�՗L�N�s��GU�5���@�ߕ�t��ɸ�8�=�UV��J���A��d�5�A�ڈ���O�]2�x�@���:�)�3���vW�S�]M��tJ�
�T<�Vr�� � %�I��Hɂ���K�'B`�EO�ʵ�N|�yV��F>��)gp�#]"��s�����E�Rx�U_R����g���Ф����֬c1�L:?�8@/�a��sȼs�\�jA,(��)j`���쌀���@d�����#���D�����[���u�6��hA%\Ld4�d8� *���0S�3��g1�D=��l@��w�C�p�f�@ʶ�+.��_R��P���'��Fo��"�TI7I��<��ZXyg��Ř~�]<Ҟ�̒��w��HI>%�}��v��E�]ci΁����'eC���[B�3d[lz�l[0n�I�5��]�1{����)L�NG��v`�S���gV��\�U�����$xd����_�n�:��y�$�e��e����Ԅ�kl�Mݫ�-qdl�J�B��q��aS/K5{���J%���ۡ|�#�i
�7�>;��M����P��4Fh�j��_�G6��V>IԖpMH�D[�_@w�!�Ә��ȹ�����p�	�����M���HJq�*�M�Q�8�3����тg�d&���%?Y���JR�O��d�Ζ�xT��8�%X�,�X����{TJK�5V��_�v�yT��2t��w0��1����(l;Z�bz�v�ߩ�G�n��Jt�CP�6�|��]̩ ��@�h'��<���r����ƅ���h�b
�scc������9��!&�=Կ����m�s�� ����;�߼�����RcZ(���F��b�7�=���`���?6��C�م�#"f�?���SK��%�j6�o7��J΄�l�/u�_t�B��1�O�����j���$uP�U�	������+͙w�n�`�4x���{���ToN�����0 墓�⊗�ERKٷ2���l�h?�`��r����}\[�d��+eV^	+�	QVR�Ї`gw(z�ִ*����
F}�a3��c� c��N7�4a���A��u_X�����jt��-�6ݩmI,��}-�?�m�k�
o"=t�/��Xp�/��c�S�!�������&�!?:�l>��k�����&����C�0����:ϐu/�xTUUF���5�	ĩu+�6ic�nG�ˌ[�;��_+� =�/��"�Vr"_��+�H��-�򗐟T4`�����Hۺ�(U4�CKd���c�0>�q�`�ď�n�V�[�z��\�x�TJ��Xt�|��9L��AɣdK#V?����04`�3wwz�/r�Mt��0�ӝ"qe�d������pH��W+d'V�W�I�B�M����2�ֱ� �L�7��U���!1��O��Oo&P�QL��Xh�3]��0���u�q�Hv;�d�_��6/�zt�����g���\���6�b�����q�7r���L#�W/�8��U�J'�9�rFDъt�Ǳ��$N�f۶���n����"�?�R�kFm�k�����C�W�u�e+u�5���F��u!B��U�
'x~�^��(y�w����Z��l�κ�-�T
�����p��
�ceA��.s��P80]��؀H��Z�HN�A�C�
����'=&lcUB��#���ֵ)} ��6��x��f:U%BLt�����,��h�-uk᦬s��HOťz��
�r�<�m���TG�p	�Y�&i�&\6m�K�yz|-�}i��\c}�\�>�<����~a�J�t]�M6`qŉ����/X�����AM7�­��%ks�4��&��䷳e,F�L�>_�@� �Zt_�Y�]�l!��Jst��G�1x�tK��ʵ�#��� ���]#��J��O�p��㵴x�,�2�m����H��	]��j0y�DCKE�����i���!(
���i6j�*1-.�(fz�UW&�S�5�� �+#�~fb{<l���\m/��<@��)'ӏ�U��l��[�������3�@�p�vdHf �>ِ��p�'�4����#�!��hP��n�����/����J8��y� AE��skR��M��[�q��HĠʾt��'� |Z�H6����f5�5�5]��C���ÃE��5��$�/m��U�y/~X�e���=7K�.��s)R���U�d1[��e�S�(����a������3�0�â� ���;&$Y_'ݡ+C`|�xź�3���P��#��$�Ǻ��Q+�@1�}��(z_/�%s���)�ik�.�ys�MTe��o�ƍ��>�
)�4r��Z�}�7D/��`q��~��gм�����}��������Y��*�[>~�f�w2��SO���Ei��qXޫ��������c�ON��Vn�N��=`��] ,��=3�"pc̙I��|����(�jܐ��x�����R����;.ns��yd�Ȃ^��U���w��A>�|��ȡ�r�cf�1>ͫ���_ҟ���s�~E�w-U=]rF�be<�8հ⇬r'4)*��R#�*e��	���B�){d��*J���RO� r]j�
!U+g� �<'�c�|U�H�Is�X(i ~�Y[�9Y*����{ 	��cA���A�<��.d��!#_�� �(*�����5���ƃ���ʳ�E�"^[�~� �ȉ���0�o&�8�؍⟌��l�� �(^��z�G2
�/��r®�J���j�V��m-O� <ل�ז2�������|�a%-���/Ɗr>�.^ᨒȤ���*`�_J1�+O:��rQq7Ee�ֳs}tu1�]���l�z�c��y0�%ӌ�X�D�A���Oz��h�=+o�J���w�m���޴��Y9�R�΋4�Q��in�[/�l�� q�kp2`f���$&]�^���K<Ⱦ��T�w^�DzD�W���'�F���"�����=��%E߀�6׀5��N�;d�o2w4�yX�*3�b1�2˹,�~~�8�w��WR?� f���a�Y�Ӓ�z��_����S}�9n-�:� �FG !�o�`if�U��_�ȣ����bU���k8�pMi:�2ꍻ�b��u�V	�e{�(��Kp�/�p͐���j=�GO(�6�o���(-b��`��B@���gS2[���d	y	XЀt���V]8���T��G��g���q�S�&�`:ݧ	{�E���}�� lp[�&+��f���?Gk�2Z��2Í�S�IP��������؇��1�\}=�,9���%��M�����7�7�Y��D�6{���J"�q=���D�����ڢ�>	D��ɚ].!Y���ALxr����F���w�C��\k��4� b������X%�m� o=Xa)⬛���1"�&�� �T�8O�����3�E%�[�{�{���YR%x�;0�H��0��4��4C�'�@�
8�9�o��?�9tb�^�,:���Z��Z/��÷-�k;�-��i[�T)pp_7]�	9L�q$�d�f������b�:nl�G���lS��� m���c������������Y���Z����NF�5����	��&-�9�	�����k&� �Vɨa���'<��ЁI�?���(�5�::[✒��9^zpu�bK��y��j6]�*4����L�ա�\��j!qR�0��. E�/Wm%��]d�(�����#��u��B�I��M�"q�s=�{�y�������;S2W�aP��꒲�
�Qz���lOw�U��W���7h�p]2@��g�ڜ�7@qL� i*�k`��>�֭diK��+��_�ץ��QpJ��R)N�GY�Txy�R��U�5�9\ls&���T��O�]^_\!��Jaxz��؂6�d��	�R\[eQ�B�1c��|�.�-�1t�����BXY��İ�}�餹,4�UD#��P�=kJ�2��ހ	`�ǵ�)��iU0�7eg�N�&�Tc�J{���"-(}�	+zd!m�%�Y/��2�Y�\�)����?�>c��:��J/���p���9��P]��0o��F�Ӫ�<^hb�o�q��|��	�X��^ꅬ���W�2�A��0^o.@~��e	��p��A�zQq��5��9뮂�Aj����W#�7h�+5�V-n��N
c�����
R�'��غtA�� ��4��a5dU�k���n���i��*��ۜ���f� '�#�AU�P N"�����%3vQ��b�J83IjU�_��w�0?�UDMnk�u"c��km=/0S����t#�yD ?k�C����^s�\h����?8e@�����C,x�+N����T%�o�����z�k��r;d��l�� :|?֜�-a'|��Q9��+���y y9�~���1���g�H���e(�fYd���vzl�
<N[�?�^g���|i���3��3пѧ=E]��{o.y�[����q�ě�h�ڽ)�g_�c�X��w��ݶqbH���@R*�Md��)gh���w����K��a�/Za�D��I�l=���o�h�FMy�����6kK���(��b�6��������)�ֵ�g����0ݍ
K@�@���I�x�i+_����[0�; ���t�+�x�������a��A�Ȗ<B&m֥xaL�5��fV��3�P���N�)Ra!��k�Ǎeh���r7�e�G��mO����@v�]Y��ܟf;���⬏f��@z���c՛*:��̑���m2�&�<FÑ2�dz��/�^���s�N�Ӱ ���Lla����-���bh�6�
%�}JiP)g���F�N�)܈1�C���S~Yj����-��y^���W��Uw�-jq�:P˪_8_ޥ����ϵ��r���J��x�$��0� ��tC@�6Ǧ4��;p��{Ӓt���0Z?��1��t�	���{{�l����~G�]*2G�r^���1+��ky�R-����I �^������G��G	�༒����&�f����گ	�
o��x��\��+�/144�c"Y.��?B�'���%�X	#�2x�}�����$*PY;6vۭ�N�R��Ѝή!)��
�/��3"~a@~�l{�X9B��t)�7~k�.f&p}�	r��y�FR�)U�z���L�b���&�nz�0�Ơ�ȠAq[�~�p$r�w<9K�dSw4eD�qdn��^�42���q�8�a���Z:�z� e�yK�I<�
��׶ID�tf���V-�:��� �lI��e|E�LJa)�9oL��c��1�]����4�)M,ҡ�����9�{s��PB/�n��m=�7�|��g/�M`���L�T�?)d8`ۇ����(�;I���֚`jg����{GF�H 5�~f����=��p� ��z�s��a���폈��fɟ��O�;U�u\'=4(�z\��#�<O���Fl]����f��<y]�������"H5���_�,���ڏ9�x����7�rxDO���"��>���P���\_5I?����5 ?�F{V#� 1��Zb�Ʋ�B�� T���S��JH��}�u�5���фu�'P23$��v��Åz�3
�|%�����9���E�@D���3S�����f%ms�od�s�ܫa�+�Cp8�+���,V����3�!v����&+]�'�檻c��@�`�6��?ӆ&|�tς��[�5j0��2�Z��	0�&u�.|3��5��@�Dp.��p�%�[���������:�҇�g�گ`s77�8�'z?)5�B���@��	� ��g�Ʌ�������"Ͼ�أ��_�\c3�=ߪI�m����<���о$]�+�����T0tG`bTnL"X|V�7�䶰�]o/��t�~�dX�w��u�E��Zѕ�p��we�q4<m]������d�����Z�?��'C�f(�;l<c����a�r��"7>�T�,X(A�i���S��'x}JqRQR	8��Fl��I�m��ׯ�5��}��vi�o��u�٘�1��v�V6������1�@��Pi���"Um�\n<L�/��
`n/ޒ!bW�E��5���H�����(�:.����P+�-Q�7D��$q<�uS�JެB9�w�^�;���#j^��Y3��� �6�C��9~b��[+�絥k[��)Ʃ��1XG� Sb�ñ��5n{Y�(��ܮ2�������|b<�ucz@Z�\�Bo��Z��/*R����� E��!T�	���Qq�����F[_�:�|�k�'!���T�oB�dh��V(�D��[P���6UgM��q�;Yѽ�nZ�x�*F�1�s1��G�k��������ٌ�#6��|�<U�[����4X����OD�Т�u2�[ɿ���c��v����;��'�2���5x�ͭ�9��Eg�D̺����|xgAH����O	睫����b�:u�.�>��3���@���3Ґ�=��2y���yjDl�YX�>9�xqh��CRDX`���Gd�gd���&��يϮ�E.�|�=�#C�
V�=���pO�*��'��b�IsNƋ�z�E/Q��zt1�r�꺋�>/�����Q�AC���Ǆ��no�2�%�dn���í�Y����b�Į�	f�:����m.Q�2C�I��)�\n�囶��z�� ��Pt+�D[�x�.�hR���*W�jFa���Z��;�9���o��b������uU_,��� ��M�2�|`����:�(� �S%�$v�T8�hY���6+�4��<b~&s��UL�'� V14+r���W��-��lw� L�D���N}d3z1@�aCl�ѐx^�>�M�3 q��`mdmݟ����l����������2��t�4�-��ew��ڼ�"��
VO(�7�����+�r� :��1M�BE2^���"����)���o���5���F�����k�">aP8-[C�S����q@B�ʟ��9�e�#��@I���P�d�+���t%(����Z'f�~ x��$��,:0���w�u�;1vtn�w@P1U��=� �w�2��P髩=���AB���?�n7�V}ٮ� G�Γ�('�79b����+�L�:�ª$�u#�)��b^��G��K�	�TyD>���`Z���ɄS����-���8��ݐ�E����N�b _&; u���)R̷�*$�����k��������y�<=�8o�&��E�V�l���=><r�%�N[�O��r��F��N<?T�-�ɶ�6��!%�B��: mƩZ��w�Б�&3�:��7�΂���/%���Ԣu��b{������&R�9��;�=��́���
Z��-�+^��j�H��%� ^���`:����2yv~Z��A(�QyR
����l�J(~��F�ЎA�W4o����\��o1�9��{`Q	���fۺ� 9S�Wҿv�j0�d*/���r�w��Q�O_���=
��ws���!�=��.HE���
@hw��!�,�����,ȟ⎉칅 ۦ����@K)��P��˃$B�?9�҇\SO�Nݒ(����M�2���G��_)>��U�!ёO��$�����gtq�ֿ7�n2�oi�؞��3���&�g�t��˱�Z�m�����;��aWCw#���#�	�UX�̃v�tSIf���;��š]Q���v@�ؓC�Á[� �1]����I2m�E�!aA��������_D}�rA������pQx�QEQY��K�|tcj�ǞZs�����&M8�$8xD[=Y�N=9�th��p��X�,�41��V�N&��x&2��?��D����l`��*_��Vڍ/J��BwƯu�J#���I�s
��l�7{���^I��]�q���O�����3���Nm�d:Ӱ���&�ٹ����t����X_'q�"�~�s��h/�
�=|��ER����?�E�;U�
Q���.�A��=�#�ɐD(�;:c�ra�ԃ����#����t8%��i~>�#Q:���pŰdr[��2zL+�-e��|0K'�>��C���gC� ;��4c4&&�|I����R�N�X�X��/�%�6�m]*a����?nx���+l�b��5m���I�LΆm��vBq��6rʦ�ڌ�x�c�qQ�K�N򀐍�6D�=.�?r���l0�x �S$����:�zU�,/�㺛䨁�$���tE-D�b�5����e�<|��S�^ ӵ�}�l�j�]P\ǧie�w���}�:�0=��}J9Y�g5�K��D�J���-�:���r��u���|�待⯮g��E]�xw��-/^�2��H��uT [z��p����-?A�\K���<乕���Č�,+��R�k��K5G����e,G�`JM�N��In7z��}d9:��K�B\���.����,:�+���]�fn"h��hh?u��H?�ݿQ�����oL���ح���1M�����O-y���I��(�ai�5Y�=Yd��W%���SH��ĶSWD~P�Z����]e��T�)��|d���ت9%�"�>������HlF�B�q^h%�6��<�#9ُ�$K�W�]�3%)�/\p��p�}����_yn�
��gV��-VW�Y�`@λ�<���9��×q�8�)�>!j SU1~Z�q�RA��_�3��J�Scgՠ����J�y�P�6
>3������f�	��e���:6���� ��kg��T�)?L�Ԑ �&�H:9��_y!�-v�]9b3q�=�4��j��т{<�����'��a��^ ���Td��0�|u��0>�r�7W;�zo�hB��M���ߛ�O��E-^����'>W���XR~ aJ��f���_��b��u-� 1G��SΪA��&wݻ��ȋ,C�c��}��	O�iS�*��s��`(M�Q�ʍM�h��`��mg�~ �e\Ϧ���{��>
���B�a+��$:�0�jM�����-0',-F��t�S���'��Tv.N�~,a|a�������;*����!�R�͏����a�'p�:j�H95>Mp�O�M��~�e�Ls�t]�b\b�7x�4�x�W�`?���{�J���Fm����@ԥ]\j��a@@�$��a��_(�T����Ȱ'#�@��:�P����-v�X�n�II�~�M��>����"+��1�tXU��E鮍�!O������2�l���zq8�fRO�a�~V�ʄ���|��x�����ȃl}3>&x�&�,��6L�K0j���˔=��}]q7k]:P�El��9�-�x/��9V��WM��;�(AN^cT�̟��2,���)h�>2�j;� �OY��B��s����RڽЗR!-
��v�᧤�P�ĽU!%�tP��{=�e�ܼӇ����8`��2�MAEj��ȷ:���*Ix�Ѳ9V���W�̲���hdE�{"�� k�-+��s\�O��s��i�7yr7E��du+��H,�9h�����uxxc����,�f��2#���G��)��� w��C��n���k˪�v��}j~��<�|�I=�%�yʼX܁0�+,�;��W��t��"�����c��Ž-C�AC�U�X�1��<2�v`�/��"�8!t�һ���R����� �b[خ�L���P�����FD嵀=QM',�ã0(��CDmX�_g��.t�",�<� �;L1i��]�V��Op��E�[єi�Ux;��;:�W�"�v�+H٥�J{�S��%��%vHA��C���x���,č ��}�:�\���u�:��4v�mQ����q SOtdd���g5Rt�H�o�d���0I� x�� ����D��]4c̗^�����@P�/���C��S�\��r6�\�g�Q;/Ҋ�H{cG;�6Yխ1ZM�w�W�A6;D�AveL|���hO!6P�\ÿ<?( n@R'/��%��	
�Mf��Hp�Z�G������bq��
7p�������㳷0%}T��B�����W�Q�#����^���_�f�������u�*ҷI(GqQX��$�^�W�I�����J�L��,V����	c/��<� M�ǖ�p
;?k"�r^���^��{��V\rM#���Ԫ",�j�qX��a'��d]~�)4��P2��w��'=r���"�v��44�����{-�װ/3"k�P04�'pW�b>��R�ۑ���6ߙ)�ڝ_�	;��Ꝗx�}�'�26(ϥ���2�	�O}MA��l��O� �p�+)��Gt�#F�T�*C�*^�Iث�^iN�����|��
��JU���].���GH�s�UV`����z��q;�8�y?���j��&ɜ��Rpg6��v-��M��8Vz>A�[hr�n�=���Q�l`����|�̴�i��dVm���HL�HL[.p��#ϯko�#���*��dN�3�M�]�$�JnP"�z5��0o�z��܄$aޥ��-�E�+�� ӋU�^R��P���� ]6���.J�X� k��z<s��3 ޹�Ho���H/�*e�b^Ѵ.5��	�+(��H���KXC�˅<�C�^�۽4{ �K ��T>d�zrr��r'�D9�y_&��Q���ŘX+��8L��lCU�B���nmWt�~<���@�+�p��kw#Iw/��Lj��}�vW�I&O��v$�cj�O|����T�M���K;$��O�^��v�ݷ"{ݲ�87���5[n��/y|�:C���K�~?���K����^E聚�Y ϴ���X�ߵ7c���m8R e��\uu��'���Ȋt^���!��b���Y�\a�E���X�7�\G�q�����otP��/����	��k�Z�~Mb�Rr$�s�q�).3���zd8��9kխ���FZ������7^iW�K��1CE��7�k"vo�!'N/�����ஞ#���&R+�cw�sY���Ɨ�]�I�`Em2ߍ��Ĥ8�3�!��x؅#��dѴ�U�ktU�i1����@)�k�?N���<ǘ�`����tkט�IO�K����֨�E�o��*�ꑇ��vb�_�[��t�޼���)T�J���s�U���}�ۈ�]u*wO�V(����������m��uⅯPN[�Ŗ�/{��<,��F�̉j��-�U,�
�b��d�]����B��*��c7�0yo�ʚ�8��A�N�[C����j-%\kd p�����}�,��҈�u�Ii��h[�K�[x&�)�����'"����d_ȣ���^H"NFL�a�^8���xI�D�!��z��Cۦ��R����ޱE�
�yD����6�*�fc8kpwQe�g�N���t�#�&�*�\m�H3���=���81ǡ����1	���ki�t��"�����]�TC���ɦ�{Wy`�����}�*%e���ѱ[/y��8;1����g�Mz
�1R� ;`�ɭ�`ȳK���*\�s͸<S��H�c�;����v�pjN��rW+���YD'�A%���ě�0��k�;p��a�Zy�������?�_��6_a+�����an�O=SY�]�Dw���m�^򖵮�+���4B:�V �cdɲ��*���n�OjtK���d��b���w@s�p|4D�LT��>�ɕ�"���3]�p_��>늰;kS\hͺ���.�Q�D{���y�$YU�����_+ϭF�,bT�A��si>n[�e;�(�Z���~Az��:M|�q�{sSm��Ë�4sq��ԩ�����pMM��Pz攧C��"�iG�{8�����ɚ�חb˥���r���b=��p�Y4���oJ_��$�P�nʪ��P`uAJB+ީ�O� �(�ܰ����ɫD����.��W�I�j��7���`�	n)�}ᕼ�Jԁ3]A���{�(U�VU!ꠜPLX�Rl�O�uQ����5�J���O�B�o�@���&$\	����5��/�;5߉<[� K�a[�������qX긦�P��Q�C�á��x^1\��������'eAw�q��(m�_m�o���,s|e�����4=�/hLQ��,Οy��Z�g�f��6�aq&30ؼG:�:��U���L
P���d�2�C�!�v�D��|��gH�g�	���&r��
go���%��/��_��m������b@ن�E��"��?Q��_��+�A�
�h�	RʀvPI�
�n�sSsކb3�d�Β���%H�"�Ѳv�M� !�j=�I(:`-��
�5��!�p">�mS�`^+��T�I�xf�L/��|�Ȋ�9Kb�D�(_M�_�#0��$8���hQ����h�K�z1�O��!ac0qu��Ex���b�br����/s�j���ZFɆ,������k��X�Qk�
�0i��Ƈ	Ɉ_�N�$e��Nf�`�B�A+v��K�o�k��������Z��Y��z�'4%,�� ؆�L���W��z�ѽt5xUT��qW�J������l�t�����wX%�|�z�9��LK���>�i!mV��C��1�d�1�^T�m�q�����<�R7I��*�L�w�mxn7��y�\�s�Q���/�m�ڿ]�(^ӗ1�+"�A�q������y�x�V�}猖���q�]�%_9������4�j�c��ذR��L�I��f�-�͙��u��a��q�p½N����x�"t�c���=�>�%��p�e�9�:�v�>;�ӊ�����$
8���jy�u7hWQH݈��b9n��$�/z�	��aZ���>2SL�q��@��=?X��1MP؅,;��#i�N�y}q�i��0��������-���_i܍�/���Z��}x�g!=��W�zW�4�&A�B��f��A���=�dkR�j(c�N�$�o��E��)L	�ٞ,�ٴ
�tJJ�k5��4{�*�6�7㲆�{2ۉl>Q�Rz(��U2���o��|1�5̾<�>�V��Ď�^�Nm���ؤ�P���Ę���p_!�,(� �&f�������w꿈�Q�Ͼ�$�L�.U��7�j��I��[$|��D��8iF=e�4���6NV�qo�l-<+�d*���$IFg���L��XD���DHr����D�_�r�����qcAqS�d��+��]X{"�L)�Sp;żp~�g;n�-��Qh#8�t 	��~��y3�X`3��9y4�H����H1����R���P������ ��nI�@C�
K+M�%?�H>����!����_܌Պ�j�~yfU�[og��	
��K��Θ,�`��}=�{��y1"){���� �?�J(�������N�@��%�^�W������I����A^�74-��9H|6$sA:Q˛t[I�G��U�n-j�����e� Y@�1�V�Ax���&�a�7�M���#�pY�qX8X���&���t��:^��
�(e��ͰW7����&����p�U�z'��g3�� 7ihָ\'/���6����������H���g`�������4r�+�F2����22�$(��:�?O����}��֛M�
枣j6I��S��t�c�P�9��{���q"UQ\�&�ձ�e:>���3�",��L�b)_P�9/n��a[\o�\�� ����3�w��Q�_������L�BT�!G+�=C���hyA�&�g�)��\�~��\hL6�����d�����Gc3m���6LG�y�x��\���B����mfI�" ""�{����%��-��k��U�����[�,L�������/��,4�)�$��T`+�������'u3+��Ħ$��/�^@�����#���P|q��_ʇ�;�I�"Q��/�.�jj]ݰ�_
|k��2�%���#��-5�b`�f��cg5X�U�����
=H�^:�z���R�� �=k~�½��gz�rY��	ǵ�s,�KeW�^oKU�8�w]���.#�HJ��/$gR�!`wUn%&XW%�£
�=�;�'-}_c�y��5�/B��v4�]��.��J�P��sm�8Y�P5Ac��F�0����&b#���ݧ�JO*Q�L�ه�I���(�+�wN����q^���P��o�OD���|��|�_�b�d�7�"n�FH�y�*������xU��[��Nݒz���&��CΌ��x��L���L�������5��tlY2���� >vo��Rzr��/p"��8t��wۘ��D[OT��6�-jKp�%䖯Z��g�Z�$Z��u�
c��)�4�ׄcu����xbt,�=��c�	嫬g�)��|Q�,
6�ߕ�K5pM����;[�o���;��6j���=����Ĩ��U'�cp+�ھ��a�;�fH������`�.��3�R�D�#N���9w/MQO+�"�ذ��C�f�|��)��F��z"����Tm85���*�oel�p+ t3)��x�)��R��h���~����o������j����\Q��o�@����9�
�0�el�fT�<8�����? ��Rٰ�:^L�Kb#�U�~~��sp{��iMoӹ٬��F�%0�I^�?��݄��D��v���$��8�P��>�*�A����-M�,�,�g
��5�S��T���I[І�����ۦ��w�}6ď����~�H\i���+����}y�Q���-��[����)�9^
�.��A���@U'm�����Y$�찳*L���93��z!x~�#x���^Yz���ir�F	b}�ΰ٫[ϻ�胚�iP�Z?�+V�U�Q���a���Ƿ�Kqa`�*��앇zf8z��:��d��!m��_Qû?Ո�,�!p����v4����,�+��'����:�GA��٦�;����85�J��Wq3�p�%�_�X��.�z���͐Be�!��G��B�#J\�ɯ�.V�J��m�xW���QE�8؇=y����S;�i�w̄
A���@���v�T��MRL�y�gԴ�H���Jx�i=i�TwL�d�W��kΗ$T���nl۪d���i�d��������y�'�'��g�l��v�SIm���1S��Lo��^!Sȟ��aO��)}�I��n|��r8�� 3Oc�o%���Y��ڬI.v�N{QB�-�[�,�\���U�m4��f��>��X�-a㻓�@*�%Cw�g��P~/��/D���ff�X/���[�k��uhRJ�o4���1��3��� 0�ۜ�u')p�`3�3i5�~���H�����^қa�Iz��,Xc�{|��@R7Ĭ�`w�o�*��T�,:���xHh�W�p	O�w����2�0>�����0иe���v`���P�����eY}��sU��@=��O���uA{Z�)}؉�y��[�z2)7�Տ��[�����텚+�-F��ڻ�8]�p�$�e���2e
�ypf��@�5P	Ք����#:� ���r鷵�����d�wv1V�D�D� /!�	x��W��/g+����(�0��c�Iݞ��/�L�>i�M� �Jl�����!�=�r�H՘aPqzvT�l���P�9�KI��m��7K���0!��BF�ߨ�n�@��V؉�,w��mt����� #��T☼w��+ew��3��@��y-|6#�n�!��Ɗ��h!c����P��%�+��FT��~u��Q=���V�>���e����`f�ք"v�h3�NS�<Xf�������o%�a���h�e1Js%BT��vVǘ�p�`�>����������Nzuvs�.?�� ��_ �g�iZ[�'gC���y�L�L>v!��p�jj��H���ZB����%p]�O@m���q��mN�=�?��������: ~/��բX�(�UEh�3�˟	>�\w������z�΁θ[eǑ����H;���_�fzġD��Q��Vqi$�5��8XbR���/�[��r�Zk��v�H8�`����t����	g���+�sc5�慽��� ͼ��J"����UM�g�o~�0���1���$CQ���['�T��=�ݼ�o?��4 ���2���P3>�Zf�j׫IoB����!����%H���Q��XJXJ�%n+p�%�-�� �z}=4{n��o�**kG�:�s�!^��n�޿}jA��Y�������F�8�ۤ��t�>��;��O��U<�z�aM�;�$8e��+�צW)�c-�B�9MI)(
�K'��#���oI�,5x��g�%�;�zo�oI(9���g$4�r�|e]�$�N�fO��-1+Y��M:�����<��:�.�m�����A�;�`q��x�uk�|�����@�w��^�u-f޲�϶Knq[	�O���(iK�Bc�*��b�Q�}�rS�/�_�����f��8s[�T7�E?.�F�UFB0׆����)a�F�o�'��v��O+=d,���b �[��Q��[(���X���s���7>�5M���+��o��jN�;����0C�?aR���!{qF�F�n����R3%v��g9���k�����B�����&�b�rX/c��-�m�2�<\ �����������K/)^��}���'��r	�"ȵѺw��q�m%�0ˊ�j8 W�3<�"�aZ�3q�Jf~�)���д��Z��2Z��� ��Ux��A�c�����\{�L�TQx������F��tn�z���sU)��$�˳�ۄ}�2MA���ˣyL��F��
�]�KQ���*�h����p�'���9�(�!�m-p�=G`�u����0<7�+�v�qx/9
�?�s��ړ�������E���Z)Ŕ����޸���|��8%ؚ�>	�}c�A��A��a���i��-
�*(il�-qK��/I���o�0[�%l�����2Z; �{x���w�>}��;JD���|���a�
컣n�}�V��m%�j[3��1��&���ب%�c�b�p�zL��ƊE/���dY۷�F�I���R�Ğ�ު���k�$�ն�0����$pt�ic�"��;r�X���.8��L��?�*l��q�u�yg'&M�Z}����7��+��*����V*S1��4���_��gl�o��ܙ"�O��)�O����zyz����ҷ�)�|��D(15�k|K��llLڥX��=�t�؀��n��WX�}_P�T%i�iz��u�M�JIS� ����0a�<;���̞z���P!����% �����ΐʌ)�$s���
�?���Ԩ��2 	[�m���!��X�1�i/E��Q/=mGv�����3U�Vο:7zj9�E%����S��w�L��'G�}�:��cj�"ÒY��q9�K
�.jf�"���,->*�#������͙�۝�B���C���صN����h��d�+T���i����U7�';����_@c>���<��Ņq�+��(�{/;�$�`-�
�Ӕ�Åh
���#��|���[�v�D{	�9��������e��{�AJ�s���ԓ�#]f����Q�kYs�G�àД���p����%��y�ߚ��z�؍�n�_l���*�
��	�t��+3��������W�����'����д���
��駕���}���Nl~��,(@?NpΎ!��"غ��ū���̚�ٵ/O�A���#Q�H��M�9�ZLi%:3�_zR]x�g0G�uÖ��
��h���ф�3�O9C�w!�H/G�x֯}'��_�ǜ� �����m�pkR�����٤z��Q�$!��vn���p#�=,A=Û>�?~_�V�?�X�Gc%2s�x�R��H����$�6eS���ꗟF;�,{��x���2�,�H�kKT������)Ft�D}�i��+]�Ѹ�(:5[w��rQ0WQ�j�wI�u��`�h��s�C�H���R�E�@Dز)�j"q�C2�>��n�u��32�3T��2'� �S������4X�k�x���r���֖�qn���,�,�0���i7�`���#�L����׏D5�r����C�ij�<.��� �q� qWC�L����f�}XR�fl4Tp�^̖B}���rZ�|Kz5��K�~ǒ�vq~��J�Vi��_��#��~t\�M�eN�](0%�^(�>#���ܖ(N`��T,�(	���,�=v��Vd��g����������_�u��<�6�cuPPA��e��&3#}Y��c),Q��̆�d6�wy��	�tX�5%�n����{Ã��0U���m
��^�����D�=��s�$��/�Y�[�9��[x���`嫰k���#�[�w�K��W��-:S����������aat#6[gg�6|���4�65^�A����˧'�k�sEs�%>:�ߵ\����\�����I�i��I{�A�s�j��<�f�ۧ�.Ɠ`tb�l~n�f7�Y�[�t����W��'�4�:2B���G��8�.���!J��w�5�����O�1F���'�k'�֔e���8�f�,ZGt�ix��� ��i���s�,�@�7Q�)d	⺙���3��CR�l�ѐKY�.�mw�9�@
�E�b���(Nx+�~�W��b8��A�]*d���Xۛ@��S�ZdmB�l����둙�^754XW�2)�y�V�ܤ FA�I�A��ʕ�IA��d�׆u�\7�!���t�0�qI�LPAF�/�!J�D܊ߢ����h���_Gג��F0s?�N��'��7�lg�`����Svi gKY�F��&1pD��+��JD�|��4q�ʒ�>d	>:�s�z.�Ǐ*�/�jXs���ūS뭞Җ��F�I��PQ�k�T:	]�Ɯ�oN"�l>�OF�i�n��h~�Z�y ��4 x)���������P��7 �60Bh��@X%�ޛ�^Ec��TѴ�70xnG1{o/��$�-�W�m�,� u8z�_&���m"+�
�)��#E�-s�\��Ty��RJ�Eǲ�an9�(^��[f|?bS'����"�l�Z�zz3�g� *Į%�זNt�*=�q���>hQ��.+Ӎ�������Go�(��n�|�@�
L+��q��.�a��SE�8t�ۚF(5r6*	�a!5��{c����s�Lvbȷ��V��T(uue{�V;)l��w��)p��Z��)�ۮm�z�	������2D�����A^�٤ �6�L���K�	ɮݱ���6��yZ����:�M#X+����W.;Qb�v0֙�� ~�Є�"s�:���ı�����klb,X�4�w�^(=���d�9#H#١�����:x��0�����`J���K���4#}�����#>��I��jjs��� ��,Kf�f�aIA#�^�wH��?`~i�Á��I�d_��2�b&,D�ߛ�z~���H���C���y���"�2��]p��B�� �I2�l�ٸ�z�m�\�q�;},�U)zqG({�)����iVC�u�aK�%�������t:�>ԉ�q��i��1����I�:��ym�27#�w�%�<_��~��r�>5C��=���3�P�jJ�+a�tewa|���4(	��ۚS�}�sZx��{��C��.S>��2[�\�W$�`V�(J�����G��v�S'�v%���Y��sN�,��"�p���c�5 ����w5�� �r��4����˨�DPW�n@2��"R�=]3KE"���B�/�78/@���E�AZk6��]BLO���}f2pSL;��!1j���`7�*��{�&�@�oP�-����UL�fH��q��V����+���~)��|�ln_���D��>d������&��`��MÁ�٫�q��[ת0��}] ��)h�@�T���1�|�������uH���B|&x��V�T�݇M[Z��p"5��N��2ى�T$���~l��[w=~���,����Dq�L��Nw6N)�}#������<��i�қn)w4�X�{fk/��O���	h�^ʓzCz�ݒ�(i�&%��G�h�eٸutp�:�H(��S�l�/T~p0o�y$4���]�È����;L���Q�-��`^�:@�_�7l,t�|�v뗮�I��{�vȩ�s7�ϙ��j���;��Ï�+�LA�澳"� ��?����p;���Zȃ�(�i#��y����:����Z�@��X�~��66�%��<��-�F=x�iSY�1���ݖ�T荎3gU��y�,~�w}@�����cԂr@��P�ڼ ����s�gL�@Va�?�����(�x/���>.'��V�ȋW=�=n1����l�.;����QYy��������xp���j_�І�{����Q��!�`����{�o)�u+)f�͏��=+�ԙ��-p���Ӻ������.�-�؃�9=�i�:�?�.��h#�lQ���6���So��o��G��3�������\�s9�!'�6$�\>��:|�vB���Mku��b�:i�7ԦP&���	��E�ԗ��aS�����~Q��X�2F��:p\�g�.ۼ�&�����<�J��57,S@|m�Nz�^GR�M(��l���ɚ�'����LO���>E%�b!��\TOy����KQ� �d.��v˦�toOs�x&���i�������Cw�j�?�#C��5I`���;p�6M>1� i�6,�&m��p~k~�v����]t�mN���� 2�9��mX����g�`�FUN�OE�~��C�y4�X�(���|4��y̹����A��uֿˁ\cY�Ȭh��B��� ��<�H�%�Y�Bvm���&�l�:��`f#���ߣ��r�QT��$R-"���~v�Ϸ�P��r��Va�C���(��$L#���424�����7�v������P��c+WЖ	0���w�zp�
�*���@��)�B�H@ES�~���g,��\�~41g��W�da��+�K��R ���d ��9�yf�U�q�����j�� ����ʱpd�̅�-��c	z?g0�N�ꝩ*�`oc���(�^��~�J=��#B��m[��q��l�����p�
��:��gb�V�C�[9����Αh0�P/&�Գ�l�'^�<�@( f�p�P��-�WQl��*oP��x7%4��6�S��~�Xc
���C:v���"ߴ��>�vt:�?�塯"C��������:e8#�P�՚��)1�I��a��X�	¤0okQ��tM��k1�F&2��V��[K���th�Er ud˪�Z�c��%u/B�a�g�B�U������RIS>�e1�R�#˦��"�i��|z�D�?�.�ɞ�0H����-�F���{�s�[�+{���Y[�wz��,�qv����~���L?��F2��[�%J��!�A�7�{ھ���ŭ�0N�%��)'<���nщ�-#�8G�:Y��$w�w9��L�&~f3��'M��5c���N�7��%����I��B/��0t�5�*�`����[�':Y����T�Q�b���[�����yd�-L*C�%�"���X ��a�6s%��4����U�g��B��,F&̖���l�¼$�N�Tδ���2G֓o?>�+O� �Ъ��vIhc� �<
բ�)6ȗͽ�:R/��Y;]:7���g��$Z�-��(�5o6�r�@M�V#H�*|7�׹QaE�aq<B�;�2�8�(���ō�^Isn(r�O�J���