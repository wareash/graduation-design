��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� ��5���5o�h?\bv������Zr]�M�wM��a!��6���R�}���h���ƺ{K5I�*�q�p~"^g�3��j���;�ul��:m>s_`�i��wi��2������hL��ۭu�+U�u�.R��_�o���%�t�|�H-�*��I��x���yiI��`�iJk��B���e����O6��k��;�q_�׆�Y+�M���´}��E7!��J�Ż���p��_U띕Pݻ@�݅'"`&�1�`t�z��yE�W�z�Ͱ�NBi�YJ���VM���T�y�f�rf̟	�-M{�>!:D�N�9��!ċ��A(�j8����n[	��W�u#kNn�.0��$�Gݿ?&i�h����0�g�kq1�;���;���D�,]*Z���3�>YɬK��w�c�hx�]�B�d��ۈ�b���Y�C�.�e[�芬%!-�~�Xa7��ؤ=��7X���q���z�(��Q�P
�!_m
��"y�%��z���^�PS��N�T;������o�C$��No�qP75a�yHp.=su]�B^��9�u�oP���Y�VƎg�嬧���^ʑW+�C�BW�52K�?$#j�PXƝ�LGG�c�B�V�s��l�$J����*���1����h� J'HUg�|��P�������M�{@.YT�Jb�#�Bѓ�refU!�7��A!P-�O�Yx,5�u���N�Cي$#���v�հ��.A|:��Ec�-an����!������^�,3�"��ӳMp�T�֜K�� �#��/~�� �gvWRl�L�c��l�\Y�Z�'��R�"�>�<^���?�/3���c�_�]�EP#YDc����5@'�/��r-L�������^e��pH��G ���3vO�)��Mx�ܞT�z̀�#`�Ye}�8���c%�{����0]�������D�Mj�Z(j�- �5�)$&�<��yM��$#� ��	�؀����΂):���_z�pQ�.Ӆ���I�=&�_0EJ'���	.���q�U�s���='��@��Ђ�l)�&������Ua��8��x�j���e��L��A9�*����Y }���4k|>gd�܁��C��`d	���/}r��}�S!�R�d'E�v���N��m �(�������IG6��M�ݟ�!�r�"�u`f��w>- ������h.�t�^Ϲڜ
����1�� W����%�krC���W4N6�8�Т';~j1`V�l@�
�h�{�T���j@�m-���CP��gl�Jl�����o�(�ӃH�w��J���Bi�G�:5����f�y��A�1�@B��28���`�Gp�y������ `v��e��8�|C���j���Q����ll���.�<%���q�\y��ؗ�vJK����e;�È��1;&�7��]���~��������M�@�`X�x�R�`���<�e�'��u]ʌ�<�2? l��avGef�+h=�@
e��j��3�e"N�ϯ�ag꿾��+$��-�﫿���5�c~1�%K�Bj�d=�bn]�Bt� �SZ�jx�Q׻�欛(�)n�饔X�e���F�',,��$�E�@���&Q�����
t��¬N��ȁ�+�{�<�R5I�ՄX���A�[i�WbU��y� J�D�3y��m�pN� �پkm	��x�R>��Z���	��,�-EZ����n:��Գ�ް�@ <_�ԍMo ��p$V��!O6�*#��T�"��o~"�JO�\�\������M�� ���2_^Z����'|��Gdh���=TP�W%�Jo����F^��~��u����UЎ8e+;S;//�L�n� Q.�].Abrܸ�P���qwo�-���8r��хS�5�׬�඼��\g��+��A���(�8{�Q���5vX&4p�6t�7Mv6!��xm���^��u�,$�29�y����M�i��<%S�5MA�0�@�����j7�@nr��a�g�iQ�T5���{�(W���U-�c�>f��f�mVؼ����14�sjsv\�]f�H���ःc��$f��u��~�ǩ ��bF�`'3>c-�\֊(��祩|��	4�6�Nr�X��(+	V�^����2T�����[�,���#=f��C-׉���1 ���Ϩ:(�L������!)����2�"Us�G����L��_An����B��S�wST�3�#�AqnS�3-V����Z�~ˮH�ٌ�i�K��p�QuS���/7@Eb����4��^u��!T���=ɸ�#X��Q�����NK�y!�:�ƒ��nm��X�X���y�uJT~�6'�����Ez�3�{��`Ħ4A��i�k]��t����� 3���#�R'o��R	���ͥ,�8��]V*��X5��������Eƞ�@ �s�X_�p�b��\�8���L�f`3t�������욒�O�G��3f]۴�~�AN u�4�$.�c��[�K�k���!M_��aA���)c8��nH���G�[�VT�%�c��Ġי�ijW���~*��`�	�/��w������r��,��#Y��c��X�~��׸�|4-��
#xB�	� �XАN�;�3Q��sE���.�E`n��Yb!��&�:�<I���6"�6��I�3bK~k����X�����I���3N�ھ�=�4bl�f>��yvON�Pw���
,^9)r:���������H=�c~ȈL�3�}8M����xi��"f��,�)��M|�B��0�ف0�*2YY.A)t$�)�7gҽ��¨���uA.�Xd�Fm��gԾ:D����s���l�>�d=�t��o`$�F\�� _�{����ߘ�	�1�fESq�4�!��c�33�yY����2��^�d�7	d�h%�wwz� ����H����C<B��Ч�4����zZ�&]%�G���=�9��[ڣ'�-�@���b�鄡a�QT���3DY�+9�������8�۹�Iw�=(����3Ƿ{�F��S�=c|h�C$а����Z�Ug�)�hф6��8�:�ˉ?˔��ǈ޲�q`����R�x��.3����w�v�mЙ�a������^�d�$��`u���eW�l�a��q�U$�i�i�r췓8�!IS�kA���Ů��^��k��6]���\\��	�&�~h����l���7�a��I��Yз�Ͻ�����a��C'��ۭC@}r�qT�a$��{�E�pX՟�\ö�ɴmUϪ}}ŨA)����r�n�ARӽGZ5�)]��Gt�Z9N�����n���M��pk�$̺&)��G	60�n���G��9M��S�����!�F�@ ����Y�[b�颊�:P͚��d��Q�Ml��LG��s��]�&���*��r̀[�L�a .=_��8��D�ed�]�������Z�=L`M�=�ђ�~�Fs%��Ts�,:c��
0������/$�K�"s��~��p)YO(=��g?b�A{�9��îF����Oh�?�E'�����2�ԔAH����`��Hȣ��%s�r��j=m�K�X�����&�vm����ȡ�#Gɧ�Y�"�T2eP��5^�I�- �/�,b^}(���v-�g)A����9bwN�h2����E��-����6���K�R���q���?��fG����հ*�2C��z�
4��6�{Oh�u)�x�Y�1���M]E4,� �r-:D�軽tU�i����Iڦg��>?����T��8:��(�*���y���m��"���2`[��/(�4��t��G{�i0�$��`��}w6�|��6��>��勱�����YcF����]���G�5#^�k#��,��O6j��܅I��Un�V��""0�a�-������'����{I���[���5�Umo�l��߬�|+�}g'�S`�\A�<E�̥�SI�\�& �Ŏ�ϼu(6G�d�t���.��aZ��L���]��K:�Cc�$Dc�3��L��G�m��Jfe�87l	[�*�k*d5S����К�;�X�Z�|�	�et����'&�;j@�鬀 �!y��j�Aq7F7}���.��\��fN������·͋{ǹ�FR'D����ME�j��`1����'-��L��f��z���=Q���v^^X�;x�uQ���:}&�a�щ+T�����rB�o�&�	'��;@�y�KͲA��L���;�֚��p���	�P<D"�]�3!y�f�x�-JʒP�9��F\e=�`z󜞿�.tBY/j��I��r��
�Md�R�4t��I��Q|�;��@����Ŭ�[�$�N�S�!��f�� ��JX���~O�޶�u�;��I	��虩b.i���{��#LN+�{D��-�<.�Gņ���Ȧ��#;#�Svde��H'H��ۼŗ�Ve����t,�����𔁼�`�(8Z#�
R�rz�6x@꒕eCT���G��