��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|n�\&����'ե�':��g��7�SXk��Q\���#^���@ؒO�;��9�(���Ut!�\/=����o�/�S��Y�vT��N������Xv~:��Y:��O�*�<���%ǣ�	WWnn��+,<�iB�Bܮ��ҭ��F�v�w|
h�ە�����݊6"�
<����nڴ�[�l�&{ƥ�P�T^����� żri�Թ���h~�R��w� �x���';ly�(�c���ə`Cd���Q��RWƗ�Z��*n��|q#	�����He�l�<��zVgNmGLG��ַ���sx���~�o��]�T&��6L�;E�<���K%��Qc��c��H�RkJ�0�iY{(������z�,�&.L8�$?ԖF�\f5��Ө�Qva�?0�X4K2&�rZ~�%Z% �fCY�̨��,U�$q[D�Ht�H�|�mJL�d�-�K<��� .q��9��kj�օ�kĘ�����rYb�H�>�^8 �@Ul'�LQ��^L�g���8�B�k����\�ݫ�t]gG�e
پ��-�n�#8IT��u�^����W�[�@��a�L�������(47)B�8���;o�D��*�'n!�̵%�&�b�	���A���حG��̻�Ҝ/��_R�O�$��^Y� 0B+��ʺi�������-qw���>�T��Ձh�]��[��kp����@L@7򮒃H�8�xl:$�Y�ʂ3Y�uK������:�D��-wFq���%�+�t��l1Va�g6dS��	r9a�nNx��V��3�J �cYߵ���G��c��A�$�¬�&U�#j�Уa��ɠ]��}ܝ�g�#�:�g��l��,kQ��y�TcC��!r�P+�� �A"`˻���<R��b^E�]�h�Duō��W���K���^�N��a��W{��q��ǻ�����)ÿw>�}��g綐�P/�+3�����ЭG�$4�L�R�7�����qM�����Eua�Ano�������{A#�`F�W	��`0��T_���Q�$F������u�C��'^78���i��,�)�*��~r�r��Sɵz/f��߂���	�O�����>�R�����R䵉9�=���J�W�y�J�]o=tr��s���'cb�0��r�B'�^Լ��:l�Zx�@���{Zڎ��\�w&Π�������i�EO6�g-�I����i���X���_(��0l���s	`0~���E�&ת���Mwe���.O�RG
�[�,��V�<�XI�2���S�3T2�;��e#�Nk-�ˊ6���L�R~�&�+C+�`֨��f�-%�����H�_�BS'��%s�C\��GZ��m��M6�����K�oP8����z����O62������+WGx���*sފ�|`G�f3�o(����i-�r� Z�3T�-���
+-��xG{�Vթ`��%3�'��:���>�1{T�qL������l�������%^# ڍqB�J�i�MB��+"P�����;&;��LN�\�����^BYëԄ�Q�ͤ��n��)vfzFv�V5�\l]�> �Z��Ђ�D�1�0�<e�}����X R�~��ބ�����{8��0��+f����j�g@��wc�M=���G�`�4��c:DXPM�ʉ'�v��!��Pw �&�QB�َw�d뛩߯E'�Н�!@�~���#���kd�bos���:V��������z�*"�H���GFn�\�O��sF\��04�(z�5�0���&)�� _��`F��u�Y�8#��/g���z�u��ŋ�&fXp��o��:��-�9e�?�W��I��k�{��j����E���E�n�(C��B��1�Y!�<�N�57����(��O�0�i �~��4��x���E��+��$�Rݍ�|�N@C�g����k�I���=�&�+��J�{�P@��j-�C�n�Y�V(�a�7c���;���?|�8���H
̌3W:m%�vw�����it��	E��:T{:�� uX�dA�T�	�g~��͠H���C[�8�N�_�3��Q�����\{�?̯"`B{>���`8#n�-��v˼a��y�L�
�T
B��עV�YX|˒�4P�-!�)�:��ޣ]���aY�xPG�bi�;=k1<tZ�-��e>�u�
f�ք6�<_�����r�$f�!��昡��$���5(kRW3�eAG�h�R^����(κ��vS��+�b�!��y��dr]�]���
����e�^��Rq�8cn��$�������G|�Cѱ�"S�=�#�T��+/A�	!�~�$���YQz7�vR�j�!-v�I�.kn��Y>�^�Y@M��zs]�v9�Ρ���8+��+~Wا wm�<�ݜɸ�{��Ǿ��W�7��LDDbz+�7z����髃g/=�o`_=�G��H�@ȋ���H��z�:	��4	�t����q�f#�!��̏57�YH1��G;O�J5Oa�J���i��*���=�%�\M?#ײ����k�D�N��)=��`�K�/��������jf��4����]5x����V�c6�̏/�f��*6����Lp��"�*LV��c�(��������f����v�Ceɉ[.]z'�}�8_�E����8$R!�Z&-��9e�2	�7�0i�����4�� fb��A���� �R������S�R��8Ԡ�$w�On�i�S���S�}��O�����s���p�ڑu0?�S��L|��&ļ�@����]r�%2��FK��ɣV>TiF`��ʒde��=�-m���EN�%�c݃9ؼ���L/.�va!�ˠ��,K�vM7#h��� *b��J ��#��_�Ӻ£.п4�,(�=����զF�&
��ح�l�iT�y���`��	b��q»��nek�M���!�����^�	ޕ+y/E�
�8|�?'[�YfU�����k[���v��ɧf�\ͯ��2]f�yX�Ч��eB+����i}+x,�����nU��_�h�:��p�x��?�����Ѡ��*�o@y���W�zL���%PS�'��X�Z�-���e��+Ⱑ2��h_(v/O<�^���n��Q��ω ��ob�+T
�ݭ�	���ɏ"�Y�� E��&=t�MYD%�T�G�f����[��}���06;�rb>j����0�:#U�~լ�Lރ!2�rK���q�TB�O B]4av���cͤ����e�A֝Fܡ����_�	��,�	�������G��Ol�$t	� ĕk$w����|_��Ye�
���`���|���N��,0��B 7�3z�%@ͺoc�wJ7���bHϝ{K�5Σl�G��|!�$�͗��9������YR^G�l�$VW�,fL�^@u��FW/y<�$ޚ���dj�	���\`��W�*�BOܲ��}q`��iP�J%��?DGv/=�$�� !�i�NUH���_��* >��x�2�`��)�, ��{���������+��������g�%��v��m�0Z�f!���$OB�Ǻ��W:u���w�Yih�x�kWߊ=D��4������h�A��: ~
�H�˹hi�a �b̙s�c�p���ǥ�+/�.=X�.��`�ǧߒ{n�g_���߉�i��&j�Q��
�鲊a���z>%=,G�f���S�w΋'EV���w�&��g�~t�vW�:da�RG�)g�i��H�J�����K�AY3) ������}�vH06�d��r�n�_�7 
I����e�{gq�s��I㨛(�+�*���fN>X��,�Ic���V6�{����{����H�dfo��è��`;���,ÒXw`����d���>�ҹX�V@p�=qӄn]eՙ�&��T۾S�1����Rw�@���&%����7�鐮���ÁC�?.�t�'��y��C�,�a����w�Xw��
~��9T=@
Y��d�X������4�<��H9�83LXXnٳ�Hm��GL�U۾�y�')�rk�����7����Tܮ (@�� 5��ٿeN�U� ܗ���L��6�Y[��Ӻ�m	v~ᩭ�� ᇸ�M��5x��06gӆr�C��Rj�>��Te5���e���B�E��Wr�M��pv�Q�^�,�����J�/Y��G�3��xHgV��;�7@�h0��ͭ�Һy���ݮ�eD:Ne���ܲ��8���$4��ei���]���g<�Ġ$:S)�{�0�]8�o�$��#5�a7�?� ����	n��7�U��5�~�A�R�?�C�4G�Rժ��h��������B`E/-J���sA2|ׯ�A҅��F���H,�<�������?\���N�U��ct�&�C`&$��t*8������N�y!�	�§�;�	m������`;/5�[&�Lf3�?�w���̪�O���6ue�!�_��r���}����I8=/��?�f3Fr���)x�����Re�L�&�S���ގ��'�n�R��)�R^��)1O�-�TՖ��~��eKCQ(�����{	��[�1�����K^������c	������;�;�b�2Y��"�a���oM�Y�G;����{�PM*��I�s(4i8�	�w�>ڟ��MG@���@�����l�o=eK�uqq�	���{<�������z�=)��˦=1��MV�����}o� �j.䓷�<�v5s
Q�i�� ] E�(zA)��2V�j����b��R)-|���B:��|}��
gI�9����} B��<�]�e�6r.�n�I�-斸�߮,��a!��2O��kp`J�%;�%� ���H��#��X��,�!M�iP�xjƷ0b�cB_�H��aDDt~�$�n�����y�$�y�b�ne���� �Q`�*�U�knP��h��%�¶p�
������4�������o�*���p@*���1���u(���v2�|���iN?w<8��5�5�c9�%�wƋ̼c�m�P�@>>&�rN*2�!�3��i�F�0@��0�G�5K�y�ދ� �^��A�4�U=�d�,Б�$c������Z��W�ډ�Pةs ����Mۡ�Ts�2A{��t}�A&a��.���>D����$r'���2c�!��T/��l�Q�/��o4��˸���������H�nYM�¨�$�7?rQ��}*s�ۑ�1
�F83m�Gb'����8�HC�~�Ȯ�N�D�5e��dIؗ�.�({��_ĕ���_]GtӤc0t�-�/��ˑl�RЎѷ{qh�[S��G�@z�|��dcǵ7�gp�6Hb�׉��1c��Lq7���l
�9p��BVN��n���V�a����n�����9���|�z!��¸����c���DdCRL��+�\Qђ3��4q�C�K:��~�i �c��ʢ�O̯!��Zz ����ܼ�Ty��}���E1���Z�:ys8�5�n��	Uh�dR8��F��Q����e��<^���͕��j`y||`>\���t�԰���E�c65A�XԪ�*�}��-�0�{ҙb�?�t�B���\����q�d:�٦>C%D���\NF�)�B�T�����p �n�`�Ă�΃���lb���ߘ�HE'��:�˵T�7��B��ji,�)br�թ���%D��G-�/c����\��L��_OA1�p��z
���x�
 R�)�
�����l�$`��~�f�a|��m�x����HE�����s�XH��+;R�&�1'5��3�-\���"��LZ��A�3~Fy�M�٘��pm�^4;7ɤ�i=��� ��N"��B?L:s��H�����-P�� �; ~�+�<��6;�C����]������}*R�x�G��f����
�Vdw]��K�u��)�.H��l�F�^�&�)���ED��{=?F�@��Ú�35��-#ڛ���W^s
y@��9X��}��N�w7s*���D��P���Q`?�5ԷV���Y��R8L���lܤ�{��|B���M��u
9�m���_p�_�C�y��]	04G�����p��3��P���xE��`!D���LAE�WZr�Ӻ�u�vG����N��X���w��iQҒ�~����L�9W�0olz�.��%�ڮpVj[��˄�E{�3+_5 ���Rvb�Y���q$�
�gA�L ���Dg�%���� n;d��Hs��F�i��m;}V�3�ulf�I���x� ��<�0q4�s~�J��� ��-�Ax�����1�w*�gez��)�j�	[�]0��6�+^J5]�V��ԫ�S��� ]c.�K/{w���9���S;".5�z{>�"�~�9(���66nuN�A�����s�n�ѻ�Cr�y�9��G}��	8B E�{�Θ��o���8�x{@��ː����n��J��nL�?���ʌ��3D�W!14=���#�f:(�i���� ���m

 ,���י)oR��(B���a�B��g�ٟB?I#��'��5y��L�����7�����_B"���M���\M��3z<Sd���"X5����b���B%��S�K^+��$�$?�b.|8R��u�����̷��@c��S-�T����s�uI���s;X���k���(�a
��G�Gv�!��j�C{���������ڌ;�qԎ�M��/&���҆:^���G�y��f�3���
ֽ�z�wɳ冊㓤z��*��&��T�f?�ݭf;�|��k������))T���J����	D
�O�I몆-x�+�C��(V��x���3��+��S��ն��N%7����|75��_C����wR�q5.�#�>��E�2�r�����EL��?�%ڠ/\��(�b��֒�$�7+��[ڋ*j��O����v:)��ƤR�Ⅰ3�nޛ�t����t�}�HMw0�H� #"��F�����m��Gj��@�M�|���@�2Ge�>�Y=�r�����z ���VK(��:,�MA���$�
����DX�2��ؐz��*���q����K�Q�'�`N��P�%�g�ھ?�f}�n(��U�"�Q=)O�*�v��W�L�Q̄W���cʹ4#k`j�y�4t�6��Ho���vnb]!�$���e��dM^����	�Ջ�m	�P�v0�j���>�(
�߷)|홣�aB*�X�{[.�� 6��m�H�V����bk��?߷q� y����=�d����f�ؾH��`Î_М��UHfi;>��0�Pʂ�:
�����0��75~I�N��9�G镕��"XS诒R� �g���F%G0<�Ci�l��4r��9�/$I8X&,�I���w�G�?:�Y�p�N����YҺ�ȯ�?��2P�6A)���u���Ǝ�j�T<��~��CD):v?������f�74�t*y���9g��4o�M'��X�o(Ύ�F����L�#Σ��>7յ	�g�Y��쭒��Ѭ��e�5ӊ�#z�9c
*���a�6a랣9M`�d~Hu�c��N��#�D ��wuF *�P���0�S��<R��S/婷�bZ�_��2���ɠ�#X
�J�XWX7�L!�Y��u>��SOq��No\)}�N�eXd��{����~&oȴJ��w(2��S�89��fy6�`�U�������RijJ H���! ������ֿ�^�=z��Ŝ���.-��JR���5z�(d"�~] &o��H�A�].��L`�q���|��W�$g��>�&�=����+�A��|����+�h��1�2��pd�s?��*�Fg�Ї]�_�a���E���p� ]��H)�@�a�`߮v|˶�!��qÌ��Z`���\+y=�'Ln��ܓ�:o��u/ZA$¯��R�s�U
�{��Fb���2*z�	���Q��5���p�l%8Tޒk��>h�(��Q��dش(\ ��v�ѧ
���^��!���q�:G|<d�C�%��P�HoKA�΃إ��u�皎�n�K��h;~ޚ���P�\`��"'�G~.�	o��)��R���j�u"`(Y�CH���W�%��0��MI��iC�y���g^;%+W b�}{�j�'�o�%u����r�b�rb��,����RF(l	?x�jy,���V�҈�J�@C!�_	�n�&f���<1&�Q���G����Pr���JC���)�a�_��8�����%�[����4�m�-j4��eޑv_��)352H��}�� �8���Lꐽ�����*�l�:t(��s��?� `�I�? ��P!cI���l��J��U]�uJ���7g�]�qcE���T8G��0O7�ȱ�$H�+��_Y���Z�_���t"���M%/�I�0����ȇ,���2�TM"�2�}4#"b/���� �&6�Ï|������� A�L���VhW��br�]1� ��޵Hw��kW��B���
��]�������1#;`F�k�̇��I�?Ҟ���+/\­49������ׁr6�g"s%�F!�#�:͈���F�Y;ř�GZ��� �r���.X�b�����!���e#:y���{�
>�4�U���Ѩ���%�V6�?#
<2�~����A�; �I�|�\��x���Ai�����M���*y,�ܞ�/-"ߟ5����|:��/dL��gf0�� Ͱ�?>��q�{�sy;-��<D��*��F�|�0��5���p���;b4�U�T��0d�g��*_!w̴��0�V�N�Z!�M�@��A{�T ����g��GE+�ή�3�]�c�8��R�`�2�J;�?z�;�X�pG�O����Ƃʱ�槔����7��)!m&+�!&kD���ZӲa�{�cL��ۀ���זns�҂m�"�jsH��*�v��4�-���8��� ��`�-��+�����)���"�a������4��)��_S�����纯��&�8��}�K�x�74b<��Di�ϋ�����EK�~��V��nPƎ�A������G��UQ*��W(���r�M\jD���Q�n"B���Q@-/K֓�!�����*d���8�1$�'�q,�	��ͮ��X�^$�zPh��c0C�晡�qa;���v���2�a���=ύ�y%F�ӛ�_�Sb �d��j�Dj�|��2yO���*�>Nu��Y��������C��e���*�˯�,?K8t�����m��;<>�����#�N�z)V��u�,�n���9؇r�H�ߡ~��:��zW>�ݿ�'��Oُ��%���!�j�G'C�`��҆l��l���qI����ЋXS��bDW���ǹ�(�o��n���jW�Ƭ����@�,�	�IY�;z,���?�y�˳���"��B��0腹�#Z�p�@Ǜ,�;08��|��vο�'��ߝnOB{9ѽo��=��n� 
#���C��բ���&[3�R'�L��pZ;#�y���CYI�XB��Ba5��$ѫC2n��q;����lkm�,#���_���R�`�uqܣ��=������n��˔�V��A�}C)��;� �z/��4��l��	o&��r6�"7?鸻B��������!���4�K
a�V4c4.�+&�,Q8�z�2�TA+;O�˫-�5I@?�$Er����빩Y���#�=���M� ��^�G]�|�+D���t|���n_�����Z��1Z������˼�R��}���%��MW�_b )o(�~ �b��Y�s�~VZ���c,��r4Z��9"���蝙1��F���k1��piZ��x��q�ǝ����y=2�LW����,�<��_C��[y�{���!���S;�����၊+҅WhS���Go��;�x��YG�e�	q��s��|�
��h�$vyn��=[�� �x��E���� g���k!-�q�>p>P��b�+�#z��~ޙ[rlֺIn%�C�v,��d`�[INF5\��Ӵ�%�Eӄ��5�S.�*�V����������a�P)Y���r����Rݰ�����^��Q,�NwB���Y~٠C/�7Y�Ŷ�4>TF�fYjF�.gg�G������:�0�Oj8�L96����zV�K�We���W<��YOw�����5����#�'�A<����Dl��|�5f��-�
ʾ�>M�Q{�?C �G��q�� ��r�9�Ok�G	ѽ؁�:��(�h��!<�%�����K9N	z������]�����΀ RS��1%�:�@���XY��K����m#�=A���㤶Qa�J�&���6�*Z��0�/�k#����(KgkP�|�1^���;L����P=�hmxy;��H#�ǱdzYi�^z��Y�fᰃ��z��.��HxmXU�Ơ�q{k/[	a��ۆZ��ގ��۱�L��ᡳ�g��~����	��<�xHh?��X�r��ޯ!��f�N��*���u
����'���p̏�C�E�:E �0L{��TI�Q��akJK�i��SFro?|� ���S8I7���/�#rs���W��i�b��9Mm�ٞ0s����1F�ZD��jڑ:Ys�ӒV�h�9Q�pv[�
�-'5̻qJҨ/ܳ?�B�I�6J��B4o����;l�ZЄ]xwA�i�KL�&�Ϋ���k���U�<W"U��s.��{��i�L=ɓ�xΧb6/VИ�V��u�E�7rp��o0�~�bA�e���k>tV2�H�8xj�`]��X�;-����lo�KBkO[�{r���=�S�j�����?�����l�iMG�
�pR}�B���s�ѹ����W��VOv����w�7��-q�Zn��cv�n�1�1f�)���9�.Tc`�+�i�a���P��9�7f S�=GYu`?������k{�J��6�ы�k���	�~�:8�L���L]�3�0	t��E�t��P&)D=�w���[�����%,w=�����%>�m������h0B���3Qt���Z���9o6�������6�؎��M��s����uc�0\�ï�E.)A�ɹ���Yk!S���[ʜ�PsN��K�,9��m(��i1���p����h�t��y�^4��?��<��)qY A�_}�������{$�%�I�]U��3� Rr�=�_ȋ�|���wp��'�Kݳ?2�B�`�����풀��Vk��'+˙�bp�G �@RFV�w6f�GLp	�����a�x���y"8o�l��Y�^/� ��4%��7�hFʌEoEڎ�TE9��C(�C
�����Ԑ�<��2 �*�����H�J��)��O<�� �}4�J.4Hj�������Z��i�~�\�lJ>q�䤓'�}��k�U�9���'����u=��e�f�440ر�m��V�����3ʍ����H�O�7���[�������B��:��C�Z"���+�5*���{�IF_�����y�me��`/�J��lM���g��^��p��G?(ac�Q�3�����o�g�0g;�yJ*��̺�Us(�/�ܮ�V�>�^
߉Y���L��߸H�+�1�I���{9ܞH�ޕF���\fe���i����"�yr��6�����>p2\�܊7N<|�Nn| ��^�K]X���)tg�,��wӜ9���!W0��ޫ�����4�t7$4���t���i���3� �l��-	�9H���h":�A=*M�*��~��v�|vg��Lޮ�V��7X�{����_J��Is��B:�=#�iu���Dk���M�ԒS�Jæ���zer�%�|4Ԫg��� �J�IF��=kW�z鑯��p$��ٚ����(�*�20!"����,SÎK�.7-&���i�ݩ���8*/K����֤�K�QJ3�5:\��E�ѹv'��~^�כw�F�r��q��$��SSz����p�'��]<�rc�#Z��R?�^K���g6s��e"Ȁax�[j���Q����R.�B-�렺J�����o�����;��pl0 ��ȹ���E *��ॉn��Gх��P���(���H�D����`-�/"�:�&z1��sK�Q┛�8nK���)�^�|N��	�����Y�#�������jRSϒ���E�g�mR3�k�d�7���0�Z���$�~��^��u�|s�n�}���?�:�6�,�D�`R���63 �y.�2=B�=����-�֢2.P�����GZO/�T��ղZ����'!��>M.^R�o��Վ��-�v��Ϡ��g�Y� /7$�ud@���Q1ל�D�����l˞L˲W�@D��S2�"���~N�}Po����5E#����Ծg%S��2T�"R�tZL��z����Kdx��+$��a�MƗ�����Z:��q,� ��h��e
 )��<������C,ݫ��KϨ��#��L�d3����y���6�����������i�ʊAW��X�O��� C�a��& �k�곅�$]���T�U!����\WI����Խ^I�P6���{�t�FPo�{�ŵ��I���������tߞ�v��3s�9p��@Д��ԩ)p;��g�����u�]��H�/���`������*$�J��9h4wn	J�ŵB�	Nd�l{~�_g�;t�
�9��P(�G=�u���	��L��`!�B���!�� Om�꓎��_�o���5�Z�4=a�O�/�H?��9�[E�.�n&Tڏxz�	9Y�R�X�GH |��5Z��L�������_M����K�F���ڢ�9�����A����{˵L���jC κ�B>���Ry�u���V1�@��bAJ�ƥ�cd�1�D7�� {���9�vx�H��xV�=�����~�`)��
v�9	��G�*ݡ5%��_����{Mk= AkYC'��#���{=%Uf5"�:B�TI�KF�۠xvP�e�Z1]X�o�![�Ҧﻔzn3����,�A��ْ� �/d���y�غ�XbsǪ�+I��P������<��0��$��v��G��԰U���E��>*�j/��Y�zD2n2�sc����j�oe�!�	|��z,��pD�P�f[�:1c�Ľ{�+{���B�c?�8�z�p}���CR����g�o�ްxJ�±�f}a��`s4��	�4`������� XA��ƫ��I��M�6�&��(����>�:��n�f<�qH)�g�P�<N���wX��b�Wk�d��uǭ���e��{.��ywS�7H���DC���I�����hU3&}\I}�M-ٚ]V`��~oDc�F�+�&������K\�O^B��� �W�6?V��@��lA�yf��_e����P�w{ec� �q��s���ⱱO}s�qÃɹ�Z���T��fjRj��Ʈ�D�����ñ�Å�A{�O%k�(I�hS�4nz�)b>���m��:�����p  �T�D�pQ9ʼ�����h撀O�rzsID�����@PȏM�mv^H���%���~�����X�<*4���H�I�����d�mm�	�,Eo��r%s�y�{Fe#������� f��<��c�T"��Šy��u��˄�����fȂ/T�J�$��@���$B_���;��a�����T�^�l�mH�S]m��s��H��F6�m�4�F9񐢪eT*��+ba4~�u7�zZ�习C�`�)�O�\t�:�ā[�R��0O#��8�Ezq�)��uPn��]�*�	FZ��r�;w�W|&�-�kwc�ӗ��q����B�(��b8��O��rT�.��ܹDN������9Ξ�OΣ�/@g]Pj$+,���g��/��em1�w��!1�}c��!S0��`d~�`�&9��"�Z�!��L�Y�0'�6���QM��P�=Jx����U:G�Kj�Q�v_5́���Q���P��E��X�G�����)�G�}�q8��Ii�Ai��[	L�R/=#5A��յ_T|�S��B�Ԁ)����lYߵ%Z�Z
�Wuv}I����B� H�_�d�t/�	��oQd)V��8A�N�B�*��3[I*^��P��3ͬo�CM��M��zQ
�#m�ڟEɼP{�
�/9#/G�X�%���4'��rק�QKb��yf�r�>�Z�Tf ��I,�o�Mp���烱̮Q�ư�@��h��6�s&~mH�#�!��U�9*B��|8��W��x��Z�����M�g�
��eW
�40�w�k�/��ؒZ��Qne���`M.�SI�����S,�[�:=�{�U�狠(IX#AԙQ˵`X ��	���:�g�
Т��X?' Tw�J� ��̈����4`K<�w^qe��~�b�4�-�?SD�+ac����'�~*!9�	YuOz+��&�+)!F��I9f���X�&�k�v� E�7����ʂ�	����4m�''���$��?S�9R,���z���v)Z.}�e%f���K$���;�;���o!}c<�?Xڮ���,Qأ����̊��G��,3��R�1�$Ow��l����kG(v�|�o2@�E�;�q��!G�����6N�ED��<�@DP���K���w��HM�O�)����{����Y�s���s���/����d���o�+���t�.�a�P���e����V۽D�i�E�&tYy�Q����O�{i�S.�Βd1=���g��l)؊ueɭ�:愯�BVx��"93W������,���[���0���ϗ�+R��O�ǭ`%sЮhH2A��οw3��T��B����P��Д�_�Y�;L��A���,9
�s�� B����*cr��)������O�3;և�n�~�A;��U�{����,S��f���vy�	�No�|���v���CO�����M��� q À2�e���4/�ȶuǊ���h�r����|,c\Z,���v