��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e����d���f{��@����S��>���4{��ת�AO�Q{���~�}Q_�=�+TҒ��%�v����5V4� gz+���B&�އ��_� �k�-&�%#_GCz{*������m�h~�������9|��Gd[y[�dhsD���@q]G{�<��g}�?��[�i���U�f��!��D�qP�� u�5���Xvc���!�<�|�]�D����'�UY٩��(�HlVY���9�|����pm�D�*�qE�K'�zXv\:eX���][���/��~����F��E |�U��N��RQ.��e�c��_!�3<�zW�$hD���8c������to� o�D2�MAK�5�z*�,�zk�+�dzl�� ��?�E{n��Ib��d�B�:�֡��Hm�;��A�4EZ��}�s�g䌥eH^��|�T�U�rb������'	s���a����|
bWLEo?�g��yV+���"iM�Q�j�6Y�$�BG�LB�h���M�����I�VG��4�J����/���&�~^��g-�9�s%
R�CZ�z�S�t�!G�k�vs��Cr��9P��8�f^"n�#�s��	#���6���Sq�:��+�ӄktY�����$��3�U����akPL>��s��TZ�����;X2�0ż��3����x����ѱJ�DLBeo��1!�tܫS�c�ڤؗ��j�+�W$rG�yb"q�&;��!�������ݙ�/ȚrGaxAu/طZ��c�D�-^{m[����	�痶c����w�Uv�����ft���<����� �����B��c�\����dw�]��m� �c;�s>�1&Ε:X�~�k��K��h��:*����b�'%�g�Q~>�S�,6�����
/>@���
s��UV"����+Åw�4��ƶ	�qE?�0��w��Aݢ��}Z��4�ݒiL�����t�Zt����X�U��?�ɟ^��U�lPS0����Bv�DK�=^�$��X�}�X�Q�uy�b��H���̲��0Z�B5���!��9P���\��֪$��y����]���)���`��+�L�;�)&�8����|��ݠ�� ��[HbE�&���h#��|.D=?��f ���3��)t��+Ĵ4�nk�pa�өOɷ�L�LX=��T��4��c���q�;���9Ђ1�
���{�Ԑ�W�7#cx���Pu�ѱ<ܬZ����T xL4�wH���FI?�[ԯr��{J�;"H S�Z��U���y"�mX��	�t i��sv���v.�X��o� �p�49j�Æ���"H����-�qQEgW���a5~A_�����3�)�܆��9�g�A�ށ�JL,��[��SpʼzH���;��`0�	�f���1��������qV���C�(S�b$�r
v�d��
�=��XD��!sɒ�T�멵�����}L�yR|�ס��
��h�����(�hq�|3�[8��1�!�B�`}�QIި���&TWy\����d/.c��FC��q�[��(�7�Sg��$0]�X��'Tg�1�m4����R�m�3�W|��$Y��r�	���&H0>ӑI�c�_��/i'��26�{�LUIa0��ZO��;+>e �H=R-L��kE���d+���s�S���30���5�k(��B6PTt��6ni�i�E��uS��\6�ޒ��AH���TV(�"�t�(�n��la�r�?\B�e��8�p7w�������A��3�ن�#����%~���E�UjӨ��*퀹����\������_��s��Ј�`�^k�(�%M�ĸ�#�T�J
Y�K��YS��<w�4����7�D:f��"h�� Y=��v48z���R��e\�ǝ�vT΢�����\��8&}�H4����P/��o.&qΠO�b[�f��-��aԀ()B�;��A�:mݷ(�畨�ҧE�>���-�D���9L!�6�� ��� {ۃ�2�)5T��22[䜼�9��\= ::D,�^��t �\�
�µ�s�I�Y��ǫ/ ����Nc�р3�b*��+w�*�k��tu�4������*K�_��V�޼­~QQQz������,s)aH���L�T�=�&��|��d?��o�iyK?��8��w��Ԃ��=D�T
˕�� &c1�&���l�U��Qځce��n*�;{�N��^���}��v!4O��Z�=�5y���"m�-�����}�ä��6�LU��+���:�FM�(�0��"�B���N�?��1H���^�Q쪀r���k�H�a��*+��C����1cB�4�,����fI~�G��R��;oew�+ؽ�X� ��]F(�����x�����w*���C�,dޚ�-M�\�]J�gNI�����gk��Ǌě�^,�}R��D�ԷA	ݗ�x�-�]Xֵ�w�@�g`��:h0���8e�����RI�+���"qYz{&Y05�)$�\&{'.����"\p��c�1�S�_�n��^Un�8�E�Nq<�!.=�S�7��7��)ca�r*�5
0d���O(���
�L3�ּ8Zʘ������8����>�7o��Mm�x�|�u��Բ-Щ:���i}b����	a�n�>�G�׸��wW�e�;*m���YC*���������;}]�#�ukk�@�,$�~������V�/3P���O�bo]���֨��6ZҞ^�Ux�>v�}�93�OY��a�}��ѱ������G1�̀��_��H2dH�ۇ�"v��?p*AXb,B��{�7�g��4��l��#`*�S�-�M��7Ƞ��׊�?�ؓDmi^��/�8f(�7�+G�)X��l%�Y��r��L�B���  ��/�U�]��D��PK�J'�X�Ӛ:F�Q��S=�߃c6��*+������� �c��a.���-�����S\j�n�p���&�vX:ޑO�Ɖ�	��&�k���I���X{R�~ȣ�� �9qI�����⾹���A����������A�����O�{�M�d��f���!�`���kv�s�Z�K�R�d�C3` ��`�K��mM(��27;��R�f���\��K�9��ɍ��oQ��L���ݨ��W����+�qd����d���x0k5ȫWA!)�{���/���� tz���?=ZĔ���
"���ug'�������X�|�IvlD	4����hk%�<KK�|�$��� C�͈��e	W�t��G�|�B�-��KC�@�s�j��ν=pئPsl�6/�C�Kf�A�^t��[���䲂��?6���q\���t�����Z��g#�����م�#<�0��&7����,?�F�|���� i�bRS����������[�Y_�v\�a��A�hܚ�յ�";G��R�icLS\O@��p �Tn�����H�{&N���T	,^\� �t�|�V{�Di�L��$�=MVm�S)��BI�y��=���,��/`8uG�3����v�ȃ+C��#dɌ'� ��;Ja-��Qx,�.�|�f�@+Pk�l�ڳ롐_�/�7=7�9�`�E���m߮��4��>>Z�����f�c����\A���j٩8��Y�N&�#�́���)�F���VtRpt,�iDv/5�9=������2c��O[-�|�Ь�11���"�Ӯ�m�K�A8mI[�^`̃	َg^�r��Q�\����+���Mz�5�>7d��l�҄MZ�n�)�B��)Ä���c�x�	0����C���D�76^uK��G�x�]O�p6���5���ݼ�X�ϴ�����jY7�>V��=b��pޜ��u��/GC��e�Qr�n+��2es�#U��y�;�de3�cS��J�.*����h󈊃�[sr�,KYծI���!��VW����ň��."#lf���\ǹ~*�m����
�訯F8�o2���|��A�Z�X0@J��T���EW��ч�g>OQ�Ke��T�p�O���]J�^|k6���y���1M�r�� �:�Sau���U"��E�4o[�!�.u�T(���F����� �����=��^ �:՛؞	�گ������{pc������+�S��Z�G�L�_�\����L�߬W+�CS]g���(q��H�))�C� r�K<���'��(9��z����΀1{Λ5�o�";��͹��������J�qZ�ͫ1�[����*z�̖/C��r���(�rp�u`�O�L`�0b�'(D#U��f��`��P��֙X��$�I�ʪ�	4�g��߻D�&���3�ө{��.����7� Au�yh��CXz�f�r~���_���m�]!q���a9�c���O�p࠱�zOLO���Kfi\�-��lm�V�x٘���Ϥ��K���1	&R��f�È�ģZ;����+f�,j���-�HFF�0�w~�^ ��V���U���Ku���'�f��\��gGSɸ	��;9�j+�uIU7o��`�QcGt<�.����yAk�w`H�$��GIPk4�Z���;e�����dF��������4ETUy��٤�L)�r�����T�Wl�����L�1��3�UT�a)�,���,��[8��v7u�h5�.w��-�4qw��Tzp���01�\�=�; �"��B���Z����_TP�'���ș�w�M��iTʒH�C*��y�m1�64��6A��ax���:f]�na����13��Y��&{������y4�����X����b� EH��E��.�	?v(Vd�o-�J�_��Wh�j�([���zoDDf�y��d��<ҠƂ� �<^΋W�
jR�`��DU��=�
e�ڼ���R�	x����$g:��tKI0���9G��Ʉ-m��]��=�lG�YQt�����Ȩi\e(��m-��	q�8*��-WU�B�oaT����B��7&z-6�[ΐ>�>n�V����@������py�³V��V��^���Ǔ����㪌r��ʥ�M�+�>XU(�Џ%g?)ڋ�	�^����cwʐ�m�n7��o�%^ad���Q )���~�������b�3a-b���p��o�KOA����?��3̆xN2o��Ya��cf�g��$[qN�@��x�@(� �p�)��2���.b]=��l!-�6)b�OM��:Ƅ�O���~�W��N)�K�Bڳ�5~#��P�������Ƽ����A�~ٲ�؞Eg�����mͲ�N�*<_8�4?������u���s��/�1�^��9"3|{'���23G;����S��&�6C��dC\�Є�z����4�_t6�6;�K��es�^#���rt�;���q&4	@�J{�]�mYX�eV�I
L����{��'�#�$r�]u�jױ���܍����������b�+a��u�E��p 	�����8-y�LNTP%�� "3��8Gפ���$��y�q;0Z���dFhB�Cg14z9G�K�YK�6��,E*���������2?����$��bϼ:�b��~Ȫ�3�!��.3/s<,��0C��eԳ\�4I������W��)$o��u��T58_�Ğ��xF	Z�
'MQ��=��	r9 J�]^Ѧ}�Y�� hwп#x�Ό���K�P��7U����x%ރ���7/��_A�,�B�k��f4��n�Qgy�w/p'�쥲��\�A��]�,Rm�QU 醛~��-�����Pv[��>��C���3l 72p;M��D?�
bm�,���V�t�8�[�P����tP*�H���hƑ��ӲR6�Ǝ��V�>W�:�JtJI�*܅9�iIO3}��:U"�X"�Xo�r�}��d��#L��#���.#�F)��nk�N�
isp����]����Բ�[W����.n��"�����T��ܿ޾�`CQ �{Ň��n�_Ʈ ��v*��%�5Lo\�E����H�zX9αʜ~�C4,o�w]�Q%�����V9c��~k�]\)�
��-Y�Tc��N-|c_�6���"�rw�CН��/ ;�Fu�X;�g�u��ua4#��r�o��"m�ݞ΁��F�\�x���m!��?4���3dBuB7λ�3�^�>7��_d�wK��SԳ���=����A�h0��t�?Z�;�Cd�bt|�ׄd)I���?D��咐dCJ����HPj*��'�%�֡;�3�>68(�9r��i����Iʅ�@={W�dqX�	��x�Y~s�H����yF3��C.�bO��p��"�v���|�n-�+�qy��*��(,�Nx6&��=x�0�a�kK�#������+CW3"��H?�(�H�z��(Q\��>�r�M��B-D<J$��}��Yo�����1�*5h����p����Q��ڿ�$�G�<��mmu���S��Z��ɖ�����IY"6�P���G�IqI�9'�g#6���?!^�n�!�b"_Ь]ҿ�<4=�Dڸ����4.{Q\��1�� �6����_���] *$@����B�U���]�3�sx߂^㚓�=��#�����1�s��l9%uy��&>������x����� ��Tā揅�%%Aq��� G����'�6;���Y��ś��x�$x�_��$�K×]xv2�14��{���th>.�5��W�Пt��Aw�p�����LsoRM��ǩ��t�Ż�$���`lg	BK���M���*��K	�	�6�G5�\�6*&��o7�>���>����|�KeO���Q�BS�E?!��PS1�v�$�s��xG�+�Kݮ������=+�{�B���u_��t]E~��Y��'#��9>�b��X_ƣ����_�[R)�ՖO5�c��&/u�
�����N���yg�
�]�q��y�qA&3f����hI��9�\HD��e�
C�'��O��W��yty:��֌2nRH����
�m�c㲆>��mlrN��WE��r`�&���F�|*پ�.4Ӊ{}>�8���:Ħ�Dؤ�?�_
YzD�^^�mӸg-����5���}�x�HL�)���^����P���}Qa�F>��_�AYJ�� vPa&�P�8�n���9��]�/�vQ���V�Љ����R��ё�R��D Y4pU�
�ʴ1��&���:�.u�4�����&I�l�m���1"+4���:��3�,4�Z���/�,��yY_�vaP���o!�wog��m�K�W%�`��[K~�1��q�U��`�l�X��Sč.��*0&���$y<�?#���ba#jC��v6�Wϒ�	�lk�p�ȣ#R:�������%_	iL쯽�Iq �tޢ�j��,��U$��f�o�^� ���A�v_��^Eӟ�J�= �{��e	��Q9�c��\��2�"RC\���sytQ��������l�p&R��5އ8#Y&����f�P�8�/L�/�O.IB�m�6{?v���[-�>����C[�?!� ;߲ryZSzL��x��S)ݾ��:�P��9j�:���o��d؉22F y����R$=��"@�mI���`0P�F��7�+���k7EX%O��}rW�:f�Ո�B�`�q:���`�ly���V�R����r.IC{q�oA��g 
e�>]4g�O������a�{F*��f�~ܜ.>H�>)B9L<U]2`�Hr.�IՈ��L�í*�-	�0K�� v0�!+)5��ѯ�~�C���*ӠV���S=%Iq��ut�E�Z[>���`����a4���wm`wt�n]��\�i�4G��wѿO7/a�r2ѳ*���hh�E�:}�Yz��M�, �h�����s�״:����`3 /�=�n��gf�3�T-�x���raP�骅+��mǗh,"�!U�+А\`�M���>��V>B�� �FM[��.�����Y]�y?�v|�u$���9饎�ʡi��Ш@�ٔFxgKP���N?��<K��dz�����T���5s�l�*������~=�Uq>�m� �.��D����r�w��.d�7�FK���%j���sy�L/�{���(IɁ �@af9�/T�$m� �!���+(g[y�k
@���KB��-���eG�~��wa��.�G�/����+��H��13�=C�r7�즵x��lL���)("!�E�!���d��2��z�(�B}G��_����ɐ�ٮ���'��T�������>&�\�?$��{1[%C�)��=��b0>��+뉐)X�|��4#��=�g��4����u�I�V�}Oa�L�j�oA��/�p��CI�d�6���Wt��p����v$UD&K���~�!^�8â�Y�~��P}�����a����]h�{@�0N!;��f����O�ǹ�%�eu�U���W@���q�^�9+V���Y)�~U8���(�w�[{�����ℙ>z�M)Vu�	����2�Y�G=KD#h���;M�3������{��g�⿛��@���#!Q��#�8%~�mGA��6d-��{<|3�?����#�m��^4�����l���W���L�8���Wլ�^,A`�I�Q�[ї��@W����`zEL�p�`���Z���p���(�]�C|���k�CiN��ɣ�z.��:Օ���m�w;uUŌ*J%(�c�+������W" �Q��@w���J��@�'��#�B�o����T��� ���E��u�]:p X�lӈVB�o�������\$҂�1�����=�3꺳cL;�:���bw3�xwu�'�^&+�j�iׇS�o�%N�s�<��v��J�0�J~��h�_��,�mH
������	?�h����cs��m^�p����|�x}�q����ߺk_H��CkDm�m�M��>$��!���;5�W���TҌ���
�gJ�c|����x؍E5yZ1"jݘ�F�|lDA�9V^Ȝ#:I��D��d�fҼL��0;�Vv{�����F�J����8�OƁ��A�2]�Vݙ������f\��H�a~{l=�
�֋B�� QZIh�n�<$ W�~>Zx^pcԋ��@�a@�(K}��z|A�<|r ���|-�
��>����VC���֮Y�'��~z�6\s�&����~"��*l�%��!'�d�aZd����7)+�$�����#�UY�P�"8�9�������P�gZ���uv0�#�=:�4�������d���AÜII�g���uѓ;���5�=RH�,58�I�rU��k���+Y��v��V��j~A�35E�iKUx�E~W�b����b��rB�,�ѡY|�=�7�կkz����O�>~Đ�hsU�311po�9����Psϕ��LqD���/]����]�º��.�k��|\��X�|��oy��c��6&�W��������E)���s�_k�Îʞ��q�R���N�&�a�>ȝqeZՖ9*����"0�b�W%�����ݸC�d^DKC����8��	���z�EV����GI�a�y�pļ���<8����h~[�b�x�$b6��Fa%������Qe���8�"k���%��Lت����GQ!��\`M�з�[ �(�)*��&I�'�X����iHN
l_!�X���%6o��	i$Q�W)��M��	I���1.������s���O6־tge�7I{���8ߺt5����qde��֖��D��W��WF2A�R[v�}��ͅw}�h{|��O��LK�*�C, Tg�e=�h��
\o�c3WiP��X<m+
��`[�>��qɬeJ����\V�'<v���c0V�lۖ��B�t}��\�̅�+}QO" ]Xcq��؁��O����Z|�f�'e�F��������.Z�~�HuFW�D������Jk����b��g�C>g��]��=p�4�&�ng�PFp��9������|S4�~��֨��W�XWY�)b-CH��F� ��?�Ss�li� \�2�i����!�G�'�������P�Kj<⼀K����ލ�N�$��n-���ǅq�D�� ������8>:�KhV'˷�U�hJ�r�ISmT�sI��w���2��Dw~��dEZ=R�l�aDQ�&����n� �K�_5z����KE���A�uZ�Z���A��)~a�o"28Eb��o��$'� UK�E�����O����5FE�?�x����ب��R��1h�@,v�:�����>&���&��S��?���؄�6���D^��z�
2�S3km�!��:�㍹�q�"!t�8�T&$��j��'�YnG�|���Æ�j����Ǒ�&`�"Pއ:���N#��������*X�R�`�ӼQu���V����jE��&o��T-��:<Ƣk�a�#�����v:��s4h^���:Y�"���;V���^���/ G��ryϤHH���^:U�[
H�GV� �s�㶄jt��o�y0|��η�]�q��?K���1�i�z��
R!L���Qd�� l���q��`�Ya(4J_�gD�.A�����|�����P�Cl1�k�QE���_lhEE�**�^���?C�L�"K��!��֭�2��Q���P���ɭ(Cv���ܥ
C��Y��%N$���!��-�h���4s?�1�f�Uʑ����C���ƛ�r� ����/f"1�0�M����u��S���ش��;]��Ec7
��=�g����ښO��lτVଘ\�"�/��j�6�i�m�m\�'
�\Va�,��o$�/`T+�^��#����W��F�7��ĉ�ď�KH��A(i�Q��d�z����!�M󗪒�����9�m�����O`�vB���X�(��3�_f��m٩C��Ǐ���<�G<lޯg|A^m����VgC9cVv:� ��Ӌ��eH�h�ф88�������:��"_��̽jJBtr��j����]z}i=��Je�Ԗ�G]ҷa���)7���|�.�Ԍ���/��ןu��/�H�$!���X�><�Ϸr
�ҺTN�����ՠ�p�a?-�D� %#�8���N�$W)tE1J����lsx�*M��?E>_�P�<���A���A�4.(������H+���rv�. ���I`�P$e��સH�eG�*�U��j5�Ќ��� �A����|�X�I!Rߚˬ��C��v��t�^����q��(��EV3Vh`#��xh�_O4y��J�Ke��
nɺ�ބ�v-(�й�Z���i��݅&���� �F�(J��$+�l��Yh��x��x��u��B��R��B~����_̉
(��3�~�i�gX���e��zIk�<3%~�����Shgu�>�!�����#�ә��(�ҖĀġL^=�����Lƕ�����ɾ�Vr $�i�ދ���0D�[��0��8�	휗އ���\|�ա�;�ʺVQWǚ�w�I1=87r<�#�Y͎~�b��|��H8O�v_����MV�v��Tp�����ɤZ���"��EX�j6��,⟻��������V��� ��@ UN0�T�́�IAT$��|x�y,*�2=�|Q%��T��GN��bs�Y�읆;�9K�1.C!zTZ0*r�S�����N�
���W�z$r{�d^X��m0��8B�A�]�m�Q~S>׺G6]}�V)�_Oe�HgR�@�p�T����Ly �� o��.���!�M�-8�`��%k7֊�%Fw(@P�)% �I����A��G���j\2l����a�웠�Z�����6]t�N�z�h,W�`D¿�Fz��㞬��%"�A峦�7D^x��\�;i(��σzCT��[�zce,:3�<�̨4pv�]0ܚrX��ށ|M��n�|�hܯ���xx�˹��@��^f���ﻀPS����	���{>��J9�����4�m��>�z��;9rj5���� ��.�'�0����#ĸ�AM��� -�������%us�"I5<cJ� 
#��\�#��Mà�n-�2qTp�WD�w����qu79`�a$ ��^�2���=aR`���=�^PĒ����)t����J��t�����	��c-���s�>���LI�)�2���lORr�G����L���)�����n��^O���`���}��1WZ�5�C@wX�^�w7Z��ID}�"��5���5-�˻p��2TYM��j���|Z��{��<@Rs9�-B�����<B�ˢZB�U������S�ŀ[���j��N-��V�琹���7�~�疩;�yA�ι��c���E���4��4-eD��a���N�s9'"�$Ni�I
�o��;*��o
v3���L��y>�)����S)Q��WC��l���U�6��<�7��ީu���L˘�`ւ�3<5�Z�ÉyJ�#zf�J5�����VS��8~������id�C�<��B�@�2�iY�ɗ��]��0F)� �dGS��_* �pFNt�h�d��8��}�O�p�)$�c�v�w����E���:3�*Ry]�,�f�sa��lՖ.�!��W��g��	���͘d��xI�g�j�]#�̜n���	�j(4�(�W��9�1~�)��pGS|���1��dE����7g$�V�~���: ��&醣D\]��z��9͓�_q��^/y�u���@G��R�<�������D��L*D���I��!���?��l�s��gp%^N���d�*j�ç�ϓ���lgO
������!`[��/�K�F�N��
p��Ԃ�oyf�r�g(�\�[�4��*Ὼn�7�ur釓 H�Z��C����f���㉓�NN�q�qb����7D���W}��-^��xm?s�H��T_�UW�%u�keЮ��`z5IG{"����W�E�$��[	� ��)��zS1am@c�Q2t+���S�ʹQ�����KI�	�h��"E`k�/	���)Y=��m������$��Ɏ�&���fz���;�9{�KH�+O���XA��@�����0�' ��u��CZ�.�\�qvElc�:g�z6�]j��As�Ԩ�#��7�(,��B�S-����>�(61���9�:���
�#��A}~YQ��|I6}Z�O�^�e�� 4��`8��i�d�%c^!~$��J�O����/���>5ڠ���7z�nA0�u��aG�#�[2�q�+�d�`��p�h��)�p2=�L��6y�p)�V'-Y�����/�����+���/0|W�y�R@6r ,$	�5�`y1Mˣu�����?F�"��=nekí���T�~Z�X���jҠ�SRh7�6�4��?9ۣ�Ћ�iE؈Lq
�Lk�ȘM+����?8I��l�{O�77�b���:�CO�i��#M�N\��6n.kG�-[�th��5�Q(������ƒ�/�H/�u:1��#ȧ�D�+�P'��;<��;H�O��~q��&X#�þ�J�[Ģ���|WGs3�D�Y2T�"	Z��mChN�4���&����'�->�T^���d�y~�'@�iaڹMBǬM��Y��獮�P�p؟����gM��vH������<_V3"g)�#���D�?�/��D	�݅�"9�"틺�U)Yh���l���zg�Y3q���moԷ�<z	��|)�M6,A�r>-�M���R�7��Qh��$ȡ�!��8 ?y�]Az��،X]�jp��,ĴM� *���ra���BS^�q�]=���[oc��~��sԏ�b�}ت>��)�j�8�П����J�Q�x�>DE()�&�М�]�4k9.��U�	�=HkvZJ��>�PJ����r�r$�X����L��؊E������B
w��SCr�kS���L]��.j��೪��cik���%�H����I]n}mVĩ6|��x�:(u鱛�嚯���O\�J��@2�
���7^a"�X5}T✬��r!�햪���A
U�MFX���݌�?���
}���'j}��mZ���Pl�Y�e,ǵ�5�@�<��r)��ˮ2V%Wʧ�9G���J�\�bx�O�`�Uա{bA�G ���%��A�~�	�'�k~��J.h�{��h��Gk�m��*E�<S��߿�̣sU���h8	��b�(t�
��i���U�X\N�88G���]�-w:��tjd�Fl�@u�\�����-;z!!mgi̽UmM��Z60)�����w�_�w0��J^JS��^�ג|\w�8�DM��V!#�E��U�x�za��b�YZQ��d�� f��>���,��hP��.G�A
�d�cZ?�b0E�����r��@��#��  �[V�PB�$}���{ܳ|�p�Q�H�r64�a������![��qLMIQ7�w����]ݛ�ns��Ã묂�e(�R37����`������4ᦨ*����.�ʵפ��W�㿊z�����%�[����H(�7�:x�$�F��1%.�#	qƄ���f���,�%��5%���!y��eGD�V���h�����na��c���B����!��M�o�Я���=q0����?�M�1������z�Y%��.�[��\�ly��6j������74 pJ�#��.�p͙�jCU�����t������y�޴MGB�]G�u�s���p�RuG"z+([���$�_:nȖ��c�e�
D�*�7�$�f�()$$�Rn�<9{U�u�f�~u��ݚ�N4�[>��Z��{7d�,pv?��������;*Tt�5��өL���5֚@�qT���K��1�A��:|T�]�� ����CY~�n��g!l�g6���v�1���uT��h2e�?k<��C�����Lu�4�e�ی�2S��^]��3�q��7�	�tMA�e�˴4���@&��=E9f$�V�ä�!���&Y��\��woh��󑲂�e�ɦ���-`�=��������ZܦC��ǂ��Wݥ��U�L�-��NizD*��M�X��JǶf���q(������g�)o���-�]�+�*�HԐ�H�`�k�
��ph彝	�'~E;��y�)�2��.x�7�1'�������l*`oZ�P�R��:�k��#�^�v$��Zj�-��-u����2�ّ��s�kVR��@g�ڔܵ�U 7`�._yZͣXG9�_BC�0�{���f��/�'Т��U.߅V��#-aӄc{������t��I���;��]���ϨE�y�b2���F�$CV$,�{��2Z��eW�iAN�|��7�	�El�W��#PU$�W�G�hq&Z�K�"+�A�C�[r�C�_:C��m
 ���\�h/e���9W����b�{$а:�ʮĊ�,Ug��]��,�I;���h����E��v˿]_�8Ѹ����˜..��^��N�Z2�z�</�̿/  �`�/�e)&�t�zTv�Lp�9������&�Yd��@�:Bj�\`p�9J��p�Un'�;��2���.�&�e*�@
D��ƥF]V�|J��V���4Z�e��Pb+ߞ%�w��01�~�;k���sޤ�bw.�r�܌��@l��,Au�$��D�ƍ��6����HAS)流���cX����@*����`B��Fi���%!NWBh��=A�긃6G���h�l�|F��{&%r0���d��+��������p��"�����F��Zyf7�tǥ�����B���߸��LS��z�c���f'����o�O`eƦ��2C����d�������4�a%6�H����%���ل�{B8�s1,�!�A��8��d~"fl��Q�`1�+������{}F��0͜K6��d\��O,��3\͙�^�P�+}QTD����V&���+#}����m�G��	`T��>%�zR�댶��]��!��TЈI�^�:ioŋgb�����%��AÙ��f%o*���\��,5SS¦O�֛}�l٦�H�^P~E��&�#FJS����7�G��;���g�R-��ᒧ�0z3��]�]n�.ΰz�%����lg�����uEv<�O�??zM��r8�HJ�E�9Y饖j"�46?}���?9Љ\K�v�b���5����7-�/�UK���Sn� 2�æC�ˬ�����?b�KX�F�w!��\@�5b�j���t�٠�4>Lq]��bB�'�PK�0E�+H���{����4F��$Ң@%n1�B���K#噔U��/��� 4Ζ�Ç�ֻ�q���>�'F8h�Q��!��$q�z$�u�B��Tҏ��,�[E�xp����d��R:�!p�|�Ih8SҢ�x��x�G�҉� P�K��*k�������EjRh�����fuXI{��m�������U�W��@� ���+��<��)�6�0q&�J
��[�ǰ�����7�T̃����'�8����C��Ψ��[�f�W����� �d!"�ìNj ��Q_�:GwI	�G��c¾�_�B��>����wn�A��K6���7��R5p��ϸ(��R4�#���}Ud�zNaN>U�%:>�Ȣ�X�p�u#?eϋ*�۔� �v"�|ԑ�aҏc��جKT܌����SgO�0KF�*weY3�<�V��/C{K���)V��8�mp�e�y�fd7��.�U�k����%L.�*1%3��A�$��P�K��0�PL�m��F?�H�S堃sj�ǯ�P>ޫD0��9����S[��%l�/w��%��w���
����f��\��k5���U\�G6�7V=���X�[��w�C����q�=�m	�$�ɷ�8��S��-:�r̛~��_*t��{f���s��^���S.��dEy͞����;-��\12��S�[~��8��*�^{%�{�P�����td����8� �IX$N�s	='H����eß��q�d��iՁ��QʬG�۬PǟVy�(�� ��$0��OPI���p�Toˇh��;�jon��Vq�J�@YjR���v���ĝ�qFr��K�"��w�gyQjp��O�7o+t}��Do0���p�gA'ƙf��Q�E��:�����{k�u�8|�.�W�V��k��A��A	��0+/g�)��LR�ǂ�];_�&��<�sR�NN5�:MԦ�c,�8 	��"���H՛&	*`��YǓ=��Q�l���sl)�`3�nl�z�h2S�7���V��I5�o�,A���#���`��ؙP����.ԐM�_���ڴ����tCվ�p� {��j��-�[�paUW������UKNˇ&f�t%WRM0(���p�/A�D��M��r�,%Z��[3����X�C@V�.QB#�4�e��g�
��:���r���(go���fp%��zX�c�&��B���Ւp/�A�b�k!H�Lj��3�	��]G��}��1 -��>�)��5 ��,�zK?O��.�v8>��Z��?e��r�Jj�qa�A�)y���0���>���@А8����Q�.Rq4Kǵ/����"�_�Xд�l����V�j� $���#��D�
$�/�B�oY��wD)��u��:�
q��	�Π!��49� (�I�W�}D�%y�i�Ĝ^ =d�Q3����n9��w�ްqĐ������w�x��Q1�Xb q�<S����h��LPʕ��x�	(��b��5T���$�?9:��;[T=V����ś��@`�D�B���͢��b����~��m�;Rm�������atE��S��e3�7�3,�F���{r�Q����C9sG��&5.���N&�&d��: �qzw
J�߆����D�67�I&��.^�ϟ��40_��m�'sb�3WAo�tI9g��"�)��q7�'�m��K3��f���
$�4P)4�z)�A�P��mٍ�_7b���\f�IV�I\�+Px�yd"�cow=�2���6�HL��~�r��F�ቛ��'�;�V�p1�|y��?"�/x�a����]K���L��=�Σ�2d���;�v����^۸�r�;��&����.=��;��F�zT�ef-��Y�0�Kq�sU�nK����Ϫ�ZE�n���DDۥ��q�7�z��u~�*V���ז��J�kw۶�K�l!�*���V�Ҷ��l�Gh��ݥu���^��_淽=�����DC����	g�w#o����̲e�i���3usqH7<�Vo��9���H����6�ތ�?��Z�f��|+�gl�ivK��k��+˶��V
u�����+t�SI[	�%� ��BdC���׺4��S�`8�����M��#©���jƺ��\l���}Z|t%��#�����Kτ�\̝Lښ��9+�3�,'�!����v��|D敬_�_1f��j �qRR��e��	W�4�_����TaFg�=�"�@�)8��g�95��a��W�ۏ��F�}) ̯�<;Ζ vBI��u -� �i���~.�ِC�|��K��������e�k>{t�^�������;x���߿��~�[��H�e^�tg�V� ��=�r�ً�8���U���ֈ=J,�x�
���@��bC[I�QZs�4�'D�RP<��
���0N#к�/�O#�e��i��yOի�}#��T,`�2t-ڇ������i/�J��"�u�뱸�6�aG *���5��D!5-
��>�m2��`��C���D�Q"�A�y��90�|pԹ��^K9Rf`�]�:W�g����L�{9�_E���;�5���T��n����zWy1\���{�x	ְ���`�S�:ѨK�n�<V��?���[v�16�d��m'oB��?#�lV�h�"	�"7:��}�;�p"ԑ��X㛥ʙ7"��g}�"�Je�3Vޏ��V�}���	�)��;��&"�i�:��_!��oVN�s�@F�K�t�_]P�
����%�{��!������]���`ZG>��߸=(�$/Fw
�"[&�� ���!���
Nʔ�7��M�_���U�g��=��/��9T	�oZ��[@T�n���,��5���7��&i%�ǖ���R���6{CE�k��q����h���S�۹���ST{e�k���v'�������M�)�ܨ��ͪ���2۟�2��Cb�3E�"���fAU"�M_��$E��n������@��E�M!����5��-:���n���?�+��"� b�z��k@A��L�����E��h=�h<_�<�
��_��	BgPr_'ʳ7�{����<DZX�F����0���P��QGRkՕ����R�Ꭽ(c����5U�$�y�:�4�$���-+4��e��<��F��FX�0 &͓N{��>/�����)3P��W�7�WDS��Wz�~055��ɔ3۔�&"	H��\0P�˰l��#ޙ=xP8��\��b߼_�\!��Ƣ/2��jM�=��ḳ'���7�d2TJ��9�Om�wg�>��*�U8��`� �׳\. �s�_{Ɯ�7����S͌5�7Q�������ޏ���N�A5�,�!�#u��¿\:��K���5�%y��'m������z��N��p?hG �d��$�q�#k�A�[CE���U[��*f0�n�����}����#�\b�'S�긦�{9��,���U�I�s�2*����]0Q4�d��>��]T������z�yK�=����
�PSh��=i���(����#�<�M{G��Ne��D�"=�Ӄ��巽!�U����t j�fSd�:��U���9j�4���%���gŁ��穽q��N�d���>����-َE����_4����~H�u��DI�:|�L�Ҧ�#��ղ�1u�s��d����(�.aD$�O�U1 \����R��j�3��
�jc˕������C@�bI��� F��|�T�_������  ��@�.�Z�=�D�[&�(���������RX�*w�=o�0(
���<����hF��2K�ڌ�����SW���2ܨJ����ʒ���D�1:M�5�%�6�̫1E�R���y�;��?���:"8^>�Ÿ�e��(u�6��6������A��R݅_rB�H� �5o@& �H_4�ş�q��e`J�d���;�B�؈�
�.�%k�	hW� 
�,���2=���M�7~���3ɡ`n����m��Ͳ��#S��XҨ��k�M�%�:����Ir(Kޗ���Tީ��_�}"�PUd�_&���!1���!C_��*��C�b�'b++R�T��k��x��JV�ӕ=�0��
>h+uQ�#G�/�U5X��*>8�q о+��%[�,�p?��1�&�|�͓1L�Pu�>���Z���#����p���͜еH����b_C*��\~#F)�S|o����sМ�}Z?I��l��& X��/r9<��<��4Lݕ�@�@(a�twz�gK
j\����&c;h&��h�=@I&6W��� D�e���AZ����X	|�d_#e5t�y~N�~�mk� �ؑ'��vN)����w�VXY��vK��a�j���1�,��R�G�c\n���;����L~ǱX:?����gˊ��:عe��}J?�oE���5<�&Pt��J(�K�Ѻ�j�����GX���K���^VN��\C�>Kf�������� @��{�
R�}�ѻ��� 0ؖg�Ja_�uj��»�Qp�Gj��"p[sPu�;��7��kK3Be�!dI2��y��h�P���~����U}�#���:�/��B�s�J(1���&��&p�ްz\c6�ý)�~��C��mVV�j�A��a��lpT>�2�H[��0P�Vx#%2�O�/d�	�������Ga7�t^6�|��Fc�[�E�u��hP�@.r8���O&aY@�}��7p
w_�q�fv��� )��V��*b@��"[vH�x���#%�اI�|S�$0�@�����p�9(�wҔ���R�Jv�ϫ�9K��90_?,u��l{,�ņ���C4��}��׌[	-��S[�[���0%��t3T�c��=��+d]e�%t�%*�;߭J�O���N+ݿ���!��ʇ����C��s��ߌ	�<�C������ja���lK����w��%(��Yu�A����Jn�&2V��N@��|F�&�2�]ةC9H��H~�*~(I>��VZĩ`��*� n9��:�v���8�L�k��>�6�~OJ���'@HSX��{>��������<Z�Fn��r�ڋ��*�5Ú��Q�2*����Aٔ4͔M����+�Z�$P�C�[��#�&�耟��cApɚ�|b��nP�(k����X��;���Q'�,����W/�iۅt/�3N�a�Q��,gA���
9�оu���+�V*�T���Q����r2?@�y��ι�<�IW@j)����OxQ�P!~ʕ�ﶹ`���%�����f[��_"6EI�o�`��5f��.HZ�,aQ�Mt�:�2k��W��'�/�ңz*�`i�d � o۔�������굃1�rLO�.�}�3 �s���_�I���*���Q�� ��a�0�$&�`��|�,��řa�K����Q��G��-�u�n�~E�iCA?��p��`:�
��8�f���v��e�ɧ��,�,e�;��G�|���\ÄM!�/�ϓ> ;�D��W�6��x5H�g|ɹ���$%�I��xϡ�o�7l��'c�=�K,U���2�oN��},�X6�$��+�
"Z���.���(M�����|7�J_��ڕY@eι�~��c���C_� ibU˖�>-�"ۣ���$��t�5��FF�X :�Ý�Ϭ����Q�251�ϩ"�0�%� 3�,V���;-��N@�/އ��{AJ&�w��}n!a~��^ZZ�i��E��?���A����3t/�;[���?�����u�5ڎ�ȇ�����Ay��Fz=�>��[��&H,\��*y8gƂ�1���=�("������ ���F�S?� X��h�*��T(���B �j�٪QCU�C
~7%����Ȍ��c3�r2������uXX��A@iK�9$E��m���_�L �'�mC��.�ix��tVHD�hUr+�X��_rf������5L��d&|r"[�MxK@�3D�`��0�69�\X(:K���I�����"5ǩ�)L�/���5�I6��;��eY��Ն4$I}���zZB��<��\ٞ�&���;�RϡEx,ހ��FHC�����:� 4u�C�����!b����5��Wn}�"�$��M��U[�5����n����~�}I����X��P�&�^ �o���;�^0�ُ��A9�p&���}����y�$�@	͡����1�fO�2�쿋�,:��j��p�]�㓤f);
���I��S���4���d���],���������f�a���i��l_]{6��BA]X0گ_�{��SW�k�??�4�%���(�t���tʝ�@��a�k�i�BX=9u/m�%G������i�M�V�k~4Q��X�J�#�I�O��T��Y��X�]�
�H��v����:P9�f�U���7Ah���-�������u��`�_'��x��hBNVO����ż;��9rw	�Gh���Ai�Kh�\NzJ�k�゙�{Õ���I��>��5��
z�j��˔\��8���������>N�1������Y�D�1O�2b�ص�uG[����ן8n�*�i���4LW���b��+�)�H��� 靂������^����D��K�&���{'�y7��7^v�/yhf�̆����μ�9�i�����_pSI�;���Щmܖ����7�~[F'��(��G�tN���'�˦�ԝg=K�>[q$/�vF�
%b������˭��N��n)8<AA���1�32�X����Qx�bB0�~R�k�v31��x��ʶ؅�D�Ԍ���Èi�� �$��&�\\�_Y�C^��d�-��-?/Ů
�\>"b�8P����Wso]ᛸ�?4���D���g]���t3^�P�vL���3�����7�
Ԁ�Ӭ�������>a|��_����iBu�e4���<�������WtS��A��s��f ��,�ٌf����@l�=]��������i���?���X,����}�i��>*�yX�騬K������!��V��|jo��0�\i�GU���kG)�h��l���p�gpyt�G0Q���8q�ͽ���6��a��Qg<���� T<�-i'�W!�FA�1�'!�C�)�#5?=��x���3ȶ���} ���J�ΡY�9�#��ݟi<Kk�F�I�Y�.�5~�YQ�>i~��+�������)xY7�36N�ۇ�����< &T�<�b,\�C0�$�@��kDா�*џ�|��*e�ǯ<v��=KyȐB��)k��mH��I����/BpG��#�7h*S��{�6ēX��Ϝ�1�NJ*��<p��z��`!?浮f�l��h�9��h/nB�
F-����`5��YA���ς8��o��TۡbK�N�'Zր�M�c�V��P���cw���\�'���] qH�H�?]��#(�S��Vq	���E�T4]����-�pA%ab�>�����,܉�b3�g�K�2���n�kj�jgQq}�Z>�����_����T1U��%~Q5�m���z�����w���v��|�Ν����a�����E����u ��M�O�3XB��PK�	�e>�L�R�����c��Y�{�m<�X.���$!���gN�R5�`;d@.z��� >�������Ɨ6Rg��y.����_��8��FTD<�mQ�
x��Թt�0����Ao�F�r� g(q�*�i��hP����2�%kvaݻ{���V� ����
�y8���ؾ����)ӳ���vik����H2�N3�r��.
��_ ��x�.8�j4?C���qî��rrw&;(��9�եc�Y�? �S�1��W��^ftd�OX2V�H�#�욽��t�|�bgf��D��gf�O�����>h2+4Rb w�ik�14S+�j�V��oMP6}{�}��k���A���˅��<y/�������2C?4V��@B�%H��H�Z�\�Ӑ��UՀ$(�fGY?� K@�5�j����b�ç�h4S)���U%zsy��M!GAZ<�os�tE�=��}�/�(��L
6��!x�1����_t1�7�;v�j�k����j�7>��W�9�P���/��1Z�jO��΄���4�ae_��\�j�*�{vd�rR�GR���a�W��Z�`ӣ�A��^S���&�����1ߵ�2^���Ű�N��'fv�V���%j���X��Y�t��z�|Y��'��6H��/ό֞��*FCe�L:)����-�ftO�4�܅����T�D%^��$�?ۡ�G��;5�jW���
L35,/#�:���.�	"nrrg`B�������j	�/�Z��w��q�Cz������@���\̟r\mR���o:tE�9d�9�y�	�9"��OL�oN�OJ��lj���M)�B�F�Rw��pP��}����~Rc*�W���G�p����`�H�[�������Q��(s�8爐��,H����,�V��N�i�v"&���#2u��ˊ�D7�5T��TG{)�%VeS�<�moR��RrN:��U���L���cBT�٪���m6l�x����'x�'���l�QF`�Ɂ9���v{�H �9�������(ΰ^��J��>�e��S�wj�>VUe�xnܿ����D���zV�_�)�l�ۊ%T�Wol�B�� UK
�	��;[n�X��>[u��E��	UfS�<>Z+n��XKq�A�#�U��ƃ��!ُ�e�Rh<�[��r�k�٫��C`J@��k��BNdR�et\���(H����1����m�$߉:�0r�\��"�]q��8q^}̽�gc�6E��S��=��=T�8|����;`��v.w;r�d|i�'��y�ٍwvUz�ћx�	�7��߬���I�t~3W[�P9��r���4���@�3��\*m�H�>����_�#*1�<�$�l�R%5	��o/��/����燸�'\��:�&���T� 1�opڼ���̎��˧�K������h�����x���a��O�Y���,yP�҉�[1,S�g#5�L�V�sqe��$$����w�z�G0��@R��z=�z'a�+���a�͝�y=gʸS��ƺ/���4>�B*�Ѝ֩���a��֝�>�=��X(W�GO�nЋaw�[�6)��4,Y�O4�d�uwOZ�oHΕ�wu�Sm�w�F,f,�i�����k�+:����ǃӽ�D�R!*��c����F���n�MM8<^��;<�������R$��.7�[���5^�����|uPn�`�T��u������LmJ��̇A�Q��k�g�=�>/ �$j3����@�m�AT.��+I�V�^�\ݼ����6��#��� �W.���e.����u�ZDk������<�/P�y�f��~4�S��C�5~�ʖ�X��%�����Q,�'�J\�#�ONkmm�ة1.����j��xC�f��Qր�-��?����چ���r����|�����h���*.=�&f�Z�"o؂/��Ѵ��-P&	���V�R�Dpr�D�bH�)`�E�N�֠+��UM=qF�UvK��Ob�s�)P5��w���1J.l# �M��"C�M��=E֒џ�����#-`|��a�x` 9Fd_�w	(*�_E���а�+�o�Oם�Y���"���E�w֣ *��FFx	�Kh+��1m�Oc��.. O��U#N3�ֿ1���9,+ V"���s��"�m.��T��>]����a]���Hl�5|�� ��,�Ԡ8��o���6߹Թ5+r�Wc���vM���&�920|�&O��X\����:���/Yr)��e���R��}������*A�X��96� (�e�`$kI:��dϾ�?8M����wXы���g�x��T��%�� �#	�ھ�H{��5-���3���YI��{H9�v;��y����s!"��0�?h������pL��kP�a��ݦ�C���Y����jd��S�X����ٮ�t=r�i���F��O#�b�٩��S��/&���*N���{=;{4����'���1;�n^��}2�b���ͻ9O���s��2���z
4��4<Җ3�m�I��ҭ�������mDfMR��&R.3ԭ�+cR�k�b����6v�d+Oì��)�(�,��[��y�ѵ� C�2f�;��&��m$�pg��w�������R�b�-@?�3,�W��j���n�,�)���H��*��h9��F���VGG�jU�H�c���|�וy��L.-���s�#U9��'r�h*8�n�h��]7�֚VI�V
���K�- �rZ��`����z���	,�F�nӔ��.��>�?鷵d�T=�C������!���*���4J����˃�>�����ng�_�ZLJ��qQϒ
�'i1���L. �R\�U��{��"p����O���vκ����&�*5biX�+}-c���^�:��%.L7�A��8�J���� �Ȥ�~���ª2�=���8���[,�
�w�P�1WB�Ew8��aѪ��ݷZ�'� ���d��dP軺�V�W*"K�%C<�&8#�'Ma{p<'s����?"}@h�}�RM�r��Q��֯e�Ң� �|����+��0��qV^A_waG� ]B�,X�c�1a�s"B��5a�x�ز6�t���B4�����=\�db<HL�|8��T�I��-4��=�����cG���NL��� K��J$Ʈ����?���5�@�Ǧ�q�e�1|�96rGȑ��������31��h�c��I��9х��``Cs�z��Ӄa8V<T��o��גQ��U�n��6��x����M�nQTp@u���:����UV?#�ݦ�f.Ɨ�	� ��#&��hKf��e�#:VY��9�ҽ�o?�ST�����8F�آྰ��C!��ۗ��[��`� .Cв�Y�~�Qx�{��������
�~v���E/��}Ԍ���Z{�����$�M.���I{��w��ovV6Ȼ���[>�1�É�( ��Jĵ*���U	0Qi]�����b>^&ai�����$fD`�����k���xÇ+���ާHdcFI�D�(�c��_#.c`5i)�K8�?�ִB�Iی,�|���ݥ|��ލ���I_�p��is{�(�����/�	�!��z�L�1�7B�4u�`�z8���ʥw���\��w��v����L=�[��2+7�w�L�΀M��*�h���P�>�&�sEb�y��}J����H>|��������c�E͟F\|l��XZ�F�v�;Ě|�7j�,��C�b l��W�����
�l����n�K�4�7Q�]ۥCM��a,$E������;�����"���u����{�v%�]��G��{ah�5ő����|�T%�bz�K�c� ��r�?��3C�-��CC6F �uo##��DF6�e���-&j�"�61���j��4"sql𧈡�Ep�%��h�y���lN�Fc�B�w4���?�J���ZK���@ba���C������"��f�E��N�� \@f1u�� �2z�(����,���k[^���)�/�N�wv��,�����\�?�~�p�2Mn�S�C�l��<��b\ לT���[dn�q`; Q��� YtV'q Rp"#+��U��sR��bp��?��E�}�+.���ᮓ��Ӕ� ��>;���+�l�(s����K����Җ����佷�H܀ヺӿ��"�I����{ �Mo`�H��s�;OlHg)Q^��`˛�Z+�Z�
��m�35;���ylm��Y��UdNN/�r��`�s��|��j��$	s?C{��yD��&����ª�x�?ҙ��|>2��O!U��4��K�)����t�-�8�8C�|YvK����)'`�`<BX�QW$סf3��ٻ#�"N��PZ.̠sXI�=x����4]_�씕 l~"^��5i�ʷu;\5!y7�$?���G�pIN�������P��4�G�Gi'W��5F�P� ���#1�ɫ�Q�����Ё����\���������[�����qEw���Q\�V,�����h~�8-�R�n0���t��hk����N�	7�a�Q �	{o
:�K%GlaQl�F���P0J.�w+MIU�d�W�ƹz�f�=���L�S0E���''6�-c�s2
f��� ����q9�;x�kB�D�,�ˉ�r_Ey�t����,F�ƒ�C64/��b�+�r�Z��Z$��o��Dmp.dG\��-��p<e�3�W�F8��F��5&[�����Vb�|��W��L��7!��N��$Yiҽ�d���<�n&��lb�H���_h� ����4!Z�t0�cmR�����lЬa��b�%Qk����Z�V���/��X���_<����P��,u���P�*�/�?2:j~G׾���B�<\���.Rk�z>G�:J�%�\]���+1�s�zfSgn�g��>�e�v<.ox�9/ѵ�	�����pU�Z5�j�l�HivػM�!YKD�%�E*)�ѾV��\?F�v��u����R�:�ƀ��v����A.�LB�Ʌ"��a)Ά���p��jBr���}�:ٺ{�JE����D`c��Ztb`�TF� `�C��z��F��\sԴ�.��vw7-����l���.��u@�w�����/Pǽ���9�&���L��U�(�+���P߬V��_TƤd�zdGCֺ�e�]
�U{m��7m� �2���[=��2 �l
���|!��� Dv�Y��\���70�v+g���H���zU�ŎY@��������=��ϊ>Tᵇ�>����jtYE�����x�X��`�R�4~���14��2����c�z ��Y
?k�|��Zk���u����vE�2�YZ����^ڔ|왹	��_,$\�E��В�"�:y��/k��{"S(tn�̥V�K<�?~�QO�Vw.��ܠj�8�:����sk��xk�Gc u��GU���r��aH@�	ѽS��<߉/�욜i���G$�����ylO��B�fd^���BMv҂�f_���S1`�4H�qA���I���$�!�;l�w��|�w>��CvC�ʼHֳ�ĤP���3�~�`]��P�o�m}�P�<�;vd�.j�6j�l��8RdoH��p�%���m ̵�?k�gD��.�P1�c���k6[�7�(�n����L,K}�}E�M��0mg <��t"���G%���]�T����&q�*k3u:���ɡ^��SZ�
�F�o�����&��tb� O�ԫ�kQI7z����o�y�W_�si�X�vDk`ܘK�}�l;_;|���r�-�$�����=�J�Ձ��7}0�1���^���P��w7�;����fH)�[�9&b����_}���r�=����&�2A`N����-qK�3��ĖRV�Qh�t�
]XS��+IX�I��MqC+�󷋓<���s`J��|����Z#-	�"�jX��
 l����f�����L�b�i��[�ү�/�޶�,�iF�ݠ�;6�����ܤ�&^7{���b?o�m���i�;�����B������z�z
�6�P����&W�M�������j�-�7�d�v�n��fFN�?�$�#8ÁXIID�P�iHg�T5����{�fH���]&AN�5��D�e.�9�ƅX��3+��B�-�x�q���B���K�_w[2l:ͦ�6���1�a��ͬ���>dl;�E%�Y������Ո	��>X�D�4�M���䄄�̓��E�M�l�Xn.-�Ŝh�m�#)�E4�pY���Gnd|��z*x���@�2��l�A�,Fl����A�j7� ����8ͥ�|&��R��j�%8���C-�g*ȋp?�������#�	��=�J
V����Y���6�����Qv���̎�6^���_�0w����k}MZ^k!5�[ ��Y.�7�@��I ��a�C��}�
�wC�9Ԫ9�u3�FIc�n�Rz3�Ћ��SKdQU'��W^':2v��_�fF�f���5�`ω���us�+ji0e�027+'�>.�u�@C�l D� ( ����	�v��J$���5�2]Ua���(�ew^�$���x�_��Σ���i%!!睨�ݸt��B p�[z��sW��Kr4�U>�3\UEevt�>1m�ZH�bj��>�٥\�D�k�o_Do��&�Z����k��W���zUTϼV��&�k���Y2 Q@MXR+J���}���mm��.3�\�UR~�\k;_"�@Xc��äx���y�51��3�V��]��|��O���6O��`16MY�Zހ���LpOu��M�RY��,�.�(�NA����
\�wv���˃i`3���X��k6�h��� ��,��v�|X%|ʈ#��l��je$�����Q��'����t�p5 �R'o���bJE7�*0T��+��^���	�v�L�&�C�gL/�^���\�4@�_��!.[t���w�E�wj��(�%��gd	Q'�U������W�Ojº@;ݼԠ�)g�jV�05��.�g�l���,���{G$	�g�z�D��0�
��)�Zj�#�`�Po����r�
m!�U�8�P����J��(<Ho��τ�ƃ�qܛ��Ǥ�@֓&ɴTR�;&���?Ğ�Q����
�n�+�:V�nuu��p
t��B�Ԡ���ؓ�`�����GT.�(4��g�>����K�*�d�T��Ca| %�U%��4�e���ҟ���,b
�����[�:��U<z��p��mT�`���k�Md����%��i�-z�Oې��"-���Z��.O� ��@=��fU��{e�߱9ω�6v�t�I(���U��s��˘A�!$`D�+�ۡ��l3 �s
��QWx��)�W���ر�ɫ2��;��2�'�P+�e97��S����a�Ѻo���#����2}	(|ͣ��u��u��:i�k�J�S�~4s��$��&:��.��j��?����'B�ƣq �-E��A+^JO��q���7�ؘ�>U$JM������#�8�N�kg�F����8G���@5Cu��N�|�&�����p9�u��os �XKI�=��FT�!~�Y-E8��Uz5ᾧ���wah�V+~�M�V#1Β����?���n~�3A9�!"CEֿ�u/=��6�^��!��a����	��NDn}?8�̊R\�\� �B2��ᑉ����ͧ�_�XY�a��o&�FK�J�Bȫ�?'�or�V��`uO����M]v1(ť�zjl㞥[W#s� xu�wJ�i+���7��(@�'W�7�`����l�̝#�ܺ5T�z���Fd�O�t�(�Ձ6�yf��i���ӓ՛Y�����d�ˮ=���v��=/�g��ާ���1�(<���Yh���Ǐ=��DC��^:	�F�ZG����(v}L1�p�|�c叏J�) �=iV�d�8|�o�SNDɝ�@yanp�ғy+��7�����Uh����*�q���W[U�d��?=���݄�L~=<>@pIzr;@0��9��I���}I�NoM48�^��å+p2��Kn��=�h?�[���q�"RV�C��#���FW�/qHI<��n��9�x|qX���;���v�<��2?g�k����pRH��V� �Lyo8I����d@���!��"����-�Z�۰��� Hђ�5�u���P׽��HX��K��3��݉5E���3H��+m�����ѬL�)�c�d��t��:_L�����H����!�D�E'���z+�dp��Ԡ�w9x[���Bb�7c'b��:��%����_F[�*�yL�{�(R$w��R`찚kܓ[(�}�'�|�K}���=���U���w�hֈ����U� ��=F�(Y�ne���4��a{��"���ǥ�B>�X��+S���_@$F�6�{�c�ˆؐ�������;]ɘ�Υ��h�J�K+�j�h�"f���kL�3덇�'�q�l6��B�[#
��s�/
���.|&p�⹩*7�j��L��.S���_�P*� �g�	wh���sL���
:,90�d��� j�ۧ�5\%��{3��bk%h]xժگ)��7��.���2��k'+\>C���g�Ű#)��B�~vTI���4��LY��&dCe&1��
XzQY«PR}�L(�
[p�+����A�#�䏞l�`�S�N��]��Kω(9�
����ٺ4���<q�<Ǐ�F��.�s���?sk��O6͏'m����H�ќ��4G(Q�mry� �EI�[%�R�><UG S���q��9�8A����$�M�vs�IeRۓ5��#��57@�X��m��H��9�����?��NvŅ�R]��V�^FԖ"�+�;X'���{��¢n��{
��1����}�O�^Gl�
�Q7˲ͺ{Y�%���`A����j�]6�$ÿz�<r��O e�����E+�:/�Tӛ]��܋��3�.�zˎmm�Q'���c9�l��^�B,���˦68t�̐|�*��T����U�������P����� ~z�Ő/�hg�:��ɥ�ivl�A#�x�/x@}�eI����\|�����"��1���VJ[��j�L��&��`J�p��2��qt�^�D���v�R�Kҋ��x~�>w�{H��^|4�Eάv���Ӂ���Tx�^ޮ��s�YH��YS$���rQH����0�5r�Sf,��I#����I'+/��8��d.4���g�2#�-��]](�y�(� uʃ�_U���ֶ����v̫��{�Om΀~*��Ve��t���qݴF�zk~�T-68�!9^�LJd��������}O=�=ڴ����Hy :�Y�1���0p�I�gl����|AH�d�இ�b����v�����I���v��� �����t� {D�a���:�Bf���5-��1�9~+�F\�0=��=^��>7�B4�j�>r!�7ܢF��)���Zо�N��U�KB轭���oF #��h�H7P>g}�s���L�S�����i�3�}u���v9G�q#[݊����Cר:3��tV:�ș��MN�������9ڶ�+sCp４�di�'9����3 ��D�[�1�:���&�F�+�A���J��$lQ��j�A�o���L
��箬vw�C�by1���xjE����Ƞ(fm0��M�E �_l.���
Z7���|�CŌ���� �^�#��G�#q���������>	��G�u�L�m$�Ƞ���O��_�msw�α}����L���_�Tؚ+,�ݰ���[G���z2���>��p���x���F%R�=pzq�$����T�)�˧��k[�!�'0�����}���=�JI�u�s���o���K¤G
��q4�5�s,��[l�:��YZ���x",y��F E�Ȟ�*��~�N ��{���{j`�A��:��b~��/���N��{ߢ�@�B��4�A�l.\������t+���{��6�����Vv�x����Y ~ w�����E� ������s�`<�U�'���옶��g�3������8�.yA���6 t3�����W���&����$����}C�\�'H%;N-��B�&��1��)0�v�-�B4�%皴={�� �"�m�<Lnn'M�����x~��q#v�������,}w�X�<G� �?��v�\���(��;=,��)*ꗬ*K�V?����=R�����1o�"�k����.� �k���{�i|�k9}��t�%I�#��o����7[bP��Y�E��5��hf��X��O��x[N�%>�Ď�<m�:�,�3_�I��!,�\pkZ�oX���X`3H�b�b�XC�&nv�K�6 �u���'�'?N��'Dښ_8h�2�&*��Ce7wOd����5ҫ:��YK�4[�:�A6���::/Ƈ�@���v/.��|�v�6 ������� ��O�1R�ĮD����|�Իx���}x0������N'�2���a~I��pdx@fb�!�.�.��ل�Q R4� �bT[�����nj�Kn#���@���7BR1��Vs���P5�V�8��B��.�I��_a���Tm��P��l���� -@���Zꑌ߆c�Y=pL��Tk�����5��>h��B��Ԭ�BX�|MP̩�IӉ6��v* �B����7�rZ_�`l	�[�oKo	U�_"˴z;(��5NaXV!6��ɮ�9㬌�$�_�l0�A�C�����j������D�sV?�f��� ~�Wh���U'���G������Z���y�1����oBƲ4�!�|07Pq��L�z!�8"�;�UqO�`��t��*��[�KӯyB���E6K���䄎�V�t��<�3�+Lg �0�
Vu0@�^�����Ky���F����´l+�H~��2f��ÕqkKOt9���fU��#�r�c�����\ﰠ:G�G��
��P
�Od�r���L6=���R��ߢl�$��G	��.w�}؏v��m
h�����RWI�Q�°2ԓ���
�� 9��Q�u�L�1�"}Κ������J*��x}*ݑ�o�O{�/�����Onf��B����B�M6qx��[��2�EG�b�'�*�kmD_��Y��>���kd���ט8��5��U��)�.��s�������^6����uP���y�&�\�/�C�D���8�\�I@�.&{�^�j�Z��^1P���
��Q?x�ɾ�r��(O44�����K�o�cI�T��y��!Ԍ#�`�%�7��[����3�֌������v�!�\��Ѱ���|� *#�&��5ax�w�Ubڍj���+����,�/,�����t4ැ���[��M�Գާ`=��3���R�p\]P��k�`͐y����m�l��С_R@ԛ��J�@h"O�D�*����UQ�e;��@�dw׎%�.�B�|Ad��F�]�l(��e������e���1�{��Ik��
��B��ҏ�$ܺ�H�q=��~X���_Z����kkoVy&˂?����պQ�v�ы�[܎<��@�@�f��\�����WZy��kS�}n�����ط�e���C�{�U4h��(�b��� 8�ePzR�G߁N����_�q��j�. ��N�m�4!,�y=�@�z��w�O�6�s�A�����au�	�%"z<^�켅�I6�P�����\��X��/�����A�*_=0;�g䗍��Y��49��*�z����,lA�:�1�˂SiJ���f�y�����rޝ��]X����(�$*��A/׾�`9�WTBgQ����
�n��0t���"C��� b�����V�G0ע��ve�g�&���c��")�r0H�.�E`O�!z�cH����m�V}�xS4�l�\��P`�Y�G�J(]S�s~S$Gc+{��U��~�p�����z2�ˑ6d�P����8�R$�r��>(@�b;� Ȃ8�n:�-���r��&݊�_���Ű?f]�ۨ�ʘl:UḖ���j�����*�X~���+�͏VP�wB*�E@u����I-e����X}vs���L���3rN���X�}���@y���c�k� )���\D:���-_A�54�q�}��5N� o�	���lޅ�L�
k�5�.��l��Xh�����n�m,g�ު�����$�(Ӿ�A�w�h6��G����=�$�ܚ�r*�j��6k�Q64-3M���>#Ɨڵ��jN�Q<���-�P��sT�%p�MkI�B�؛��E�mL�(2�V%���C u����*�O8�?@w���+ї&��AD�.=Bf�����"��J@3+��f������3M&���K ����Šw��;y�]�8ѧ����Z88@Ǫ�<��'�����2�8�"�����gaB��mE�;���|ٮ�1���x�9xM
.,��������&�-��u�D�
Tx�Ds���[�?�;m0�[�	#T%��i�B�2� 0Z��7'ow��&�yū�5���w_j2�Z��X��5�I�~�^we�(\�(K#�/�H~s3ō͆3����A����`���}LD�{���>4�C8�T�.G�=�+��"�^���3�o/lR*6׿'�X�j��C�l�h��^�T��W�	r�a�3�Zms�\����m_E��Bz����5��aXt�We|t���(�:�ZE���I�'�>&��|��u�MVC{�� � t!�:^�˻
:Qn�d<�j������t�q��Yk��@�β݋H��Pen��L�n����V*P�AMA��Ⱦ�%��.)ZV$8 �I�\�kLusz:۸�҅"r�ëb9��9�!�;QV���񜡸�~_�Z�r�XC���лg����?h�j�8a����߁�3�ŕs\�ի�ga�UOgiT���F�P��v<�q���,H�d�{�F���J�����/���4� hKh�����c�1�<�:ugJ�hC������tz��&AqӜ<�q��g�� ���3�Լ�#��o���g�'��<���rL M3�����"Z`�!��%�YN���Zx��;�$�e}��E|Q����e@}�6o�\�njZP	��&�征W�2Rt��f��^?�'�G��bL:r/�e�N��K���O�n��L
fS�p>S7f��/M�8�3x��4)��m7���q�\ Uz����KUe�󰈒�\�$b��Hqz���08A�:�&��յ7�Ջ2�+9�(x��
�qB�h�QX�?�2��̲��PQE��>��M=���|��
���`x^�iԠu���}_x���-W�cS��ix7	Լ.�>���<��K��}_v#ieG��X���J�ġ��܉n���  ��Wj��� H�BnRs8S �mP��qa���t$�|��գ�~��3�rOw�H�o?����2�^CE�[*�v�A��6���ذ�ow���X��6��NVk�I��~4�*���M�h�J���ӗ�)���s�!񎠋�Ww�M�Ċ�g���߈�*�~�`)�����	TuIB����,��or4�C�O�$ny8�9s����D^�R�H��	s���r��Č`+Y�ʉ T���2�����kz��}C������ꔅL����+c�2q�F,D�v/�֌H|�����E�ѻR`yڎ�.BU޹9��}9���m��"��E0��ۻ�{�f��ؔ:S�Cb���ߏ	�9���� l����A�6���uK�n ��n53A����r�_4ߴ��*���t'��=�lvÍEd��H?>����ǟzXl�2��O��|z^4Zܬ*"!�M� ���-K�+(А_�U�H�^��z�T�U?����H�}���K�ð��G	�<&勑���4f
qi�Y�+��6<�� j��r� ��ᙫP�X�����^X�:���s���H�H�{K*�f����_x��>� ��n�{��bgݸ�����ۅ�n|.5�� lU��'��>��yL�b�X�|  �x�w�R����m4%l	TK�
����`���C�'���~�6�ȧW%w����Z	�D�$6p�s�E�
W�悃�(���?��$�1�{BĽ��5@r;���S@�"D{��Y)P��[�	,F �-?~���<0�T�5^8G���N=�U�E�.��u�<���s�IyS���d��[2�^~��ۆ���%�H�N��P�$m�þ*T�.k^���y��]�ʍc�(���lI'�bM�,���y���6��(:��;���g=��t(곴X��m�'Iq	Ki�&'9����h�{�G�N�`���C���̔�Q��mOTQ�o+#:����Q�����;�(̎[y��7X��]���*X���S�_ӴK��؅���ـ\#�U!�ݾ��#���B�Up�8���D4��$|��z����H`w�2�T�6��n�N~���*y{��U���K��E	|1(*�B,Е!!}�!}�B���^Qf����껉>�\�5�q
C��噀/v6dG�l��_��v�{��xͯ�%Jh�e�� � �^%�����/��2��7ב�ߵ4��~��i�7���V���xM��,��;]t,qD�2�0������`�С@
����R-�X�*��yH��	�^F���=��(�OM�Z'�%Or�gfRс�E�qqxm>�gָ�r�._M�槸� qU��q*�1ޚ�����?��|���|��a�<{��h��x�!�Ć��.�h\�ߛ,��6�W�q�2=�� ��L$SkF�6�/�[G`����J�	��⣺Qa�Ʈ�vW�I���������:� ���r����z /�h��=��W5>�pֹt��h��*��Zr4�<C���f�=B��z$=�nR.Y�k���\8�E��#��{J�u�d�S����Z���!Å�؄��y�'��ĔMTGG��L����	�map}rAe�p���^�osE����)���z�%����[v�9T����J���(��~V����l�6�N�^����@׭���~�n���o:~�G���:�W�O:�C+��v��d� ���n��ŗ́ ���u��G�R�p6E�LklE�i�תU�O�(%U� �W��A	2�{��UĞoŬ1�z��#d�X����RV�:5;��h���,0gE9�Jŏ�CGq��l׍Es�=�@�����fE1�q7�!$�+O��dڤ�3�~��D��=K'Mʼ#m_����� {]���ð�g�P����A���1��3">���e�f�D+��]5�Vj�������};��e/�������[� �+K-Q�'n���3`��t�U$D�o��)d�'L��`U�x�W�׈�bYW�w0�����Bhz�|&WQ7T:~���5��b�!]?���ɬ/I
�4��
0?{��D��v2����Aw1�:��� ��S�B���(����%��b���g4������7��� �@�$�3֓��^���T|��՚O�+�m8��:��I�B�i-��ƍ+��~j�(ˬ���р�D��������������q��Z��L��o0+�a�4���/L["c`���ɋaѽ0Y_@���X�byM#��4$���i�_�}��Y��h.�K�������O��3Z���m��\�]$��7g(��#�#�6�Z\qEY���4���k_TMQ(/�o��{���xe�eu�zU�ڇ=���"M�@e��>�F#�����Щ�\�fdL�V��Ϭ(���g)�D(^�l�R#�M���@c�h��3z�2���=�η4���q�4��gFr��X��6e@Ձ��nX�I���̢R�/a?FP�YL�Z���Iި�B5���Ūɥ2�m��L��oWlђ�n�ܺ�+��*���ի��hPR�D���7�Bt�����^Z����9c��/���0ߢ���e��߾�5�,۱�F��+�� �D�)��A�1=V�rr-	2!A�]��kR=���c������I�dM���P?��:��5�I�pcm������ǘ���I�8�)�oG�
��v`�v�qΎw߁�WI�)���1���~g~z�p۾��u�bF������l�9��q�R~��3X�-�^�>��c�#KB�K�v�<������b:�Cz�t��S�
4�X:Nk&�3O��@��Ui7)��/�o��-�t-��@e�CQ����'��Z�g���OU�b�wt��-���&\�P���e?����W�+2:���>�j�B�l�l֤��i���&d�|��Rj�d�c�f��� Q�-�Gnk�� ل��n�n7�	�O��a��1n�H���JK�`1ZI��$����S��5lQ2�U���i쿗{������RĪF5tP��T�?��v���p[w6E���KN�/��G���N�q#$v��:d;�Y0�Q�;l�s8�u�#���QUUB@���Tz�8W�<B�r������	p�h&�y)J1�Cn5ϭ��G㰻kliF�VB�4�vXwNYg5�-��_ѭ3�9[T�%����:��A2!~��ҢmzI� 1�qY�=��?l�����vӣ,ߣڼ���E1a�+d�[d�	@�����	F�L�ܗ��=g�1}���Y��8�|��bФ�Z��	�x�G� D~hf1!sV1f�ȣ�1O�����FU��� �b�>��c,��9�]�h]>c8�YYf�`@ �`[��(`/#�� ���RChRoǒ=C�%�v���q��A��BT4c�"h%��:B�OKe6���m����l��<؇��f/�T�K�����<<ŀ���7�!�\ŅB2�sI�d���������I2����u��Y��(�Q��b�`�W%%�0>�J>ɢIl9d�{P�]�c�J�����:V�H�*�qV������ĄwI!O4od�� `�5��̎u\�e��`Jr�q�F=���e1 75�`|>��)�ڴf�n4���Nx����JR�팍柆� �\
o�GQBL�����$�{@����Se�:��C�E��R�g��n�b=B]��;x��	��B�wm\g; -ٗ"ݪ�,�8'�t���At���鈾x��g,e��/�8�7�u��T`�$ʝ��vYd,�iҐ�;ê+?AY5��vlr5� -��7��p�I��9�:��'�E�2ȸ. c������yr�u<i�.]��o[�N��-g �����c��8���Q��[[G0E���r@�@��czPޅ�x��Q�L�o(@�����Y��~ ����s���bl�k즲e�m���|mX��5ЬR�Z�E�ǲ:+\	���K�ZG�����}I�0�iT�F��B�`F�"�VW�����|�ܡ��@8:}ȶ���I��k�o��3�����/<#�Td��� ��1t��_�C���Ƹ���׮��'�	j�P�S��Y��Y^��2��v�7�@ܛ~!���A.�����r|�ū�	�~TBtR�%rk�s��t��͡�u�_,Ɵٰ��͏<e��f�_p	�tͺ�>����@x���¸�O!�ZTX��]m�>?몀-��V�6�\�|�{&�b��?�3�L�4����?�YA�odr�y^�G�?L�~S+��^�T
�yC9>7�m��!~�|��j�{f �obG.���F^�׬#[c5�*�����J����QB,��²v��eU���;��x<ҏ?���Q��{c�5~��3���N����9�-CB['uwt�����_3/*=M�m�G���kMqF���	'Q��<9$K6v-�~~�j����y~�F�pR�E�ov9S�h�^̓�3-b;
�_=���r���U"�w�%f��D��ϱ᷒��<�@!��q��LBŧ�|� ����d鏽��e�����Y��`=pP�8d�By�م���mnN��7�����*L�ĸ�ߒ����#x����E�Kh�e��Êˍ��������4���T�t��R��x(�:qH�"ta�'�4[��&�oGo�1n�n.d���UO� �$PZm��*��MY$�\���7Y�,9M�>�C8V�������F�H&�����I���g�Ɨ����Q�^-��Ay,��&sXDQ�U4�%ma�m0W��סMm�h�G�^����o��y@�=�r^�w�FCZ�����_����_m��Y��)�<i���orZ��(.R��d+���i��A�ݷ��k���[{����<�!ah���`�>��������4���������|��ji���^�7�i�J�\�G�D-@��G��C� ��_�4�j����d��Q���G�����T�c.���#ͮ[��D6.a��Wi�Ykش�8v��q�\�M�Y�<��~$B�/�Kc��mA�)��x�Gv�&��о�� H�9�0�O�;�����M�����>�N����;���@�8:���)ДT�$Mg3���ޖ>�(r��<wǖZ�&oz���0���f�r�Ok%X�����3<�]FB��厑&A��m�籲6b%���sȉ*ǽ'����'�y�?bھB�'��*bF\&���DH��/k��l-H�F�����Z��;�D�AVR�Tܥ�>�No��cP�����4�.�/�@��-���!�nCT�3Zg�c]��P�<���1��gZ�Z�� ���V�ȯ���[�D��[�Z�~�vе��/���3���-�Y�E,��ڠ����OJ�Xg ���OO:��XDo�����a����L�9f^)X���,��P!|}����Z��Idhk$��/+SH$�R9���7G�-r)X������0�9�M���ב9�p��[�b"l*�\����x7/B��߇�2��k��˱FX/Pro��^s��b�@��:?����\��B= �0i��z@_F#cXn�u������P���Ͻ;�6���m2z�w9Qdj�=nE|�i��N�m&G�᭮��K��*5�/7�>p�x4]; #Y4��H<�n�AK�*hh�'���
��kckwl��B	�9�M���s�3)A~���Η�0�VY>���5̢4�w�;�;�mB��G?XŽ ���h�h�̀w<1_�
~�����(0e9��x�=�IY��B���Iњ����o���
[̄��ӝw`8�dI��]�a�m�q�'���Uɶ� �gaz��^���,���7�w�6d�[m��D�lZ�@Nd�Pb�z����l�v��Q=.�))�~�+a�mϯl���,4���C��s�$1m����@�OӲ�JZ!z��p�%L��ř���u�^�c ��Ȑ=g�5Y�/P&�)J�H��%��ה�q/���$��xj��ۡ��uR���X��q��F$���2�f���a��i1��`���@����l�[�42����mxyWF�i��i�Ҵ�YcB���#O�e8$�pyS았�jΘw�^�!(�����(��5H��QϿ7ί����1
��P���5}��8��{[�	4�y#�nQ#���;' s������"�ǜQvw�}x=��^D�8:ڽ�ޯSy"�Zֿ�_��+�ݭi:{��A�Yr>K�6bq;�Z��
i�q+C�п��Ҝ9���sTrv�����D'%GۿNoB��0C�υW��,G�6�S�pH-���͉�h5%�?���O���5j������Pxk�� +��#�>�)x�̷�N���Q\+}�����@.yD��܋h�(�i�#Vt&I?����}&q��8�*�K�F�?`ۑl	��e�|�0���^��R��=Vy�=T�xΞ�ܘmUz�����/;�����<L���1�������SB;7I�D�M"WRMalQ�^��՝���r�t}#�t 6��9$�]������J���L��<6�A~9'���֎��"}�?�}Q%6�)D0�ï��嘆���Q�٥$"��䂲xzgE���ޜ�@�oS������تu��$�����k�b��|�+@����nC�D��]�����ܙ��>��6<ER_��;hȍx=�,�ּlW킺���h`��Y��I[l�;и�^�Ε�9��K�9U��D�f��$ܓx������L�$cO�x\OJ
�<wWh1��C�!�_��r�\t!����Oԏ���ܱ���z�i�Y�b��2T�s�B��3�%tI8���u��,�e_z�;��5/8�<��.ލ�!|�O�+�����w }�mc�cOں�h�����C�HK�P�%#-�ke?�]�A�l��w����_ZPc�t�q���|����	��	y0G�ܨ Lېo�u��0�'w��.�����#�k���M�-����Y���<w��}+�Ӓ��s�z��~jP{��y���?8BIf@A�lkyċb��o��]^��7����2,� �����V	+a�ӌp\��#o�=��?�� Փx8�J�V��yӚ��a�0S�ܕO���!|���0¹�clя�O(��ꦮ.01�10���a�3q�RM�ut�0Gh�iP}j���U��L@g܈T�}D�:�'�y�d�9��P�����#���2Q_���Rw�R��Δ��g�s�-T����z����D�?���(�#j�äV��ك`�|y��=��	�L)�l��B9=
Щf fp���2���G���O#�:���.�}���ç�#�Ć?6u��2,���SL����h
-��됕9~S# )�[~G��'fGijQ��� c�7:#�1��M�29\ek��⫯�ĥ��&��e/����P�+̉g��É���RM��w>m���Iv�x��uO���1�b�+%�/�J ?��w9��	ni�`���oϴ
�c�� �?|b#9Qs��e�\��\n�6���	�1��	�3�O�Nc�0S�D��?������!� 	O��U��J�>��m,�⾮i>o�cA�������%�R$ϼ��b�g"e��{�w�>���U�S#�������(W���W���Wb��2`�aKY����Yy�>�a0�֤�F�p!6]��+�!;�#	�[�p�z�W�V�����6pSk�?A�j��`��\�S��r!�H=�i���*����K�Kdku��%�p�Eʞ��aU�n �E�`�y���d��s�ӂ�%���'hN���A�9ҮZ)9k�s:�"�N:f$�kd�b�G��Ǵiu��UF=�>�-���=��4=�Z�7�$���^24E�������<p�d�"u� T�Y��@�&V��'.	y�ν�c�?�k�#H��B��+.��$�P�>����.}�H����l�f�9�Z���������j��sn+��ޟ�@�js! (&rݴIh�>�����P0��F�?���I:�<������(tw�D sJ;�y�0��������J��g�ZG�����^�z��QB�����7�Ij8��]��7	����v$�T'x�W ���9,r�T��l�
�u�-�$��l�t���l��6~���� Z��h��l0|��I���ĭ�ь��	NG��Ȭ4��h�,��L4f&�or����O�/��.��W� 4��>U/9��{,U�A��și�੺�Fж���J�*"O�>,K������N���q7WuobD9��3����+yk9ݼ�I��0�['�8�\?r�	��t0������9��=<��63f"���nv�H�_X�sw�6И����.B��'ڥy��6�T���L}|kz��Zʜk�|aV79�)I�3�s�9+��$	�r��׆�Rx��?!� ɱ��Yd���ܑ������V�����?c�]�6����(�����P����,/��Ǒ�9K%,�d���t����L��DJ0KZi�s��y �!��dB��۸��V�dg����]�:��(S#����r2�1�X�3��Փ��b���8��-U�1G�w�Ѣfv�0Z�ۚ��ʆ�
#�
P��6����s%�@�����K%��#<�\�*s������������*`�p�Ym=�����V�B��%���p��Z�D��@Hg% @eK��I�O�M
�(��(��ƃ^�-�'!#y*�]p�'�R|T�F�t���o���N�D�@7��^(�J��a��6���鈛�V:�X�F{�æ���a�����2:�Ci�22`�d4X�������t9ݧ�O�ny?XQ8"�W����x�P����y1�v���l��
��=x����v����@�����q;���"YLؚ&����q�6J�uT��u�F$k���@kd̇���R����][;䔩(�q@����]�5u/��( �XNo������
KS�S��*���
��";���̍�ɠ�=���NbWέ�O§_ �~������T|<�c�����"����]Z��\i���P���M�yY8�ݟ!�������hԄiBߗ���x�lP�f?I��*T~$k�6b�y�o��<ڣ���!���:x �g��;�9��G�������������>P�M	�7��oN��$-���|��l��ώ:{\x���k������U�c�T�fV��C�?螰�?�'��&{��im>�a9j�*S�j`,x2�	���l]�H�`����S{m�{$�R�b1.Y�;�-���{�c�W.n2p�> %<r��`O?���4T�ҏ�:ր�'�߀B�/rr��&�Va�{��U5%_�����5����އJ\��v�;��'0/ڊ���[����[�.���W�p�c�%�N����RA,���v�⩊��o��`�r�݃���T�zH���-�>�aY�BI�k
K�Z����t��V���.�g�F��D�5�����r��]m�!����է�߫�u�a'O�>�����S0��{���|�K���O�
��L��}�arȔ}z\��Q���������!���n�}?�k5��������-SF:��եT�%���'���!s[ZBb^�׽r2�bP��&��L*�&��+fD��C�XXWcV}�O��������8s0�T��g�o�C�u@���f��،��ظ� �y˼�x'��;bތ�&�����(�ngNЧ�O��V'E�g���K�Ԕh�a����]ߵ��B6��I�X5�Yu�h󭃺�b�T���'m��Ŋ#E�Kq�=f�ǜQ�|��6-b�7�I�@,!㜁�����[� �gl#�K�M[�Um�8�z0��h4�ʔ�Bin�=	P\���f���|X�N��CI(�P� ���H�U���,� ��3�([Dl2���h�쌥G��|{p,��z܏����|��B'$�Ne�l���J�$G�U�r�j,%΅���^���`&����X�#�O� �\ v��XRR��
�8�-��V�j�o�����}Pr�̾�i�X�z��ۯ��i��U�ª�#���K�Wl[O����؎c����z�!��z�UH����1�p�H�#���J�|S�\4!��ߡ/�������`�l��;�(��u�м����;��M�!@.��U#��O��2\�8ai#������0�VEW���_\v��9�U
� �H��p��������oi���Pr��k?x9��E��?�=�(ٕ0b�l�%�'���h��T�|,*)��{����^#� 5��_��zz����yvy�C-�H�Ch�2�E��������u�b��+E.��FOw��̢���ڏ� �ސ>�ЬY�ᮬ�s��[�1ۍi%�\�􍥾	㚬*oS�0Ùv��7nsT�N`=y��z�L=�>�99k COX2]�^�.}-�*�_T��B?Cޮ��w�/p������)���=��z�B~D_pC2#�	���c�$0 R0	�t�?�/*p�H9�ۛpg�m0�WÊ��'�7���~Ԯ�z�*a�팿Y���E)���Ԃ��tL�<��̉۶$���b���ԧP��Q�d{'݇z-�Cz��§M9���֘�ה�)�=�KNP�k��}�	*2)tT"'��WF�[�·U������L=���
;���r����J���oRYr��s)���p�P~��i�/�ڱL�w=�!8�Ѫr
�&��d��S�t�(���o=r�HET8����%Y�Z ��U��W^8P��٠/(��B&�{S8��tu��ze�V�u���{�0?C$���_^9�6	+�a�F��{#��T�!
G����5��Z�&���3I���j?d��O}?�o��i�f"�BA!o��f֞�7��e����"R���L�#�t�uɇP�J�S7����}�صǀ]wB�W#���+��0{�D��}_@w�h(�����hrZ�|��r&�a� bS��e,}2��U�0�"D-j���lE�c�\��Zcv? ���v>KH�EM� ��@�K\fdPf�#} ��c���0��v0�:6Ӛ@>�~>4�P[��9ܡ$_��M�q��`S�D�V���,?���j��Ғ�\��o?�S�&u5���L�_hS^�����7����X*��g{4hO� qη(�������G�˼{��/��K? ��2���'��47^-זּm��$K�r����uWO�'?\�d�qc�h�@��ܳ(�m��TKBg� Ed��5\�zYFg��v���/9j*/�9���y?$%ľ**R	o��3 bUmd��'�����2������N6��A�j�L��;kC�S����z��~�����J�ax[cz\�XJd�[;|��2Q�u�&P�i'��B�l���ŬϘ^/�j!����n҅x�f�r�߽�u����*\8�~�ZHe�QI.�e�/���~G�*��=����.a�q�ItAy7	� �Q�X�6�PU�onO+z�!Q���-�_=��8�Kv�pr5��f���#Ր+U:A
�\���~���2ʮ�/I�R@W�Z���va~�6	]�^�=�jiF�mS|R�Z��;X��0�]hT��7}�Pȵ�A��s��Mz�<!9�L�V��C�f��m�A����_*��J�+�����v',��=J��۝� /_��B��1�!mĝ�N���z��.E�<�E���O��Ͷ�aT[�>R�*��W@���i"ξe�������N�ަB�~�^1���} T��w���a�*�_U��Fjf\�M���do���,Ξ�8g˴�{ҳHpFJ��D�������ŷ�D.��e������)����tIq�z��j[�T�����I�:����C�$���:���L�S�!�f�b�+�T;�Q���p�o� �=s�<J��Nݡ��L���}����_u��#�ݢ���J_^WH`���9'�8P����q� j>[M����[SFz���i7M��r�����Wߔ�#�8G�������G�h?Y�$lڋ%m�@k���AT�Rt��t#}-�%e���&�j���u�zѵo�VqA0)JU�)�ǘ�'<V`�*+��'I֐�qS��t���4;��h�rC������W���
�ZJo�/�.Zw\���c���m��ggX.�=�أ�*��R]��Q���<���
ތ�E��SC�p����}��/��s�86�����}�'��h9������
3������QT��h1��I��U6:j�js"
�]��=A�w]h��1/@W:폿�<jC���Z�(��o�����Uo~WZ�wp7�W]"�X-��80`PQ�{��2���� (\�Cz�4�@���O�Hc��8�F�=@�K=v-2ΐ}�Lz��',펼Ve��lU�5�V9���<=�
��V�����Z#�&���ω���6ԅ��?��>#�j�4��Y������K2�_��q���wX}"�1)�c�4ɉ��4G��Fo,�X�/N������U�1��6�<)wRJ��q�������a˱��\7�o����5��m��.���3��"��Z���,�lG�
�ߣ}�O��,�U'j�L�)��Z���܀�É5YYl��}���oP��(y��Gt�H'� *U�d��<�Y	E7��w^�
S���B?��%r���UW��4sRi`5�[8��ҮV##DȠpD;�H#���0LL�a��hw��9��Sq�gW0󗭐Q�=KbI����r�+�\¡ܞ�@ߎ/g|:�����x�Uj����l;3��
g�����?B�G��0�^g�/p������5�1�P�	9+̑�:�U�'�q�Ew�  ��}C[U��_-d��qX�-��(U�xzW,�O;/���dtZ��A�a�ǵTBt謀���T�yp��~D?\��z\�]YC��Jz\��!MT`��#.2j7�R���(�0Uu3p�L�ӱ5j�]^�^!^���7`��x[j�`�%Z�Ҧ2���pa��B�-X��p	@X�*�Sžؗ%�~��ӓ�&yA��EP�����:}җ�Ë~$B��|D]t5U�_ͮ���)#���/�O[�P(�]�Q_ŵ �0�[va�	Z1�m�2�f\[a�Y��հ�r=��[��-����t&lF�&���,��]�2�F�P�������T����4���&B��ͩ�h�$%#(�m��[)�+��j���7�>�t����|}�.��jB�kxA�I��X��w�BxzA\x�mH���Vs�Ǣ0O���~ѭ����uv;���a*S���l5@��d�	�#,V6Q���4c����9�&��
�P�8��HQ�P�bUO�'"ز��D�;!��� Ownb)X���X��*6wU���G=��c}jm��}	�;�V$Ml��q@�\uT)�� � ��� T.��;h�"H��YQޚ�*�nlݾH�,&х�x�D���F�������5)��E�+�5L���5��P-�Q�zG��������o�D\��z����"V���d	���e��>��������M��1��H�����-�EW/������~�k.�Ј�O��(�$e#���n�%�;��[Ψ��1��tō2�p��9%v5�����n|�Y�9iS2�o���ؑ��s�3�@	���r��x����Lu�C0��e���f��͑�8	��Y�pq
V��k ��0Rq
m��䄄}WD�g���� ��w��2�:����k�ߵ!j���>�£��.Vf���R��C���� [��#>�����D�M�Y<��,Q�6*᠘�X6'��u��_�Վ��i�/({�tڢ0=Of8���5��weKG%u�j*��H�,��J\�z�U�{i�a؋y���E}/9��f������z>�Р?��ʫ6�v��\� ���i�Ƽ�Gu��@
�=$�s��i�����Y�uZ�����%d��0��DEGq�r�+�uάH|RTZu
iC|O�"ݿ<��,(Xw�0~g��j_۱x�MBbG�����_�!�X�@;#��4��ό��_��	��௷�eЭ����Q��{������5|12��������YGA!Q�p�7��R�h��e�/m����Q��n���6���?�=�`Qm�8"(��J�8�д����g�:L�I��C���/�@d�_l����2�D~j�G��c�^� 猅�Ct�n�!��?j�JMtx���v�E"�:FDfR�Q?V���p� ���	�amL�@{vuUOp/�UH#l='��_��,_J�r�zӄ�H�T�V+˭���Z5;u¸(��m�Ѧh��}H���]���E��S��u�&$���W�HL�������O2���)a�s���Q���(K�jp�u�	|�G�,�e� u*��m����P<���p�,�,-����!��j�:�<,-Z	�N`h�'��g�}CD��On޷l��I���I������d +�������R�`����M�5�!�(�U���po��_�L�b��	�Ja ���E�n��`S��E��_��ʾwJ���_ǕQ�kQ����W�uo�gh�έ�H�>G�ʉ`���Ҏ����^�鈂�����1Թ
w�j	Ei ��(�� ��^	�yaa{�t���O�*��B�^�@t��Ԛ���!�M����Ϣ�L5�h��پ��gzވ�����9&I ��Y��;k��YJ�2»Id��A�lō�۔���u�hB�FG�E*�#c��+���i*��o�!��n�iʘ������
�b.���Ȭ��Jj(�/-p�7�z�5�_uQ\zǮ�m��׷�|�ĩ����;�r�פ��6��܄��!���#���!;$�SU調���;eSK?�`�:#J-X���L�Rb�l��TUDl�V8����>�3��a�Ir�m��Gl@��xi@f�K�ѡD�}�Ӆ{���yU]�Bҩ�Q�v�zxn�;)|�ʱ/Z[��)m�n!�	6�V�
e���C/�	��7�$;߮�GQa\�o��?��t��u��.o�b��ʿP۪��r»L��#6�>�$��B�X�G��bۯ���_<)�Mi�&�y�x����<wL��G9���b�nJ|[j� w,�C"��t���SL3L�	�_,�r��JG�,��y٠��r�	�К�#�GCp��Ū۪�(�藜K��~SwX�kow�%a���4$	H@�Ur O�2�s�n�5�,���pɵj���Y���&�4�Ԧ�]����"9����\������V'\1�$`��\�C�}z��@V�:��tB5)8/=�Y֡��1� Ta�"���[)��˽`3鈖�]B4:`�E!ch�xs��i�?U1`w�<|�������@٥,��b�[uq�u��ԠJ���Cʃ5��Z~�&�-����.�S����铴t[��)� ʷ�Ԃí�?�q~fôN��"���	@ܑ�fzޒ�?�~�/�޼�f�O����!̛x�$��S*�4��Y����d���کGd�7��[E����hG�@�姮|0<�Q���VA�k6�N��V$����N����|�pL��]N]�aO�%*�Cl��Xz6�`�]\-���l7OK�u��3�7Ԭ_X�(OTH�D�ݢ;��Ê�F+/����@N#��C����9i�A�����\.�O�~[L��>�X�^NC7��@�W���.U��4�`�I|LO?���A��p#�!�P�u	���;Z�A���_m"p���F��}���!�c�Z�d-�r�[�rQ\����hP�*�z�<LPў9J�a�WC:Fx���>7y�䤫���Ou�aӕ�d� ��ފ�m�y����C����Gn'Y��0?�\W��b�\���F�i��Ш�=��l\7�	P�u+��c�k@�aLT@1�f� ���~����,{77!�����H���vW/��3σ�f�V��~ݦ�^�Ƕ�M�ݶvi��[{Q8X�	����1Q��<P-7����T���`
�~(oe0���%����u����]G�\i�v���IБ�5چ�n���}&��,K;p̠'�\�[�/֪w8�� ��_\�Q�m��3�':�'5	��z2C�.V�rzk�ٰ�*#��K���z��q�.W�TR]y��B����.��L�f�����d�tۗ�
	3��D���|��f�'J�ܟ�d��ʌ*�q�f/P+e%.A"&��l�l2�C��_f43����,|��*��+�3<t�|";�'��.��RoQ5���~p�b����PnV,�'(��꒧�˱�Q�@@�Zܫ��M�� ��SyTI4�Q��6��!�����A��N��y�`��3'8�/Q����u�S����1*S��/-�QF��(����N ����*��J��
���֢aH�������ኊ�|Ae�o�ev��{}ߠ1��H��Q��3uo�?N��F�R�w�v��b^�����=D| xw)�[�[�ZߴLe:��(�d�����(����U�,)�&����,=j�02ч�s�d�;�>�5���QA������i�=)�� �w;��Փ��e����JH�ƯE���q�	��0&�gC��a99�����?��㮌_�:��+J�����嫕W5�` �I���a���	�k�lj�"�ZX<�	L!��&��9Y�
�F?�l��}���5��0v\σ��	���t
0L.Ī�%!�����~޾D��w.XU��=7X[ �H��P/׶�7!@�;r@.aW�2	1xӀ��ʴ�a�b6i~~jGDO�,��o'�7���=���n�B�Vb�z����O�q�3���^^�NyT~��A���{u͵sr)�����qEm�2���j}྆�|#�Ԝ�p�Ot�0
����QD�]J�����������
�3ך��������og��$�G��5fuaOax?n��"�I��1j�
�wd�}� $W��YO^~��L��G�^>�?���y�d -^�?Wj}�Rޅ�{��ԼƢ{� ^sPIZO�Pt��[��ls��Cgg����>�T�����s��}cz?!���ە�S&��J�x����( ��$C9b��?�(�� �Y֗��m�-Nm%a��z�Z$�ͧ������;T�ɍ����k(����Q�R�4��#i���䳞u�+Ytq�!�Ƈ)�\���ȏ�5Z�l�9�_F���pu��w�=�d��]՗-�N FS�.1����َ䑁;	F�ћ7T,�U��}�IȻ���ӾBqnК\�[����BI% ���f����>:E�'�g�h��3��bU9�I�ܪ���k��n����#�F)!����ܤ�h8�h��>�U@���츈$�4�a��� Fi��臞��|�ܓ�g�C}F��n�eptj�k��T���������뚾`[w�w����q%T�-fb��1��$ev���,OoV�PZ�S�'��˗B�sF�YS�����0f(IJ4�p۠#������u�&�~SvXY��Gu�����3;�ޡ��1�J
Ybe��Yg�<�t�^�������5��ڬ{ί�R(�;L�e%Y�'Sے�����:�� }<\O�ż>�Z�.��f]�kߣ��	���`C3
-���:O�Z��
��C��$�K>بb���
��am��
��߼P�V���:���lpP;�0ދ�M(Ã���%�i!v�fӃ*)���8'$>M��Sn�k��0������P�W�	P12өyA+J���y�|Gg��p��},q�����mI!
�Q�:�Q3�y�֜=�V�b�t!�I_̍ㆷ�s3$��pb�&���0M2>Š� P5�Yco��w�m�!P�A���~�~N�W��W�{�-�w�:���7�W��D�me�h ����7���G�����|�36I��j�]ý�9���A�2:��߿,�Y�_��"���tA9�g  '��t�8���S{f��&�w��qe�,V�~���o�|L�tT�`5����k�i�_z���:�7��[[ �1i�1�{���z0zq���I�Pk���wt��s������帶�U\F	��ֳ���1xٔ�տ{g'~mhT�{- pN~��vO럛~\�����HA:@0q��,�3w=ɤ	/.�_��j��Щ��f��<d��"3,���A�#0��\n�\X�64'�q�"�f���0xC�'?1No���#��(�&��5:�q�%	�{��W,����[����1����8:sDٜ�������B�l�{�kA��bT��Fhnzi��(l�������P	���t�:��H����Ef��ѓ߮�4(z�T<�SJ�<0Ļ��P��7�Qb�\�{���E��ު�K���봜ä�������?\=��۫=������^�U���G]��U���kn��؏P��{��)��b�A��M]?מ:Ň���d�q�ǐ5o3��G�B�fM��^�&��1w�U���Y�X	!%��#�S�����p��+k����4�Y�d�e�B���Z�)K��g3h=�
���!dҝl�$��t�fDع]���\�9a8�tX�w��r�pS��C��>x������n�hd)V��n�+0C�s�
M�ig;�/3� ci�lK�)�(��Ц�Z���PÛ��mrZ,�醵���ݍcH2�	H^�f���T)Е[��6�?s�nv�&d'=!�s2[�
D�h������e�댊sڗ,�F:�xܤ����39��s����2vށ���)��D��ݻ�΢��m�)h�����Ήᵐ~hQs�M�OW��;�#Ƥ��Z>�P����A��܀�樓�I,��~)Y`y<�9�K����ʝ`�Q%�ɢG��E�K�=�)l�P�<8\G�Y���½/�����-*�R�	��VB+iݞ��>��>�^�(ˑ7Ys�r4,��kr��L�7F��>���JkV<m���TJ"�6kw��&�Z��J�aw�' �vf����ӳ�#V4��>ߩn)���TC�lתLx~}�ě{Ϣ]{�:��/{��Ҩ��*�}i%�R�<}}�{2Cr��nV9<�h��^����_��
a�zG�,���l���@ȅ�W��%�x�ZsC�f˔�[ c2�ǎ��C��'j;��H��,j���#��t��R
��CѸ�4�G���b9j�,`�1�C���xBƷ�#�E��5����%�2ƊK�.��"=�~���k��r�$�0@��2a����a)���Ţ�r%X��:�G��DQc���_�m%1��GU]�G��Lr��X��=(��Ao�orX��J��Zٓ�9	U0Rx��+0ͣ/��S ��ؙ��kEG���s������Ҙw}�0�)���Z�<�X�
o�Swq���s�u��{g��Q�]���qcjo��zʑ��A�nDmf;�9����tM)��g���T*jQ���P��^/�2�2�yQkQ���(�ok�>�Υğ�m)�W��1n�O3$��tx���`�@�ɏ���)��a�����c���+'Ore~�H��;�27ZH?a�'Q�hb�,>Z"�Iok��¼����]��*�`����D�g����-�Ƹ�Gn*L�/�D��b��$J@5��
���Ea}
 vk�1'Uϻ���E�N�bt
������%�z�
7�Ӹ�H'�p�ο��k�҆� ��%sPIC]+�)5�lAF��I!��Aʬ�Q���h��C��ː�|��M�lP�g޹�c>˒ѐ��7킙!8
	AB���9����j}#�1�KF]�cWH<%ַ�l���:i�Ж h'��!+(�%����M��y�JI^�nQۍ�i܋�Aʪ"5�A���!�� 7J/��AN�~
�6��V�-�c=S��)��n�.�L��l�
�ˢ�Cy�v�f��c%ZY�3�8)���3�ƯXX������W)�ABؔP㗅�������ߴ�O�0�9�;�nx�����sC�M1)�J)Q	��N�s�.\h�~�^F/���HE�Y�+�S��8��"3�����U�o�����Z�&���=%-T7��,d��VXd���ݑ��f�n)w'Cߡ9��,��f;��#|0Ir� o��C�U����B��9������S�u�����4�0눥D:�U#�S�T����骲����uy�I�����3��� a��$�H���4�j�0d�T?!��{	����p
����7^��UUɶ&sr�c����k���1����Õ��j H�F(�7k�%�T�R}�䱫n�����i�~pno�����ʴfʙ����P��t����/ۈ�SRh�5��
����r���"��;d�%�_��4ln՝��$�r�9y,�m�ͥ��& ;��[&���� ���wΐ;�{a��I�z;��	��K�6զd�a����u+1D�)�pv���#N��0L���*Q���.��d�0��L� 1�?�V2J3\v��ս�%;>ȇM�Y߹����������R}-�D���xL���:�zbjV�Wک�f**��]E��]U��ĜH`w',K�d%^ ?S |3��!3���[}�4$���2�4n�[�um��E�v���m��B�����@�%�f�B�)(��E[��U��U�<dΠ�Q�x#�8S"��bh�W��������������:b�.������������_�c#��_{�b���!�W�M��3�V���z@��wTJ�*4t��BH���W����{7�cE[+�}7蝭���)����aB��3�g�HiI3ɕ(�?����B�An[F[��#s��!6��@��Xm�y{����T�g�y��� ���S7�;�V�/�*���w|	=;=i�w�W��ԍx��rY��5̪��?���d.�	0�igѠ��*#S*Rj�ʷ�0h4<��c`(�ȿ�
�B)_�y�Y?{5��2�K���5��
)��k�܅)�t	n"|�S?�e�
�Ҵ]���x��ـ�Uێb6��7�f�����]����Ev(�h3*HȓP�tA@���	̲��=��&m��Y6�C�A��zX��y>ъ��R���ئ�C_�W������M�������:l���݊m P8�D����ݔ���-�
Y{`_��NU���N~)�:U����)0RH(��{z��UnPz B��١_�>�y�����j�m��u���+h��x����~.e��$����z�$�W	���v%��/:s�;M��x�oR�آ'���l'[�01@��ß���C�V�j�e=�u��@��*|]w��kY )��:Gt��HJ���R������z%���̥~(�?�{҃��FI)�$0����@�^�h�N(�)�޹��a.����P��-�[��dI`薙�@��?c���a;zv�>z���CbO�G�����qzm��b����k`0�~��.�$z�#&%�(Ғ�H�ڽ�Β�-SW:�~�R�ӵ�?�3����_Z�[�¹$����H2�Lu�3Kb�ͤ
�[�?6cۇR���:�G�7�xx�4��Ƹw�_���@���C�u(���LL&#V9-����4���ݽ^e@��
��_��Y�v���1B�Tk~�!=�����I=3���eZ5��&���"��F0.����7�Q�ID�}��]8�I0�o��'o=��7�G;�.���3n��J�߳r�ƃ^�k����%YyN ɂI\��5��S@�V�^�p��2�Q�1�t�\���v�O�1��:�m�ud�r>���ܗ��PşK������h�Q%��FJ�%5�af�|u����3�đW��V�Ħ�h�>8u�4�����V4 d�s �aE �o�i�7�\��{'}.����<� ��1�W��֎�)�{�0�dr�̣���t�<�#�j���f�)��'�\#Wkzcu��t~h�N%%_N�tGmI�T/W�;�ȆrR� �1y�*wb؆Z�O�� g��x~��A[]���z.,�I���`Г��)�K����9����;6��<W
Ұ ؼAm���7�OD�ȃht��uJ0�"�7No��� �'��j#���f���R.�u��ql]�80Z��!�6���������&B]��WZ�25R*v�/����Q=Z��%��� t�E���y�~E�o WKB�}v?�S=ġ�ޕ]�
5�Y��͘�,<Cv`T^\+���OE�o��$f0"춂�n昐��'��Ȣƙ
`ˌ�c�dB��@�u��X;&�����z-��Cɦ�<�iĝD({�?����O�����rŖM1�M%l����h�^��ּ^�?��	f����<F0Hf�h����钙7��%jtU���[��ڎ�S��rc�&�k�-{KK��np(0	���
���y��|A1�����K����L��Ql��Vp!�B���A㥍���Y1.��n��/T苻+��k��jJ��Q�7��cD�]����.��}ͯq��A����x��������"�3\^Z�N��,�dw�C�
�߷_Z��Y��Z3��]��G�����=�G1����?q�ĐnD$ �G�}Q�=�-�@̎>�̒�e�U8��R#*�X���y�T�?��ޕ���'涪>�� �`x�R�k@�̮�n᯻����q��u˛���I$�.p����U�EA���Cs�ոA��D����X�/Lw�"����WA� )�l31�YO?�3t�/����V�N�H=Z[U���\�ָ���\x9asS�����/Y�h隘�Ē0�#�!�B�6�L3_la}ͱ�A�2nM9X	���]��vK���AQ���P$�%�ۅ����%v�����1��c�ǋ�Á����~��]O��Vp5݂�Zў<����>���94~��֚�!�3��� zIDMGH�����|x�R^��mƋ�~	{1
��N�U�(݀ ���1 'k�o3x[L���ء�&͚��+��4>�挪CXp�ޗQ�0%��Ė�t��ʄ�������
%�JpƜT�X����}�FB���� �mu�qo$��|����KT]�!�C��b��R����d�����o�vKvj�ש%>,����Q�nT+����}�Q��/96�������^��㈲%~��Շ:��&I{��a�������o� ��Bf�V.УX�?�<q�޼ݤf���y!MwM�dv��1�Vl ��e���s��C4S3��cw�7�5a�`��|Ef�8�9Dh�?S^D5��)��Kޟ;Υ�B=30� Kt&������5�Aq� �?n$�cݢa\��D�&(��S�d��v�2��ϯK�e�ru6Z��!���kѥ�,��؋�Y�~��^�)�p<"|�YC��A%i����4ljV��Z^rggK&�S ����u�g��9D�@���p�Vj]�؏`jx��=]���=a��c�̂r�*x�N'�T*�ޖ���\�J�<8j�"�.oM
�_�2�* Q�`�����\�4i�{|Qm�����8���B���w���'�����G���"aJ�5�t9]L\�J�#��QFX'���Y�t۸����#��BݔB&����l���[lv�ly>5�w�`0I��#.j��J�P��t#��ak�.|�1�
,?�՟�e��	��;T�\�+���X�s�Vי;��i���|ေC1a�-574f�
e�LR���;�}-�f�i��c��ZɈ���أ�e�uBb�ȧT;�ު�<C�z�ubi�"7E�� �WH�B*��v�8��9���Ǖ���̶��E��,��L�nן���B`S�s _�� KC���轢�5K�����:3g��n�mƔ���K��W\��;��Ҩ^�w�ٴJr���d6Yb�g��913��|�'S�`m�1����u$��A��&2��(0�-�	�S��s���q��>^Ci�w.'*k�sI�~z(������餍D-^�����Ek�*�dܖ��ȑ�B�kO?f����ӗ���6ߍ���M�Y?����]�!B�� �w�ߎ�t�1�=�]�<��!=����~�_�X3�d�7�)|Ѡa�ɶB���c��٨��]�d��y�Ê�������t�q��m�j��Rz� O��p�T�q��J{�1D ��p�搙��4ؼ�5����-ԅ6%�מ�y�b~��p�}���!�������n�t�K�n2�R�E�i�2����t�N1=��e��4�l�2^H�M��t�Rx!ٛ�E4v3�&��`K�\�f���(����J�T�X�d�c���O1��[�X��q���������1�X���#�Ef�Pt^��a�z試���]� 2ջ:J(G׸>���i[�9Ssj���m(�N��S�v�4�5e�ʬ�q���`T��R��%���\Ļ)RX���2C��6ϖ�\�guJb�r�E�[�E�j'@�"[�p���4>��kq�;�\��!#8Î01���Ё)^u2YVw^xniV�m���5�k����,���+O1&�\'&�­ʶ�曉��3����yȕ-�ќ̼aF�Ü�rԹ�²gM��Bq�e�2���D����*�jW7�ʈ��V���u�����;��O��$+$�T�u��s��� ;ǜP��DE�.�B�{+܇bܷ&�E�A'����5|V��Y����-�7 �Z��6�bt�
7��i�߲/S��8=�iy �{J4��Ҍ��tN�6��&m�M��]���ЭIƗ
��l��s�<@�ty�x����լ���
Ha�s!�خ��W,������h�n�8<���ijR�Qez����8���
P3
��cY�9��vX��^l����0�
 �އA�kH�7���i�
Sf�h?_���4���ǗEB!�.f<��7�gQ�gUU�I�d����<�}e�u$��
�TB;���~Z�d����B2,˱?rS�CT-� ��p�3CI�#�'�G�e*�]R8O|�[!;B+�����	��6���P�!յ�4L�qe+Ͽ^�����T[�'-���9\65�wʧ����g��@O)����;�G����g�����9
�������7���B����)�|���'����a��N��Z�y��1�
T"�7�A���Ĩ��K���Se�9�0N�U���8$`݇R��x��p"���;�u�]�T�����-׾�C�����Y���/��3��6����)U���7=�ON+�ɽڀ�v�+����ä(j�{���!��^�x�ө�!e9XI[��5@L�lO�A�c,�~�������X�JƱ��:�Tٜ�G�j"��25N�%	�L�W�ێ ��o$t��� *�5Z~u��eܚ,h�_aH�&t�R��C	?zj&�l���l������4<�[2�}I�T������4]+< n��`��+U�$Ҿ���y�Y�` 6?\���i.z����-��ޘժk)4@j��(�y�M�j-Pւleh�r�4X�<��+�(���XQ�Ew���Z"-D����4��R�1��I�-,;�C��e��=ׇ��ɑԠ��ZGA��($
�#l؋��:_���N)��@�9@�W��كT�NS�v�����՛rD	�C��)Sۄ���S��(�Ê�$+�@��
w�4�ͬ��!e��g��&� ��X��J)hH�1!��5�PO:Y�֝�x4�%� �gj@"�d��iU�\{���n�0ev�F~�W�E��#��њI��N롞+:�8Eh��9d��WnMt/(�HPp_��¦�"P�b�4:����O�S��g�.�p�l�YVG�4Ƕ]���x�w�=f=tv�,���o���#��%%�������K�a�!Y B��d(�&�89����9���_z�������9�l�'��Z�V��Zb�f�O�f�-�n�FȈXLe?^���S��<��/����Z9PwF9�,�Qp���`�}Ç�߰��.m1���k��	���eM��λ�z�H�(	>08��PC��/ku�)���Bsr�.ʣ��!k���>m�l���f�,��]Y���N�A94�|�Ț�b������{8����h�F�v�4UP��k���fL�i���gya/l'��L���� �W�k�S_ލ��5�-V��n�����q|�I
Uu��F	u�\��0%�.�#��1�*\Ye����!+!mM�-0H.�<�u��ذ+�0�y�V�6��D���T=�3'l��^�����W�u�}��qճ��K����.�6Ƥ��m��6��/f(�$�k��c����!Q8T����S�o�P����Fj#��{�юS'�g��Į!L˒���9
��?�u�¹4ӄJaE@���(lZm�$�z�;���%Ļ�J��%�^8�;K����Pz���T%B�A��0xD�᪼�$#���%K�8����
��`��y��1�~�Ү{��[N����M��|!���/�a��)C��O�˝f�ƺ1K?��=��xu�Ԕ�z��C��/x�+�4C�6���iwD)Ǳ8�Jc�U���9�;Ku	�8�8��9dD�.3��?��EL�g��֋"9Yg8z
,L�_�g���幻�$Xp����E���v���h�	P�r;�&>ը��J�1�!�������i]�^A6��>�J�p����#>�#ZT$]/�?�#�I�ɰ�q�S0*v��ܐ�2��g�+I~H�� L����
������9ڜC�V+8�;�\�D�ykS���jF���I�=��L/፫��lRx �C�[�)ad�V�[�h��'���Ԝ�����<��}^�Z�^04�3�#�)�qAd>��$T/$����L��F��}����Q������� i{����arD��.��C�2Z�Dc��y�$���!�_&�Xv'�p�mG���Sg�5���?�X:� �2"����̀x�:;����aL��#�l/��II����FO��d�����2�푒�j�1�R�Еӟ\�r�,t�#�M�$��7p�T����k\:.����Ѵ�:I�&���E��p��;�c��g<�`�m������Q���6r���z.Sѕ⻏/�o�P��fɨ�b
=ؒ�3�h�X@ۜٳm���-J�@�.�"���W�t�^��q�:��8���I	��%7����/�����Ns���y���qVİ�*��!��jmG�jLu��X���.שs(q{���l���n��r ���C���X��2��5������3���F��q7гtQ�97�b g;z��d7f2�I@R�r�������tÊCC�9K�I�p��&���=��7���E8��k<�Ѣ�����.
�
�K�cG���t5�kƫ��πL4ՕC�c�*�x�,��)�d�ԙV��(d���ZX����=Y�T�:�6�_
a-���5a�9�xp����cA�!�J����m�f�csX��F{��^a)������h�{nI�N���".'s�>*��+�!�h��)b�
~W��x��y���B�JpyߌI��ա����Vo�09�1�}���y?�e��t��j��.��1ώ��l�g�0C34���*�jLs.4�i�yM���h�s���ț� �PJ���\	4��a�~�.O2����đF11�!im�,������͓�b��[)͗x�f�G/�mxY�����K�d��7��yH�Ľ�$fzVr�[I� ��a1��a�i�9ꮌ����?�ҧ%ѷes�;�[���j'd��z?�:>�kF=.�S.&�_����	�������j���w�l��;�!�����w�3���[ m����,���M� ;	5����r C�z��E޻���pq���@ˁ�]1_"A��ur��k_���c��D�2Vt9���+�i���`K'�X��l�����̅z��)a0�}�2j��8�$��H������B��Zl��w����b�vu=�����u�R���U!�v�B��r�ĭ�0�<1�Jñ`�k�1��+i�3�h����
�t�������hoO.Yܜf��Ԩ��g�a�C<O�֨�2&ˎ�F��u�=Y�}'vl�������I��(��5�7b7�$[8��d�G�z� �sar�1�]N,���>��A,��O�Ȑ�:��V
v{Ԡ�T�?�Җ*k�㋇�QB�ve��m�,��ɗ7��#Ě`
|fP8\�O�r��Ϥ�ԓ�v�haY�?7(d���� ��<X�"g��_�5���:���uWt��EI�l;�o��9�a�����D�9gl��!^�n;4�
� Qz;����oɶ)W���ԛ�倌�bl�,�YHѡ+_�.S�s���$���8���ء�����T/���8��Q��X�yy��ו	I�4�[P����?��?����נ�����z���坮��1)j�ґ�W���l����C~6�`v�� ���lz��E Ysa�s��F�h�.0xǨSNݢ;�$'~E��K>I! @��~�('	m^$c2���;�Ce?Y��k^�Z�"S�>����g�bK�mF˖�8[�s2�(�$����y�90���/��&����R���4�$��n �s)(�VԴ�B«)
�Ɔgw�ȸ1�(
�WB��a���)_c ��{�����3��޽^�@��;w�S4t�J:�ȡ��ӕ���2�E��T���tZyt�@'׶��H�����b�z�,�: ��p���側�����*��kj	u!��[�����:t4���ct���A�K�U�ݖsN!�����f��B�&ٷ8�{��d��;��M�ixE9�ȾU����\ �!��/�T>8|���M8ˇ�\���vF���q��V_��3j0Z��&<��x�h|���3�U��9�;���Tqݳ>;�����2�w,Kc�3Yk�:x��k��_y�{B�9�$9��{�?j�%��X��}��~n���	X?4�-[�=L��O��ݬ����`����x\�;�RW���p�C|�D>O�5���q��c� !�@&��j�>�@�9�pr����:��J�Fy(��H캅���e�͎zegs��6�O�!�"��!V�<�BF��饡��
s�PTs�\N��iJ[��g�:�i��ւ�is�����֯���Z{ ;ރ����������5�C��K[�3+��Kky�E�N��~UbL�꽠�x|�"줨M��@k*�CD:�oz����Z2���x�_Sy����=�"+M�Bj��pj2&u�GB	�a�"��6zZ����nҫ�C�Ѱ�Uy��3�5�5�O�G�6�8�?76>{��������.��Ь�KC�=<�B��P³ >�z�ʖxJ�k0���8_P��"&�i�q�F�*�qe!�.@wS�G�%A�ƣ��g���C4��76#�����!�U1�&Ȫ�1���H�N:�=�"'}�X�+F�2*T�����Y��*6Ĝ��RT�"���qA�]�;U��H��_�
%�����-҆��1p,݉�j���ｼ{�<��
k) B9&Qkc\k��uX��,w����I#���5�'�Ĳ�|���yz� {���$4x��y�������^ڐC 	A�7K��t"�X�P��)u:�]����b��]�-�c�'���u<�i=ᇪPAYn0�Ui��D�h#�S3ѫ��)����}lM�E�Q`�+��ƿJ���e�����,���h�,H�uX�)K��,~��@]�|D#`��n9ZMhW��A%vf����3���N�pgy����?'*�K�����m�b��(�.ym[��������_q�j}MJ��&����fRH�?�;ź��D���t#�=��?J'vc-Um+�z�#�S8BWs�br��R��g�����d��'�@�aD ��z����,Nv;T���3�Ƙi�a�(ǭ���g8(^���1P�<8���vj�Hf���z �8����n�>�bS�x�U�:G��K-������f��;��ޅ�i�4$�̔�� i�}M�����Ʀ��1z�\Q{��=��&��)�	o��V�&nJ��r_�����%����SOA�� e��~6�܀H�!ö�����!evD=�n�W���!���_qLf�����U-[�ǒ�HPB��`������}��g�b�3�<B����I�xk	�9� �>�̵B�
����R����rn P���Sk��o� $��}��vϣ
cIf(#��<�J�C��[�]͑�����p���<��jh*�h�-��[���������X�D�i�Gs9�B��Er�~�j�+N�e?7t�)���q{v���A�,�v�E�tq�]brq�a�g��;B6�s��t��4��9�`�����\���zNږg���J�=�5Q����&�����D���Pȋ�h�t����#� �<塼�w���;!���%��/p�����/Z0��]��w�[��A�[GeP�����~���I�x9_�#�<i!��ƚu�k�!3v�bf2(W��3Rf,wh�3�<a&!?]R���i0k}+jN�>� S��}J&�YzK�rJ�܁+�q�@鷗��hi�fJ/�A����$��t�R6X��.��M3f�6�^����B�;%zU(^�v?c����n��=��,73�
�H�1]Q�}�P0,u)RF��b�Ⱦo5�#ih�)�")
�?FNP ��w 6"�	ڞOw5x���]c���>H�z�Q����5���LD�
ŨO����9wj.R ��P��w��V���@�F�.��:��ʅ�E�����큦E^���t0� �i�L�6)�~G��1�ɏ�7H�0��27B�ƍ|�R ���`1�R�eE�'�A5��m�$�v�<�k�A��g=�U �k�EVm3p������ps�|�%v�=g�.*,�!IC��J�Ks�A�l�8�bĪR�j/Ow&f�%�!یO ztm2]Z��>�����O�*��EyR�y}�YW��D���l�S������S7u�l �K1j7=���A��1�,�DAU�W:(J�m��%�@�w1�'ŉ�\D{5��84˿��Ci�b��)u�s֨�"��&�g���{>>��Vu� ���#�H��81�ު�,"?d���ґ����v�8�]�6@J������{H(>��l<�v�����l"���x<�s#�A6/�j˲j /x4��p��O� -4�G��'�G��Emy0O���T�0��Oy�;��z<��:WGw+�3B;� �F����ѽ׹���A�3�î砡�J/$N��*��9����1�V|g!�5�M��F�S�{���|�Q�&i�����Bi�Ɣ�Ө�wq��p�����h_�XEH�v�p#��6'[�Q�j���==)�r�ߎ�v��%���K��q�#d�~�xO$���H����?�I%���&��dn`�Póq3l{�Y�����JI�F"h|I��
<��Jw"�01J@yPXDt���o 
(�!���n�5E�p��N��ۯnaH4T	[�kIH�~��A�F8�\����ʩcj�8	k��ڱDUW�\�OG��]�/��=@��5�CW��:7N�?R�p�Z��lC.�8bx�*��c�H�S�,V?�%����Z�lpg�#��1.,\E�S2غ�%����&I,+#�tRZ�$��c[Ig��=4�H��z��Gz?f0��E����\��%�)k��?0�H�Mj��D�{��'��)!꡺�l�����D�M}�p��\%p1.��:`D���D�Vb�b��M�-�I�
tQs����_���u��"8�]&��m�j�W���-��e	���:L=vOO�ȥ�B�K�©�S[�)����f�H� S��ې�2N��/��L=x(�Ξ"c$H_�m�MRhvfŢ:a�dlQ?屽�Q���1.�5��f��3 ��=)v�LfQ���������`o�*�ǻrc>�rৗ͞��VE���!�m��\�ىڰ�, #�ɯi���a���ϑBL9��Y8EMxk�* �Cd����A�C�]LB���u���(�@��C6s2~\�\ ��7��O�wyTVx�����Lt)�X�+�#+*�M_w��kn���*3��7�$����k/e8pr��H7�>g�dh��b�����������4)+�-��59��E&��F�t��
mG���5H��cR��~�~��8����)ž���@ xK$9�Q���T7��FﲆA���f2���i`�����X�މQ����i�I�:]g��C�4L7�or�C�%���=����P�������>�I��3�5�m����h�L3���=�d��f-s6e)�y�i^E��I� �L�U~�e���m�7�+Wbgx�J��^�ꏄ���p�尔�#v��ʨ�q�flm}��ܤ �;0�P/�
�e�=]��\#p:�B5���o��q�Xsl޻*¥���&�l`<�a;g�|:�Xs��N*��R��-�$��.>k�%�e
F��p�l�a�	Y�/�S����oj��	�x���IF�zۅי�^�-�b��|�ώ</-c]i�VΆ���{VfD:��+���c���	�U�# PU�2��}�jwa��V��1r���(�D��$�s��f��S,a!!mXuM�����A7��c��C��l}P���ū;]
V3��1#Ȓ��L|���������i��&iʠY����siKc�>�h�EfK�p�@rE)� ��ˆ�񰓆ШiN�د�di��tS�XԖ�|�&0�r��'���O]���$,Lu���:<7`����Rv�����$��a7r�`M����V�.1���߭1��Qu�by�\��("O����D4��!���>����-��t�=�\��P%��Մ��tt�!�O����̫SO�hԅ���җ�A.���'�~?�θ���G��x�W����]��)N�e�7<�i��;!��:������Z��C*�-/�(a�-�L��(�����	1y�~��~afe9�K�S�Wk��E�N��l���ĩ�|��G�'�9��u-�)���7���<�ҙ*�ugxe��5&/i�8�7���\�
 �U�6����8����`�n��u�QY��n���w8z�����[��F�1Oĝ">��z��Я�����Cԏg\tC���˭�0��lr�C�����ໄ]�ݲO�1�L�g�R�_�����)�c��8��Sfr,:�����
����m���IR�Y�#��+�;o��tW*9q�L&�����&�ua�q$��G����J�Oxq��@<}�n�]����d�յ�w?x~�Å_��"�'X��R�Ng���gLkY� 3��䊧l�d9W9��i%��Omb�q��M���+�R��H��~d�����<�vI�
�g�4�CX_�(��
�u1�ߟ,�gk~w�y����\|���(%A9
�0$���f�k�хF�*˛��j�Cc2���[c-C�,3�Ę^S��׵^�6��r,'i�;a=Q����%P�Q����N0z�l�:q� ��*���Y9;[<�<���-ibՍT?O�*1Jq���:��N%�}���aAo��ͯ�QA� �ew�+k*�0�7b��ɦ�r�e��~T�1�Z�j3-jhJ�� \�4���@�:{�e�W��N�Μl��n?X�6on�U]`޻4�T���;.��p�o�-(����\B䝵vA$+铎(����$Ҁ�Ь�������Sv�C1�{����5�M�ii�gM�(�$����Eq�_:�J,�,������(�H�r�����m�v?C3�D�	���O���Bl�����%�9i9����U:iΕ?s�Z���v�Tgx��v�-C��!��,W6��:�-��z}V�n��w��u>�K�>��F�|h��Ht��H7�h�	im��2���ڄ~�o�=��*8u�D%v�Q.����/Ϊ#>�)H�J���?[q3y��zbh#��c{��"e<�[ٿ4���m�Z̾{3pސۉg�SK���c�6"�Vu�.�i���X���[?`���,��a���̝�#�Jc��V�6�Tʣ!��"x�/T0�������K��g+>X��Ә�5bO�#�����9|��*�sY�Cd?�QR��(J����D?#�j3)&k$*+��V�$�tC.ë��`�k�4��.�F�R�e�W$�	���߲)A�0}��> 5N|�fZ*ba�e+~B
w2v��x�Lg�-w�?[�RQk���ŀ�xuf�s����w^���^�x�Z�A:�*�Gˁ������ܲ3�6�"��SG�36�Ȟ	��Υ�!��d�nh���|�vڡU�@!&�#7ǲ0 {��P + ��C46x��J�@GԬ�Q"[�
E�f�a��+$l�m6P��$T�/69�R^����k��<�3 �tB*�=�˼hc�6�"4�{ �XP^8����CÛD�H�Jhr1�z�e�<ˡ!���F&��Dh7�k�7�T^$�-j9>{Gt�����Ȯ��ak���ch�SSi�s����0ڸ������{N`��U����OXd�,q���+-@�:�z����r� ��T��~jƵ��R;oH/!�B�M�$��\w�a�s*ԯT�rifi�d�M>$�7R�~�#LO��%W�Z���I�����o����)�
���-���J��w,�4$?�M-��X���Ĥ���r��5�n��Mö��.�B�󙥾6�o|v>�����Llĉ&Oi~s���t���1�~��Z���DF{��ނ�Q�q��S	hڰ?G�A����t�`w���2'�3�Sbf�*fG9���f�������vBEy���V%s��r�?�W7h��7G��d��X=%Bw�`M	6�T�#�����hbvD`Fѕ���܋�wKkv���P.�p�$I��=�a���F���������8��4��t5V���k�G�jw'�=�S����3p'4N5�;��u�����ۻ�?̱�ة���$1^�f5�
쥗����5��d>�=-��}T}�.}�ĥ�^u��l�uE^vB+�s8CZ�J�[�������3�\+F��rR�=sL�:Pw-�F�[�C2���E�h�g�맿���JJ��ľM����k�%K#���-�K�����7���"���:�����tY��W�g���P�𐃯;;"ޠ#�jL.�Oq��_�)�jF�.�|�V�L��v��;%qu}�����;Rr�'A���N�����
��pX�I��6�.�!�wW�(O�?|��Ճ���B����0Ix�?v���ҩl���7,;�Q�b(i��j�q�]+�/�ݡh{�	��  �;�)�hx�(�&j�J��iMf�ݳ�K1���
�2ޣ[��#�,�B�Z�~�{���㣪�źȝ1��4ʐ(�1��]��<[(��E�:�f� �cY�ly���ɝ���vZ6�X��t��TK�O�ط^�3Æ�q��Pԡ��nV�hf��\��B�.Б꓀֪v�{Eғ��^�ԝ٤+o�?)��+�B�du=�{;F�V������rѣF/9��iڿ���"�2�S��ٍ�]�ܨXg�u���\��͋lGºKn<����a��Y��J���%j���"��i��`�<�{Ph=?���{%iI36���ه=�-��T���C�S��(lv���\XCv�८�%=� ~�C76�Ҥ��˲^� v���q��^:ƇuX�ظk���%lhB���n�L�f�{�۠�#$�����Ź���]#����7��w�H��5�;XL��D�����Fp�� @�Ĵ#�u�þ��U��%cCӎZ�m�� ��r��|��Ǭ} �N9C�*�Z�f3lZ#���wrc+�Y�� Xr��.�_n(���@�ч��^�`���� �;�E��q�w)��<��?[���J��S�mH�f�]N��´�e/�O(:��nb҈k�~�NQ����H2 �_�$~:��Q��5`����j��LX��S���m�3CE;��H�+%�����+)�tt�A�c���ȥȜ`����N�P���N��)�٣���1� �s&,�6�����ޜ�������qy�ue')cd��h��5H�/��g�c�*�.�i��/:���Q��c��58��	����G��vJ�,\�?�Je�B��ޛN������^ꪰQM���P<i��q���"*���gV��J����,�f~zB�!�}�ۓ��&��u�a�!H!�S�,�n��}.���z���b28U٘�z�x�� �e�CT�Ԛe;`�`1��bd���%�-͌m�N5�^L�š��pɳ=Ԯ%�K���"J~�9��q-1���%�H'�e��U�n.���o�֍�� �ao���!����a<RƷj;IP�"]���
�O����AŒ���\����W}6����_M���3����q�-������9AK��b]���O���>�Ç<��t®������~�ja�3����8E�![�cOL�q�ӧ;�/�?[J���5���[zp.�.�a�
ր�vӟWq�SF�%o�56�f���*[��D�ҷ��Ʌ��m�%ʊ�N 3���I��D���������5:{4X|��d[!���kk���Ghm�~,����@ � T�f� � �A^�L�ؤQ�*;B�����%��l�&�y{������#	���� ��=��<��h�BI�\/B���/�������6�o���}����'�L/��jb �V�0�24���Y�2�Yx��^b�f�M���zX�I�y�7fֈ�`�S� Y�����3�վ"��'��@�6�v{�Ή ��/��{@�''��R��~�D:��x_��t�p��xn�ˋ� �	n����IX�J��&��{��^�/�y�>��ȉh0|?4�q�/�����tvj=�}�����H�?��I-ti��RŤ���PX^��`���o�.yUd6���B�/��VS�?��a�)�4�O!����J��N~�s"a�ʵ�Yəg#(J�A�o�I��#m�Ҧ�M`����b���l��F��d���Os;�	*�t#;v^=�S]��&N,@�D?�\�O��r�Z	]��(��f'��7em�*c���,{�����6��햕�םʹpK2}�BĞ�0��>�d�\�J����c�W0���S�&�5p�?�k�������!�wZ��먘"Qt�o�sq+�f>�959��q(i���F6�7�V�B��z[c�#����y�?>�y���P�Lf-�������_l��ė*d����ʜ +���k6�������,�+;�Z@�Z��q�f�oә$4�
������χ�--�7&b�OM�χp,΋�mgA֫}(1�hنzU��n����N�6E�/l�fݼ��#��Y,O��i�1�S!������5͉�����M�_&�#=����H�N�K�)��R�ڃfc4��Rb�.�����
�Z�z��3yP�CA@��Ex��z$8�u�_PL����~A��ub�vj�^2��)��G��P>J{I,�Cn�گ�z��o����rY�ۘQO�{� �a[�;0�v?�Shi"����˻���H[�ܧ>�6��4;M����Z�X&��F�J|;�-��Jh}k�f�)�5Z�c�Jߵ�ѓ�V�z���52)AEq4�y6[M�"4{ck�$b����Ե� ��1��"]RN�Oa}�|ͼ�w5eb2���.���w�T�C��Ia�B��Rp�obO]1��a�?D�ܽT�U����u�����6r���P@�`�c~�c�Q@�M]��4�u�r���znWs�m:���
t��vS���2�-Y-׼;`��4H��}*����y/��n���Hڹ[%Q�0W{k�oI�~�|S镯�}ؒ���H��/@�}�]5�s�0vhȂ5�X�����w/���`Ur���r	඼ Р�q�W��JC�Yx����	*��"}�	[^6�����^�C��(
m{��o} �-
��0+�������]�f�<L�0�-yj��`���u?|�@�8�
�i���V����<A*���B�ջ�������v$�17�3�y�P��	�~�RT=�ÿ��f�V�8܃^h^	�y�lrو�ѧ��7�d�LL��D��9T��2���7����.�8X�^����6���v���}�E/� 3���;ވ�Z�K��;6���#���\:���~�,# >��e���oHQP�ҁ@[ܕ!2WT"rf�E3 �j�=����Q]\qF��0�s8�{����cڸ 8��pl�6��4[#D�!�4
�X7�#İ82�j��.io��P2��=���I��8�×.���
t�1�@�w���m;sQ�>��2���=c~v7��"�|�g)�ϵ������I
芒���@��j˅�4����亄E7��㶹%��i��. �I��\��~̂�t�����F�A!M�]g�|����^"��e8��c{�s�#�w��S�-�i�w�r��*�tB}���^����#B����;����ϔ���P�a+VЛ�����e?]9��y^Kj��Pg"R���w��ے�v�������k$�%�T���Տ�|����Ɨ������E�������Z�K�����F�͑���O4Uqf�Xf�|��h�6%>����8��� `a�ϰ�Ad6�Lg&X�"��r�tU�K�5sd#_-��Ft%���m����L_��H[����u�/E� �ח8t��Q��Ū&�Ru{^B�%N�,�W Q���%�a�>	�*EӁRw
?�\�j�xL*5���e��i�I���7�>h��,鿧�W
� ���56vM{��\<�xm@�@���ѽ���p�!0)�|T�W�7�����c�4���k����`<���}���R������"�7]J^g1�9l}Cg��^��I�����M]h��RcUI�y��'w�=�,�-ʹ��ss�
rV�}45�t�'�M�`�����XE�[�ke�;��@��Қ���Իʤ�i'�J9d���d��o:�N��5K��?s$�����匮xl�%�3�2��w��^x�
j�R�S5Ǻ��)�濦XI-U�4�/M�1�~�� �]5�Q<�1ڦ��1\њ�N@d��<fq5_��i
���("|�lIx���ΏL���L���܍�˾�<��A����R~�U�
�
��钬*)��������ર��nKiMo��|SF���j��UO0��sTMTZ')�v�[E,uQ�{UD�Bo:�9$��G�P <�9���W�m*���͜R2�twȱ!��zs���R��V�J��6{�?I�9�� CP���ױ��Vk�d��x���E9�w��U�m�z�2|�ԯ�e�K%4�`���[����D4Нr���T/߸CY �pV�bi8R5q��C{��t,������t��=��t��3��h�'�-[��3B+�z�N���%��B����n_�Kk��$��H���&���4��F�Ž5���T�Z�Y���E��d����o�:3�'YOࠀ}$²6�ũ�!i�0���u�y��-�s;��EQ�1n��/�F����<#��W�'��R�\�����f�b��D�V�Ϡr��h�_K�D���9�!��5`"S!��ݥ<�D���W*l ��СDr<�#����DLw�p�T�#��8�)^֬���(�x��vx�ہ��� �|��
�C��1�t��Tt{d�x�2�!r�:$9<�A���<e�r�󆫥�j����?HzX	����-�;��ԟK�<T>WW���P3�ʐj3o��\�>/�Wlϭ\yXS���gS�����Ud1�F�g�	C{��\��+1	s�{��(`�D��Hņ�L�6/��IT�Nq�V�S)��q�r<[4���ލ�p���vb��w�V9&6�e����{�Y�qK��1$���؊-��[��Rm����P{��ai�_�<����E8x��GN�)�*e�L`�F`������6-���jڠ��Q:	q{��qhћO��>�<�+���Qq��b�1��,C�͞ËKڄ�_��H'I,�������q��]|�"V�[�zr˪�`n�O�v�}��A��t=>u�� �#}RR��,��@8������[�.+&!�cÅ�('c=�~	��*���,uW0��nۯ��P�hs{�/�;���(z�kE�3��w_w!�$Q�7�eoDAܷ
nO���b�������m ݽ�Di��y!n7����v������$d@1tid� �ӷ����=��ٰϪ=��X����N�.�yP���������oj`�,�9�9-u�|�x0��� #2��3�5�;!��H��Dd����%r@$~��O�J^�jw��ؙ���Ŕ�K��p�G���>#��{:U����)�\g�U�x #e�{-v���e-Y��0]��jƴ��S�A���6/8�Ó�=rrg��C�k����ʂ��[C�v+�)66B����#��w�p+Z�v.�7s;�Uu�=�$��>�x�>�C�����U�zױ���C�v�Z(�8�#o�O�L�hg�g�	!�����d�����7���E�\�]_nڦ������$�U �̫��cw�؝�gl��0L"3-��������:�?��i�E���]+r�5��_�fκ����?�7��
��F��j}`B���Fc�C����4 ��s��}$zD���,�k��d�����X�k�Is�s=����5����+�8�{�h�����TR0xElZ߱�lF�i(>������l�.(>m���c���� �/��p�;�����[��wiAU�Lk��d���H2u$�$Y�EL����+�7��v�5�~Y�ƧБ��V�������cW�O�b~<��p֞<)/vy$=��U���҅�f@������~�����O,3�e���ߓ7}�I[{s�{��
Qz6�H�d|[�����(#o9fb7�-�u�C�Oɛ��	>�b?�a �C@hr��8'��z���]�Jd2�Ô��o��A-��|���'n�R�����RR�ĿקPabA���%��9��;^[��=x�_�0fe�SF�B���*�O;��#�?5w�C_��ys�.A��� �����_�VG�s���A(X�ViS����	12�RMp~�s���*)�.��TFO�)��>����}~�9���������x��aE�Sh��U���M�3�CcX`��t�����:�jy#�����g�C�诛�~f�A�>/�}�����8G��J'K����yWk)�`�W�z����t�!�4A.S*ځ�?��1���p9B��}�?���>��t�9�;m�>�'��G�Z����d�C��귎�dڴ.��A�Q	��p��Q�`v:�pd�eex:��Mk�Bw�%Q?������<2�������Л_E����]��7WN�!Od�=���B�Qz��uun�5{Ej`��� R䖏P���i��y���1�d�i�V����'�S{+}vwrQkm���&�O�c�ieD�'r�⣚ 'iƂ��*��v#S�eԂP��|lX��s��9������}=tXv%U9+�9,����%<�'������%���!��M �f�M8z��1�g9yȡ�#`������|�f��T����e�ҕ���Mh[�Z��'���ʱa��v�Dy�f̦�ø�9|�Jt����R���=z���n+�ɗ�{��ȇ�p�/�w����'0aW?2ԧ3�b����	���ҫ~U�梙!��$��i�%�A�F%�mq9'9^��)Ӝ�
�Y���D���>1�HM�,�a�����C ���E������X� � �F�&��M�p�{@M���1Ch���0HZ�e����i�`ĺ���D`���m�����y8B)l��+���b�}()h 7�, *F��9/v�;&�"�J�-��z��r�>;�B,�K���\lQ��x�f_��Dp}¹^1\V&:���+A��|[��wz C�k�zW%�ާ��I���&R�{n:)g⹬8�P�c���&п����,���w��^S����ο<�.���Qo]Xsfiq9&�'���rU���h7����>m��s$��K�^B|��� ���/��{Yw�'�(_s�4����~��9�Gm�[;A��U�
l��M�W�r�5t�����Ǐ�)��xGc�o�Kc8Imq,�}�u/���":R����$
$��Kl���j{u�W��7������f�L�u۔�d���\�2�x�ݢ�c��K��R]Wc�X��>��:���"�ʓ�[n/`�jel*���mXJ`� )I��O4ǯ�u���od�z�C0�6`�Gmܛ����(���Uj9Z��h�K�����O	Bc�`��Ҹ�ey���h}�*Q�J=b[�+&:6����U�k�z�"��A��9A޺'_o�
�Cn����s��G�LW7C	=�dz&��^h �/�z@�=8A1o#�&U1�\�sz%C�7��v�ދ(�re�#��Y��k��^Va�� $Q�j��wUe�8ݶϫ��ZS���p�����Z��L3���������C:.��+��f2!�e�9���.����0�������M�e���E�
+C�Ht�2%͘F�o��??8�+���n�t�NXJ�4^���6�}5���ة 1sl� D�~����z�yX=Y<0��>W�=�Gq,W�)�H���%�T�h��	���=��S(*b��#	��#�K*��������F��;� $���α��Cң��V��G��p��ۀܹ�\�[�hM�YÝ���7mU�}$��$U�?}���i�P���_�F.x�rW	��s|љ��I%�n�������O���M����}Ǝ�ooEzr� ��'|���kqh��V��RքL����ZW�[I�'����%�C�Ⱦ������~�#�p���UBa�� �F3�o".z���:'��` �J�Zǭ}4[';*0����G^�L�[��p	�H��?/�Ì��k�����rMZ�(��0#�3�j���XG[[`�,�Ǐ ε�)XQoX��I������p�}j.��b���p��#b�T97���Ņ8fp��iM��\�J,�;�8��]C�:|��a�t�-K�C3�3�]m�leb��i�'�Qx����y�lDH��R���~��'Y!"�R:�����Z��QMn��p��	�R��2��)�wN�{<���]#CN�|�+=�⸼O6[OFl�D�z����D{9���._N� `Uw'*Өn�Sr�+=V���]�����6�VC�q�#?bjoHT!�ZІ�9����VjX���W�����^����K�3��'Uȫ, �g9�Z�h6n��6H3���ޙٸ1�����4�#5��=�>x�&X��d�2�n֫ ��2L�_��%�;G'�ᭇ�ۜ�����x%b�d!!M��b;�r!S�,@�l�n����+^ج�;N�0<4j;����J�2����Ćc��Jo;Ҽ��d T�"�n�k�e��a����"S-�$$�#����Zt�n>��s�SY�)���kI�b� ���wb����*���lȃn��$�*��W��� ��}6��'�������j{�ER[1�#j:d��*����%�B��3��:����]�/=����]9G�V�w��X�����H��q���
*�$\y�h������J:�!,���]�d�kO����P�a�Pp/���ɎȦ����¼s�FTV�B�<h^w�z𝽐�R�Y�B**��*֞C	��mږ*��YGӘ
�&���|�l����8��l	F^����N6mK rwti����6@ҵ��Ǆ��0��GuH�[7z�$o%�+Xií/�.T�s$Re�&�L��O��\/65>�YM�����Q!��N屒�؂'��� J�y�����܊���u���l�}�#LP���ʝ�9�;����Խ�
T�_�z�A'|�ʙ����8m^#�����۰�Sؗ� ����%��I�	��͓n� �Ě�ZLK���X>XW�����b�+ �7�pb�A!���mwӷ�T3y�<�����{J��.*�fO+�o[�vc�H�� ��gAiq��;R_��U���J~-x!�l���6sJdߙ2L��d+{ZR+�����}%�1i��� U������޲P���m��gL��'n�r(�=. 0��Z	�m{�I$ �~֦�UV/[gZ���_TP��:]D�g!f�z�IC��7�ZJ2s}+m��>��E��ܗ�R�Ix�>�<�GN<~>�
he�?�ބ��=(�P���q�N�*%����U�EW�q>��>%����5S�uC����R|d�hx_j��4�ǵ9]�i��%��O�N���
�f�!�r��3���6&70�8��WU[����hnn��[޶�__Q�j��r6�De��r��8�-Xaa�<S���.Us� �߬�j,!D#�c��i1	��O���\�u5J�K���Ȥjp,��e�
�Y1��qu�}ʍ�6���n�W�����)?�-3a^�3*��+�Wfe���kGɵę� "��â� DPа�<&��3K����"�s�1r�^���Y���uc�k\x,v.��Qm'zy�4#]�{�ٲκ�q�Vv�_���ve��%�N�b�#��L8��\�ݮ��`6j�d
����B>�뾩�M<��)�%L�$Lig�y�:9��`�?4kg[��0A��+�-�������!����8|�+�ӄ�K̑��h�(�<���V��� �q�e�v=�E�͚87X�i�Y�����6r�Cn�H�����I{�������2�!v��U�����j
[Q�� z��y�C�է1ܜ�T_��fA��W��.�Р�����x���O���[N�kT��,��U�4�
^�P�q��֍,2�1ƔwҬ�ʢ�O��J� �~��~��?��/T�!o{q���:�!P����>IGoЍ�Va)�=W<o#�Z�q�})B�zӹxDU: V7�9��ҩC�0��9��&� !(��fg@��g�=�:ҿ_P1�s#�� �lHoR�����Ѧ������%�������nY�ձ���Q-h�ζ90J�0	F~M��|b��E�ĳ�����6��pN|aZ���)��&!{�4�N9����,4�ҧZ~�]�r�(�����Ix3px�N�ey�G8�~����nH�ׅO��/�E� ,�rK��KI���s�����=��b�����b���K����z�#z_���$CP���͓>q��% �iYϷ��J$��h9v5FΝ1�`�>����ʂ[B
�~W�Nٰ����k`O� ��b��H��@\�0�w���*�����m���t�wy�T��Nm��� �A��7~���m����7�{1��icx`eQ�yk#ǯ����:��L����z�s�5.֩i�D��W�sY��"��`_�S�3L�(m���J'R����\��X�K�(�����&Aߍ��@������g�Ի}���B� 52V�6��i7U���?Yڋ�ۏ���o'�sB��
J�#Q(�5dY�@�S:���R��ۈ4���%;t���2 )M�p�1�1��w��L���.�%��鎮x�)��� pGT<)PY�[�8H2��QUfXa��P�8V�.�����=5ÁT�'�^�j`%���Wp�Ț[����2���$A���j� X
D�#ȳ̴�2��>|�a8����������りq��T��s��*[�N�A���!�tްPN�_3n��E�+������m8e��A�]��sv�nt	K~v�� 1<��/�|S*N&iR���6�d��D��D�|���Y:�+��{�"�A?+e\	5�J�a�5_4,I�y|�ƱA�S`蒄��8�x��7��i���<ڶ����lU�F��<*,;>= Ji�� �o��B5S�!`I�s�l���tUi��R^f'ʔc{K��T��	mםX���L��̬D��=<܏�8&p4���@��T�I%t���Ʌ����.���v�q��\�KB���k��U(R��#E�������S��� ]�O0�.��W!'���gЍ`b�� ~�-U�O�0�kꜪ�e�Z�����=�жX����LZ�g��y������&�"^�5Ē.\8)�R�Z�V��=����z0�.�/E��g�����Z�p�Ul_��4ao����p�N�@�1@C�#d��.?��١.��ڥ-�n��t�_�)��4�j�C5 �0HO�����d�F%r���K�I�֔m�����{���<�x�(��81 c+
7;��V�[�G��(��G����4�����[ʧ\��?�L����$��L*����7�v��17� 2��:FK�1�9�B� ���զ�o�>�L�9�i���*
�O���u��._��G
�!��`R�4/�2��>��=ɋ��:|�v�>���}��}	��pyu�zJ;^�Ӑh�@[��U�(�t~���Z${>�_��o��S��aF�jG�s`�ʼ0�"�uR�XB�*�	����1�
���,�%*���=���~��Q�a��QL��,Q�t@K_⥥�X���7_nj;�]��ՉՋ��̼��3-�D��ܺ����� ���x-|�&�h��+ �$;��uᒰ*�Ń��d�{��Ά�4:�<ן�4�� ��L,�*��|;��3�tߌ=W�'b�l� �9�T(V�u���q�r	y[�P�&� N�����?���T��7_��F󒈼[��;b>��Ҋ�Y�F�r@S	CA.}-u|?\�Gf����
ޑ��oE��`+��?m�y�#�5!���G1DS��`.nC�m]�*Tܳjs�B�~R
�w�������j�$��.�����X�稰�r�w���Y�abc$�p���]#(�c�X�V��Sj�~�{���t~F���~�]!m���Q.z������v��a����c�`@�cD�-4����b�$p�\k�&n��2�y[�l�Jus�V���R >E����f�I����HR�ʼ��`��}~�wwq�Jo\ߐ�RW,�΀=~�j���!���@��;��z�y�8�fd�z� n8= ۯ����?�%�(�~H]��v�U��Q�	�ո� ��b����y�����b�n�$�Fҳ�U��>����zh�n̼������K�s7��}��w��5��g�i_�ġ�D���Pr����\z��28���[�n2�4ь��0�$���)t���Tݞ�@{�t[y��#͇�44#�}r�zde��Zҋ���T�-����"����rD�p��A���Zjȏ�z�!9�����'�aQG��:�������/t��w}p��8QQN[�W6������L���vYog���a+�buz�r�*EU�B�JdA��A�#��ȧ�e��	�Dޠ���o��3`�g�`qcR$�K�x5�,��Ƕ��u]�O���w��
OI�p-~����P��B����?ف6�&�,]&��#�"��|Йg�:&��>�h�$�����f;"�Ph-M�&S��6��7�|JO��ZYx�.Z�	�f;y��{3#�q��В@	�N�V	���'����� �t�W$��#��r=�c��w|��8/��W&4���.�qqˁ��p��s3� L��%{J!CK�1`�,�/Mg5x�e$#W
����w ������Z�
���8FL�zK��c�a�I8�r����<`߇)���͠C:��qz��D$�����d>�1�i�d����"��@�lhK�gl�4���y}9�>q}�����:?a�j�4�P��16�t�����,*k0eJ$�|aŖ��n
��j.�K�}�4��,\
�j����	4��(����X7nNb��~x s� �R9���Q_�#�IV�Ly��+O*�ZzMh�3>#70S����1��@;�/�z���R�*�z�=�n9�b��힀��|��*��x��{㏟Px�`���6�g������T��J
��K5����z�o���:��P��4N3'�m�<�4G���h\V*��6݃�[<���M�w
���r��{�$����8��ߎf�����QD〤�+�joTA�ޮ����<~��-Ӑ���؛Cѷ����Sҥ���:���{�?��G%���wW�	�;T��3*E�Y'���)~�>����VF���n��	[Q�0C���4��	hB������>�I8�A�l^[��;�1}h�ni��E�������c�G)��UΪ|._�Ǯ=�]P�<���N �f꺨��q��]�U[�	�[��,�b�m�fr���	ە瓕�T�52��
��=��o�|#�m�dk�r�u����� ����ﺘ4�B���M-��J�3���`������s�7��i�e�

^�|
��|z��Sy��C8�ğ�qq�s��_�8^�2M:ޛ�ߤa���~� ���r���V�-���%�:�ٺ��<�Oy���v�!]�XG�|x�]4oI1x��d��
;��E�"M*�``�Eב�����3�k�	?�ȉ7��\��μ��[���B?���a�|7��L�QBP^�!�r����=��{�6��k?7o�i遉*
�V3�1b&^G��@4R�B�أ̘�	%�9:.�C��Ɓ���7�$�F�?�G�I�H����s�)�#��x<Ø(�6|X�D�W�,v�� �p�<�������Ƀ��T���Qn�|�=���e3ā�ɗ��K㝾=���겋B�b�����3��>�=}\؏�b�hm�:B:���p���^o���������I Y5�ґ�&���j����־�~t��"!Y��U��F륣�e�K��]ғU���fy�k_�P�	èG�~����`~����db��>�r���2��Q~Lܤ_>dZ�3�΀P�R�c4 �4��/Tz�{*~��e�����?��F:����"M�
\G�}�h�����j���hyv�*��&�?�bom/\QS�+�U�eY|F<�D;�q���h�4���*�n���w_}��~��&�>K�G� ��\�������=xR�:yry�i����2���T����� $~Y�;���M�!�!��f�s��F@E��1�#����zo(@��Hw�ޘ&�.e��������(�=�u"�C�E���ϼ���|�撋t�k�ԡ��z�i���hG/�;"YC�����x����?:\Yy|3r��o�mekɜ*�%���ԒŃ�&�� -|;I陲���[Y���`~}# %���/h������L&�(�
��pN�Jת��o��R�!jQ_f\3���5졼S��T0 ~�Of�4[訏D�ÿ�e��\��e�b�K���
�l�C6yF��D�F��'e�j1	�ᙍ[k�������IKMxm6�R��s�>]��w�g�Y��.5����I�����0�����EmKT$3X�)}�(	���<Q�fN�D�J�7D��d��3-X>[�`��A��{�b��0�2��S���\�{�ה������,�+Y��~���b���h���B���@\[�B�����b+���bGL��]��% J�� �V"��<l��n�
>�y�^��!l�9�y���xL{��э S�WMz";�1ӳ��!�G�ܛH�p��b���q؋��	U�F�=u�(j%D���C06�W�,iTx�9\����]ע@&��m��!��請�C���62�ײ��a�����T���ɿ�7	{ĸV������qE��Kxq�Oԛ�h�D&_)��9��XG�š߼&!�(ŵ��԰=;7�Sė A�:<���D�}֊�w�z��U6?Hgͭ�۪�"�ީQ�uD\�2rR2iS����X�S���Y�Q�k�,0MgJȹ��Ne�\ x+d��v�L����j
/�����:D^%�N2�(ś�iCy�}�\_c��^镅�7��t��Nk+.R�)�:��QD� Ҳ߀�¬#�n�< �rAf�fN�!�P��r�ϡ׸�ֲG;=CY�S�t�TdfZI�x��@�.�|�7FU�k�����w��k�^���?]�%�a���?$�= a�>�99X)6��w
뎂�W��-�����[���1��yLZ�-W˝hWi�hq�ֺ������� ���EKZC�-Q���)'s[��7A;A0y p9�ܔ����^���&4���V�� ��#'�8&i��p����U��q�RS�O���V�w�A_A�v��q��!	�iH;�ʑ�0����g���G�D�C�[ 6�ƃ�F�μGZ�<�̵�m�g�]�ނ�j���4ҳ@��V��i�z��\��m($q�@}'���aҐ�J��0�>n>�=I_fheSU��A�:�k��?� @=N� �%�g�&Ý-���<k#��Yq7�����$������`�S��i�E���������U�4���ND(����{B�~�e��ۏ�zT�MP�vw��&j��ү	>��nOq{̠/�a�����j	c7���5�}R�%j�0��ٟ*���`�S22}@����q3�j��]�N+8���3�DGRi�u᫣@��rVs�)��^���<V�I�'q��ji�����.>��/fe���@��s\�f��D{�E 6��������z ���1�
��z3���xB��o�K�6܆ikM)jX$aj&#icMV��k���@��#�P��#�nD��5�Yej�[��K�#
���Ra�ݺ��3���x��$F��H)g=]SO�0���л"��&�	��X�hok��hI�
�k�$����mA���Խ{��k��|�V�apb�dl�̎�����4���!���*�yc�u�%��Kt1?�n����=�_�k��:��Gu���:����$o��p"��	��~Yb�����ֻ���ʉk]�f�_��i�&t5���P~z�'U7�P,����ursL[��t/r(Wd_a�d
,����*q6.+:��¥��OF�<_�u��(�bF�q�tY���ͪ�^ �4��Τ���z�*5�WZ'G���P��e��z��U�R2)[i[_���0x���'���qv]���+��}=���O�@�gm�~�L]��E?���:#P����9�OcN�L�E�x�+1f3�ɜs�ڨ��g�>��-c�oP��zZ:��
��&�֝�s�W;}�H�Ǌ~HN-6��+�\H�� �/�8ۊ��c�3w�Щd	�����rÇo�)�s#�����iЮ��b+Mˮ��J����t�DЈi����Lai��;J>��c/�x���cd r�-�X����@W�������^��k�*x���J�<=���iT�+g���6R��IU���~�� @��H�-!ģ��<�_^���/��2L�5(�?H���&�����5q+��%9��),%u�Rybq��n+�s9�=�pHZ�_<���Ñ�1E�n�+^��BU#���fI�箔y�+���@�W�䵩x�����_*"�+�.`��H�vC�_~���p�?4�t� b,`��o�N�T�����L�����H������od�3
]`��^3�������ݸ��<|4�r���5lPu�w����È�g���᮪!41�T��W^�㫃Ԭ�����d�ǩ�׏	��W�J=�����)E~L�L�i��ࣂb��҃r?tȗ�-��P�^"':!�E�VԃБ@"�yགྷ���x���%q���*b3��P#`��.!QSŴ���H��V��n8�}�7�؟��}�$a�aM���:�ftU�5�	XS�2��h��Bdz�Q��y�bdb��)aU��v2u������������p�	Rv,��"^��8l���t�$0��ıu��@�8@b�?���x�O�G/�3j�L�2!���{4W�X���/,�5|w!�o@vx�֝l+������q�u?�4�G�2�k��[{µu|�ѫ�8� ���%%�h"�����8n7l��M+IL�Cj�sཛ�WW�
�Ցs�z.�=tp����� ��"-�g�o����c����kӈw̆z�d-ԅ%̛{9��&H�N�M4|�A(r=U�!�V�4(�T����E���I�4�]+���$��� w�_����ʘ&˯cbba�b��;��"���:��-5�oD�]A����F�
��� I�����s�@
�w,I��G��Pb�vXw�*�4�6)a	*ݪ���"�h'paÓ������os�<d��ՠ��-W���MI�*MEh�S�[l��u�	#V<�W�]ͽ�t7�5��M{���٨5�3��l&\(J�O@Q3�8譑(3�ÿ�^V<�)�X�SN�R X�o:<�f�y�:0 �}6Pz�SD�T�)���l}x��B�tcΖ���#����Ժ��y7��(�YelLD�alIB󇵛]
9�V�yy$�;�cM���Ug�'8�i ��nL,�v=�gn/\@���j���Pb7�;���W�����Me�}c=�1iT����H��b"��<(C��0���
��/��PGc�=/!uL��[�Y����d�ö���Xf���T���O��{Q�T�;�-�u�[}�;���&��#b�e���M�_�G�[B�l#��B�_Gv�p6�,�Ą�u�����x;�A�O����JW.��#�/���������2�ľ%�z�^��m�$G�5EVH 1�q���D�����簍��~�Ԫ�g'��\�+*�͞�R�EA<��-��P��j����L��h�X�./am��/����ѭ�8l�x�ٺtJ���J�K�����p!ɬ���S��V(����E�O���*%�S~�}�F�
mJ-�a�c�.����s<�x&D��5���C��� ջ��萂S�����E�/u�J���|�b�H.��l��a#sQ�V�O#n�f�	����~��'�@�=v947^�r赐��v�0�u:T:.�!�͉�Z�0��i1a��U���>!r��s�k�|�9�Ƅ�b��
�ڄ��{�; �)p�)��%B�X�`��o����'�����O�#h����<x���٘�q�˱�&l��dT�ׅ����e�X����ؚȒ���s��Z<E�t܋l=��|(�/��<�_�`)�T;�3g��/�EP&�л����|� �bE�禥v��ՙj�U-���/WAr�-`�=�?f(���1�`j�f���HG����u�Sµ��v���pN���U��J^���VU��
��'TBغ\J&�
G�#^VA�����y�u��Wul���;�T�ǭ�f��l���-0�RZצ�-�\���ݩxa���/ ���gOZ�V�}Cu��ʓg�u�2]~`��FKw���o w�.��p����Ȯ\+��1*�!�a�nw[fж��˒#�(���w���W�\+���i��"i{x��z��ܖU>]�ԙ�U4�Ŀ'�$$M����竂������P�P5 0+��Q?��*w�?���^.��1��~O޼�F�p��bk塇�;�I�i^��anta2��"�Q嶟 �� ]CS����?c�v�bO^C�n���S��:Aa-6V�B�r�&0�"��˜F��^�˿�&�I'̤U7����p*7^>za�>�
%��8쾺F��)Ζ��S���\VƑ����O�x#��Al�.Ə>5z	V��HpڐyofQ�y��H����͕q���m��ɛ
4-|+�����U_|�&��G����~����ח�D:l5:�zzRC�zc �y[g����L~�x���?����	�#�*ͫ�R��L�%Uw���K��_8�q�,7���l��@��M���ܶ[�ڥ7���/V{���d�9A�c��i&�%�l�e3f������ �U��쓜��L�c��!dW��u5���O��e��Ἠ#\Q��M��%�'U���3�+�<�r��|���]��ic��RZ�e�d����1E 4M�G�98�������O�4�9�v�PN-	nY�}�/wB�f�M?
�����[:��CuB��H�YZ����{��=�f�;_f%���OIA�8m:��pzu�\���nZiN|��� �$9���>&}�������Ѐ�^�珴{�Wť<>o���g���Si�g]T�C�a� .L`����n�8�9BG��_ݱ�}�LR�1`��g4,�yL��]C��,���IM�A��3�l�U����Z��5��	53��n[���YIM�mY)i�?S�2�Q��NCmk����å1:����W��ʯ)jjD�vO��<֖���PL�\n5I�g�hp�9b>˓��۞���m5+"��0�Ğ����	�P ��p]�jM���JP&��ىJ% n�J�G���)ky��E4nh����Hf|��B��+D�h	ggͧ{��H�k,Vt��M��h�%���'�q��$�쯋ϳ��j�^��έ�
6�5�D���y�@o���˷؀IAV9�����?���H���_7m� ']�&Bb[��m�g*�܏��˅��Ӣx̩)�a�#88��w�E�;�ǅ�u��݋o�4��=_���j��b�Z�nA�~(�A̓-|��Q�k�X14�T,�e���h1g$l�n���Y���
]���]n�rz�D*A�Y�����x�EJ�LX�<Ǡ��-���NT�`�rV��x�ߩ,96d!S*�un�i�M�v_j�2}zmn�$�?Ѕ��@�y�]?�:*�|�=I�X]��T,<։�������������ՑA�,$�bGcn�ZN����5`��-K��>�i�TE��Ռ���e��4/օn�,D����ʗ��,dV:`�Gm�����$ΌW��p e�{{��P9G��!^�Q�����pSH�-��J;�xƏq.�|�2|i�3�b�a,��E���c3k��i��mD&�'u�̌���B�k۷IUH4cWN��c�w�$�(���9�M�+�����{�C���L�te�I#�hv��X��m�J5ț�����ᯍ%z~X�������5�y���ӈ�����x�$�ԙg�n��}\� �uTe�����M>.��壛I�&�Gq��T��1ق(Y͖[J��^@[���Һ���vxot3aO�c�������7������z?ٵi��l�g @<Q���7a�(��=n�o ��ĺB����t�l�WK��P�����N�]�VL��Ѣ��G�IW�0ㄞ`�(,���ì��d�ϦaH���l��Þ����6��ׄ�kd%����u`��={�m�2}m-�SH�9+RG���J�1��{1/��G��ӁȊ����Ԁ��mY�� \w�"Wf|�`I��⋛�A�G`�ٷ�,��4�%Z�g�[ԇͯq�>YPDc �{l#�*��L5Mh�<�d�Y�1�����������P��gI�$�;�@!J����e��P�|�D5l��	�<#��~��O؊��խ0�+�y.i��é�p^3��~g�x��~�kr2�5����NK��!;����T�w
�yٖ�����m*!C���@��G�vom�>�I�԰�����3g9'�s���9��u���3k��5�m�u��J֮Z7����8��K��G����3�\K�(��9��u�� d��~�:�1��!�?�����?#:�qa������������{_�O�x�Gm�$��&#��W�k����JIwGe!�~����U����B�k 4������A� ��;[ca�^Zp��ç�}^�b�  �?*q��W����l�������� �t�*?�2��
fiO3N�6F�s�!@���� vmS�p�J0�L�d/8�b��	.p���YC���MGy�S�aX7���ncq䢇9��
_�}�nC���G�W�qS�\B�K��ɔ�-ғjW]� ?�K���ۉao����|O��I�	��S��'-
�;Cn�2(�dC��@����p��`]�'��잦�� �o�靏Iȼ�:�<"Ų�0+�k=gZ!:�M/��Q����`�QP�L#�a�~<�=���&�V�`ᏻ�IO�\�m���s�O&P�dx*�`R�z)H��gu�����*\P����A.ܛ��U-�!	�4�
�/���K���,|���+���1\d�3�k�h�6^���y���!�`p1��,R+��x�s����@�Qhɇ�v�WrǛ�+�9�aU��H<�
9&��衎p9�K������[B
fhQC��=�ݧ�9,Ǉ��A�/�+Ǭgπ���͟�����[(FըwC1�<l��(���⮕	pC�m���A��<��������	}�7�ئ�y�����3�j�}����<z6�l�!���.7A�i�# Hʆ���S��ӟ������C�+,��[<D�>��VGޓ����·��K�$3��K��a1��)��40=}�����p@��ܾW�y#��$%l(5v�!���#a���ɎQ���zLr�&�55#4^l�5�!�8k ӈ�ό>>53�:��X<�{*8T���^@`V ,b2��Q\Ƃ�@$�)����h/�I?*�v�z��Tj�{Z#s����(7��9
3����� �+�S��8����&+��[ְ�\?w����z�(Y������A1�]�n��Z��+��&����X�s�T�F-��Z��M��ӵ�خ�h�A`��^SH�M������͉W��W�-��� 1���=���\J*��|�%oIϾMqL�ϫؤ�`O���	J���������`^��G�o��M֕5c��чq�
p=�k��{x/��s�'F��c`b�(����!l�}Di�hH���hZgW��7�=�Z�,~��a<�.��v%�'�t�O��>`bM�aM���յ2E�&�os��@ww���w���3y�g0�JI2|SpL�{�;����>����N�r������ �op _�X��g��uN����ڼ_�*�|���+%��
������X�4ņ���y�S�WeB����|G��0]�"FZ�T�╗��M���3J�R�A�i0�-�O�x�rs����7w��t}�_�R'�T]� ����<:E� �\p��?�<nd�1$3#f�<(���������� [ �˼z��p<ѷ��#�I2�����
�8 �ײ��|���.����Ÿ��}F���̢a�f8g�[�d���'��A7nì�j� a�� 
��H�[���.r�
��H��p��@6=��Yķ	�����W�L	�O��ي�ݮ�Sfʆ������0��V��@���L���������O�o!�%w�@�h�%bn�TU�Ch8~�?4HoE��k�7o�!;�	�<�=��}��/3���Ba�V^���#��u��o�Н�w�������b\ UJ���� ��QKn��[������C?��[qG)��'���Y��:�� o_�#���������tׯ2�OZ)��m7�f2Q�,,r[�?���z�T�R}dr����}�NX]�V��O��CWj%�ٳ���ad��A���Fʏ;\?Ǒ|E���W;���g�)Eï"p��.(0��!��ϛ�+ \Ф�M�ޥ��e�qį[%��z-8>�����跟�,��(�T�a=�����f8��Ȭ�^��;1�	A �eF����x\0	,}�)ɊO������
���˝��jߗ�������fS�C�B��1-�<��ې�%��c������B ��q��b�R���ZB�؀x��%��n���4����(���hw�o�O��]=�SbΏ [���'�Z�����E�a�\NSų�|i��W����^1�xr'��o�<C��U0�k5�a��d\�>3v�C��2Y�v=��0O�����Kd���8t���M��WU��E��-��-{ӹ��Y��2�ڪ>�	R�z&��Fl�tˆ��H=x6Fu�L�ש q��#Xp��cg��ެ'%�rī��:��N%�h��b�C�IIP�_���*ڦgQyB7�Hٚ0@r��B������^���Tyh��y �ũD/>9���b�Tk-H)Z�����~��kD��1!n�LA� ���M��|P��2�9��Pl��������%Ω��.fϔ�������^^
�72�d|Bb��.�ŅDY��Jg���xQI�
='��ؽZ�vU& �؎xk��V�t�iV1��q�0a�������m3\����*�>F?��'wW�>΁�k�ViN�~�X%+��>|��,uw����)�3h�
U<���I6os���x-R�lB�Q�W��^�+�x�8B�)-R�i
����#9IX���6�b�=�X`����V�^��-�ئ ��g� �����}D�Yr2�~-�r�a��P�ȾMَ�R�j�v(�V�����g1q.Mн�ܜ�Ó}P}�Fb�eF�����{qݦΦ�R�� �]>����j9}�l��oD�"��;�d@���݁c�V���o���Y�G1?R\��Dn"z	���k��C�X��=}Z�2�yP�R�ᛝ��n{�h��B�b0}�E�7P��tƪ