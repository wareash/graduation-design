��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|e����M`pہA�Q�t�J�(�N��d�[	��ʘ6rps}Ք�76=�����͎;M�w|����G��]�n ��*�)5�sQ��l���>�a�n�>]J�0E.cЇb�Z�?�`j�@`�����eR58pH�+��	I��>B��,��]��4����C�Ȅ�>�v-�8FE��UɱO`c)Gc�F}g �gt���a��]��5�V��!��aA�D�;��uP��S�Je��ET hA4Oў%�긾�C�O�8G{���:j���cp U�P��'��f;��D��,6��v4j̝ݲ31N�v٠��cZ�3�^�� #���Y�Ĉ�2�m���̑��R�bzN���-�F@|<Δ�oʛn�,�����ib�s(÷{3�l#��Ԅ4�:'�����	k�*���aկH�v���� :?E�D�{_U���S��i?>Y�Ѩa�.��:�wk�Ҥ��Q+(_\x�HmΜp�-3�O��e������T����䡠�/Sp�q��WD6��R�$U�Δ��;����ڍ
""x��b�s1/�K��A�82��̢<�yi.G��q:���5��*��c�0u6{�[5�՝eڪr�L��>:O,'F�Hp�ib�K��F]���_+Qv'�&�fu�͜S"Ma�\�2f+�2i�6}��I���#���+�8x�S�F0�@R&7]J���|��;��w�"�Av7�g3Ct`�'	��ow�9�Z5#X���:��B�p4?c��KC�����1�޼��`d�E�S~���f�u�+@�!.MhkT��Ϊ*������2F�]HrI�l/`��-6^������Y}rX��U�����ݡ�2x��*΅��Y���x�q탊���c1mq�
���	��Y"#	����e��8���x�M�֜d�*�,�;b�-ɕ�\-,M��S������O��^)qѲgq���{#6�Xb�쨢G������S�t��@'��(*g�~��P�>������g_�~3���]OZ�_�%DG֘�'��\2<�P*�A����R�� h�|�����~���菫k�5���8���l�[�fw��+�?�;i�V��ߜ� �Am�X�����7��8X�X�QW�^ji�s�)�!�;�m�� ��?���vP�ز� �5�i﫺kB������3� ��E�Ք��8,�������&Yo=��1�m�f��;p��e�+�E
m��5f{Y=�`�n+Ij�l6����4�5�L��W���K���e�Z � �8@�"�uH��|�H����Ǉ�7�V�<�j.�(!�ɳR��}ͣ�o�1��t�=hq��LԹ���19�[
O���2]�!^�z��@�6�Zח@"��W�g�ŔЪ��l�V�nKe��,P��;���zi����:��kF�d:#��Tx�'�����IEȆ�Gg��/��?E��;Ҹ�9ǝ�V	cW�|[ݶ�����ǛW���$�tSO*��)��.H[:��a���[�>"���sŤ���07=�=|�� ��na��C20 ��k_v��@�\5�����KfE�GO���ya��:$���6//k��uZlr�v�A��v�]��#0O�+z��T�YS3���X2�Eႀ�cCҢu��=�Ls;���LDkBZ� [0�*�� ��v���D=ƽ�^:L)�r�	)���Na��^��DBysS��X���qi_�a�����Z�EC��/��\�#��i+��͇�:u��?��@^�r=�ܣy���ܣ��A�7�Rs!|��˺�bt)�#��?4g�L�����lļeMF��v*&Q,<��H���D��W���f\��D�,��$���rbp�_�����8V)6Z�^�e�����&oC��k|@!҇*��Cl�()0Z^��=c�<(fdH6\x5�hX�2f{��幁�1�#3BHo�M��.GE�����&�;j[m�`�!���oJ�T= �'J�����i�U>��FpG� ��I.!zvĪ3��z��h��qM=m���������0��w�dF�hl�6�7��"�!�˘4���v��>��L���ܳ��<A��:h��t�����UD�Mk���I@jO����c.*�ĺ�b�V*n���5u������]�+G	��rb����խ���@T�j1 Y�Mu���_3f���to���j�� �G��)M��hI!�Ҡ�a��8ʑ"��/�~�e�]"݈La+[�I�����P5܂�g�O,&\�z�G�פׁ�z�w�_�����Ϙ#&<����O�� 'b��I�r�/H��(�#B��Y�~&��0���=�v*��K�4*��M���zR�MF��{.^B���H{�E
��1�R(��y��&��0� �����m:
źg`OR�}���^7��f6ǎO}�N��3|\�l�,�(�U�d�N��9��D�>KBeuz�3.���5~|���T���pU��v�����B)uZU��?\M�~��"���mT�ey�Z%GXo�R�һz�"����9	gy̈́�E4�WƩ���7�����'�=ɓ(%���?���u��01jI�-���(����札7H~��DU�;�fO�Q����sĿ��mi:� v5�%�C��yX����O���V��'��D�=��˰�n�O��seg@c3��� &z����ߴ�C�	�3�J���O�GlD߰�$),uK�FB&Ǜj�˧�
:+Ij����A�y7%ǩX$~gA ��5��|�N����QƁ˙���b������0��3X�)�]��a?��1���F�u��(."�PDϭ�R����/C��	ű����>�Cm��s�zN�Q�3`N-���)��,.���i�,�;�]@7�f�D����N"4Gj����vz$�́����0w�'����2�n$sE����!�Z6�b��L�md%�1b�j��n��|#B�voU��݊T����m��{��u[4�������)S�R��x;�Ն��x5�\J�Y67G���Z�sUb0��5��/#[�f�8�
�8�a���$�?��f�[ʖ����i��V��;w�R��2�,ς���T?�E�5�g�d�+��1)=��'Y^���ʹ8~���5p]���kÅB%�t ��^e ��-JG���֠	�w��MW�E 9����$a8��J���¤�~)I�d�I:9��gD�� o� �Z���Q���(���.�C�!
f�EIߵ؁1�H|�f)�<4O�V�YJ��u��b��g0��Ro����\\/��l�@���'������N�/"L;�D���
�����]LU�=H^��o�-��v������Oa1a)�Si�(�;�)�mth��=3��V��!��޳���u��t�oy<Lc&\##���
q|*������4뿊���{F�f2T�&��B%[�����j�.��;��>W���|�DTT,8�5<�z^,R�1��j�,�����*�G�e,�.�>?��� )M�ETۭ�Q�x�n}"�&D�M�jQ(���'�4׼~���?�'�{*�FH�%R�܇�X�f���O#d���ĹA#]�~�g*)>�'5_xV䯉����0�
ۚD�(�b
�?��i#��τ@� �/��$f�)�(�7Ӥ��sւM�՚�dM�'(��=�����������'��hP�hX
g��I�a�ntw/�Q�I�KO�v�c.�Dc�����VM��0�_�C��P����+�����u7PM���ǐ�A�/͝��[J�y]x�WϬ�y9��drB��:PQ}�s�r�:��_͏ov�E֗s��[�h�� �R1�x����m�'�ɕ�p��4�'Ì8�<���n"�����ؐ�oh��x;:�c�E</�@$Ä.p%�Ŧ����$����A6VC��P�3��v��.nO��b�,��O����<�s�_�Sy�P��%�s	���i�y�9Q������=} �Q�z�V0 �����x]۸ �."�iTmaC�����yk G�w��.#QJ������
L���X=l���R�
ɕP�q������>��1��HNU�
j����;r�NdY� ة��R�u�ĭ�YQw�ؘ���$�@���٪�;�H�!��7Bb�+L����x|W�����#����/2��q����Lk�d�Lw &'�������U>�[$	�q5\,��{��IU�3��h�!"��Q��t����K�6X�2����|��a�sͣ��9Ʊ�`��!٩}�ȡؓBM��h��������༐�eqO�*��o��3rM�49����������Fc��T�g���+҇,�w��oB6o[��	J�I�9�~�p�����ލ�5F������2��*�m	4$��/� {�{��R7S�$���4��	����&�G9�r�pZ����/@��JR��^<��ol���{D)@����S�l�7{7ϊZE��������Q��t��)��Yp�˰TK>��\N��[�+��d�{�_,l.(iBSë���2V���]����|�0�T�c�:�8�53���ɴ��Q��O%�� ��U��%�^m�������B(@�ߛ����,���*���Lv�Y)�X������kr�m	���
a뛞��d:�Ѣ&*$�,]C������Sw�t�Z&} JBY򇘥I���H��o#�hrG R'�t�~_��Q��~�ˁC�~�@֒��#�YRs�Mxk�XƆ���<�	�}h�W��ٛ#������;�� ����0�>
V�@��^a�	��v�<��;荂Z����U��|�;?��x�+۬��\� 9�����EK��՟����sit�� +F�+�,���-Ɋt=�%�"�����z�9��A�f������E0�21E�"�U��#�Iţb����H�d�(waHZd}���|mG�nǾ���	��C?)N� �uh�_���'}��4���k��������F�J����LI�~gX!�_���{���5� ���3�����o�n��Z��C89������J�6����B\���]�8(J��ۤ%����A�.�� b�>g|d��=��P�Qǣ�#���%��~�ޮ;���΍&���Z�"���f����o ���V۞��9,�8���m���1@7�'�~w�k���&ӷ��s'�%��� L[�۝�W	�{#�qL���s:zJ�l[�W��/W�K�I��ܲ�eV"tM]5�_�A������F��������Vi'Kw��vXΠTd�3N- $% tx;��~QTd�� �M����unn	D��n��y����g�ś�y[�m�5�a��:ݩN�'��k��$A�&-?q���F�M�p���Eg�gL�ul���LOX���`[����`s��X�� �W����M�qL���� Oɰ$[-+��uԫ4ͧL=��N͑G��~�a���Ha5ɜu��ňP
3�9C8��/�M�rn(�%�:޲	Gt"���a���Ҍ�1=P.�˒�������'��aq}���a�!>g���r��_r�̴�3�cȽ�hz�:����-*ԙ�E�����bS>�خF�?��b8Zz���qR����a)��M̘��~���Q]I��^R�0*b��ݰ$���g	��� ��V:�B��Q����pK�g-�ԘVk�|X�"�LW����,���u�&ZT��Y0/��(�G<�+1	�}�}���Jy��wl�RT|�@�w_UL���V]��*��6���N�=�MƧV������`ֱ�UO����[���U�&�:I��~rv3���ϥ�N�8����8���� �
�p�S%9�m}�-m��qW�hV��hf��tG�����`[o?���/��W��8d��Ŀ�"��Z�&p
$�HS`z2}��[S9�Y���K��єM�UҵN�4��0�W��+���GN���8T��7�mȢR�F���-�������e��])��	=�&��hu��8�ױJ�i΢���?�lD�Vcm�Ъ}l�&�ؿ�I�iU}�1R������?1Gy3�mj���������[��lz�|�8K���R�N3+�1�XC�5�T=?�6����.��ڨ�HlK����J�gP	׿��Ϥ�����V8f�q	�����W����'�s�?���IQ�C%�)"�Uo�+��R0��՗{ˏBQD���62�c)o��fo h��F*W�FC�P3�����: O��lC�f�޾���*Paڢ�,[� f���9�f3yc��%1H���a�ˈ5
����*Uj�(�@4��Iz��[��YW)�{,���K�z�c>´�Eg��RFY�}[;X�v_$�3��Z)(������߫��t0��ە�Fb��τ�]��&�9;n�~��v@���@���s()�D�f.�6�� ����Y���14U�Y��[��*�%L��fY �<��١`/���@ϽZ�3�>�̟-��e刺�v*e֪��ݚhV����f�뀪r��8�B#��lW>�)�.�m��2ۈ��I DS Y�k�@E��Y�qK��N��7{]��Q�o�?�]�"zB,]�&_���sx�䯙�gºsI��ϻԕV��p���d�'R�A8��i���qf�C�L j��rK�0�f�4��Y=��'�b��H��^T�peǊ;���m��)�*�e,/don�yQt���iª�� u&�$曨DY¨�@��ո��mbI� �����H�<n�ݫ��[�Pٝ"�Sxx[W�K7�a"D�����J��&�$���h��]����l���KJ��U�N��kt�ڹ�"Y�{#x!�z"� -/� ���F��Tֈ��	_�J��'�
�w������H�|?Zv2�m��ˈN���]X�l
qWl��������C�Kh�\����A��Gd�5U��<2�a�̧f+��:�ؕ�������ޱD"�3~J�C+R	P�,:�0�`�J�l��F��َ�(�����l9I{8�j�t���p�X[^YY�����%ڻw�.2<����f��\#O�������ۏ�~�\�g��� �\�
'�	�a����m��l�X�=�b#�t�7��tۺ�9a)���v;��q��?��3��7�#���A�{,�+t��#}����T�$�s���xL6Wp �T�a}ϛ�{=H����8'�����_���pq�9c�[�,Y�Y!5�|��(��%���]
��3���#�������g+��$���]%B?����l��QK��j����_Gv1�ӫ���߼�\��we>B057�����5�J�B�*́'C8�p����V\�Q���vX�m�/D	+�F)l&�o��kƋ�ѕ0�
g]9~���32�Wpi*?�)���Go�P����`?vW���%�����(�y�x�g����~��^k:a���&�-dx�`�a��O_��)=�Bȃ�J�p�%�O*��9���>&���q�J�K�;�0�q/ݵaZbo�rx, �3LqBIS��������S4�o��FռLB���#��Rr�,Ċ���@�6�LՔ+Z�5.��aPT�[�nQ��#��`~���m���/�9%���6R���e���xcw�(��~؉�D�C�>�����0��p���b��Ȥԇ��u��F�m�����+,v�=�YX^�S�Y�2ED)�a���z�#�Qx��Ed�+<"$fm�9@n�����w�3Bgqj��W�AV%�jxVɲd:�:<y������˵V
k���΍�(A#tVҭ>��~��l/)e��B�\��S��,��7]�lR���3�G�ڼz蠮��h۝���ø���+X7M���䑾G������-���l< �,E,��[2N4�T�� ]���s��j�Ĳ���쑯��Om���g��⺺��RKP����]�B^5�%�oO���׷���>�X�P���4[��MA�0�C)��+=��a?������4RR��ED|�`;O74�&�ly6��0��(��*�����xj�I��,��T��<��7t�m��S4�/��r����S��������L�yv�e��h��y�(x"8x�
�y�6gO�?�G�Q��՞��	���ΐ��-�0r�P�m��t�^�#����p3<XԸ��rJz,�珐F�5��Cә�h���ʣ웙^VJ1�\�
/��_��:�C���2�bǁz��"�_�� 3W�o��.Ǩ�?;-��S�y�doT��!7�Q �W�{T�f�ԇ��J�B5���F|0�UOg!g��*����"!](5��x�f�Ct�&-�~ԇ��*Z�M�ݪ���_K�j9([��)�r96 ?��d�����^	�p����t���YHt���y@�3w�<�3?�y���$��Ysm��M1>���̆+Z�g����H���d�{8D;.�6:� �?���|�ȋ�yY ;�P2_4�?,5�q@$�,r���9s+*���/�hϿI	]�dU�*@E�(]�Z�B���إ+��RO˄��*��4����Ӎjb���Q�6�sk�Ko�키{�,����e�R_����܇/���U���)��͉��m���^j?0<���ĝ1RtDޝ{)�Z�~��0�g�#R%����g-�4��_��=Ѓ�
�=}�ӗ�3���8��2�N�t����<3z#}z����.q�X�Hr�7z�$'�r�K�	Э��0�F7�e���l؅a`��g�7�^���6�a{�md'����.J���%�������q)`;�@ôހI�|Tt��珫�M�D���#��u޷Kl�=�&��$�4��L����q�"��&���zK.Yr��`i��<k\���,��W!�����爓Uv����!FD���`��J���v�\X�
:�2��@�B7�~�	�jh�� 4�֟���=�3�{���������c㪰g�YA�;R+���Ȓ,��V$)ُ�_9i��	��VdF@�s���m��.�nE7��H:*q@�~��ƕn�:�1 �h�Z\��EwK�.I3ȫ�m�������ZGu�#[{�%zO���~��Θ~��Dg[v��bO�JB
����-?v?1c��Δ�v[")`fˋ܌&�&[����h��JBT�Z�B��_])=�n�����,j؄��x��}}�N���S)�X=W�V��Rl��#�V�����E ��ڨS*�U��s�ƺ/!���g�\�VH���*�9�h�u��D��4�e�N
y{r5���1��Y��11���梱~����\|�e��TDh:��e��8?�3y"���ǟ@�
C��c{��x\�h)o�l'`SS7��E�pL���nA��A�8���}1hU;ϡ?IҍhV��<��znr�O�`4��4C�����v���>�!s'�%MjX�Ml?h�ŕ5lۆ���!x������mh��	j�Sdz�ʼ��-b���%�/���8��rr��jc���V�ؠ�E�v���Gd����]���k#���)m�Ҝ��ZBHd��w�)ZF#�gNK; �wq	UC���E��j��z�g��/m�:���R��bݑ�q��S�r�y�o�m	���?�/�.�h/�'�YE���SL&M�
Pd�Z�= E��Sp�įvD4`������hk<~`	 R�V6:Q�.�ƫ}yD�g�b�&�.<���pN����y�qsd)2s7,\L�d����E'�y��Y��J��	\9M��)fh����6��	*&��4�&�?����|$��J��y�ע�O��a��|��!p�H����xq�2;*%�����Q�5X�qK���WR��{j!F������cjMi(�>4*��Q�5��(9N�d`t��膌��y1�
����2ٗ��Fi��џ��?�����<E�^,I��
1�ӯ5��}%LxM�)�b�!S�>iG�����U�g��-w`f���$�f���v9��i���t��H�|,u�2Ǡ%l��6�[�3�}63��Ž=�G ��$�mI�:�,�4�73leg���>>��r�^�Y�c]�1���?�S�����Q�LA��yߠ'���uS" ��@�iM�5������{Z[H"u��cg{�Q����ST"��]�T%�	�7O��#4�YM����p�F,�����p�9rW���2�*h�_y���{D�n\ﴀ��Y�ZJ*xr���o�z|���{R�VUg�����yR� �33%�T��5gz���h�'��c�i���q�A��dsAW��ǆ��Fi�����`�9� ��[=粐�M3Nqv��b��8��\L��^��C�W��F
�~kX��T�?yC1y-�.O��� QJ���>9*}p �}�<�UϚ��>�Ig��ν,��^a>��v�k��hJ�����s���<w^F2Y�鄤������f�:V""I�@��:L�����|�G��R�Uh~���ň�Lm����I��+��	FIoA����0
*>M󄊑`�6̯?s����\�Bz%yk����ԻgB1�ݶ��ȻԖ��j�h��j�0|a'-�ܮTq��.�|��ۧ}��+rQ
�[���`?��{*�k�%c �D�����Px��^��!�r|�
j�P/�[L�kN���o��D{Y;���?з/v�ge�YG�'Z�m5�rږ,�$���L4�������B\*��)
�.�Z�Y��BW���a��`�$��v���Yx�f���� ��l+���9�U��Շ��^^7��DU���"�쟬p�y)|Sv��O��C�$��[���G�_�=�d����Ȃ�
��;��]xLz+�[m�V���^e��0ߔ��Az"�?u̪5����Y4x�a)"(gq�>s�6���눊�D��_���ZTs���qO�����o&�&4���y�Lx�OV�8��3�z­mn�?.F��yXa�.�6A�Y[��3>�2n�OU'�!Y���M�����,&��jv�M6��\�؛H�	��C.21�@�L0���Ar�|:��b%�$.�d99�Mb�;��Ci�'&<-S���В�s�K`>UR������=���#7�E|<d��H�>DW�J_k��EFZ��-֛�
l���]%�*m�Щ[/R?u��Ad.-����>["�����s'&�����E��e�woor/�����Z��!X���]��}�hW���TB8(�y��0�j����(�7�������;"���@�M=�B�8V��<R#K:��|�!��!���᮲��������J9�{��ZW�+�-ﳾ<:{A��b�QG���s��$���}�jk��c���q�O�|� qN���ppy�h���
����z�`7ЃᘂF������VW�^�+���D����=n�W�G�H�n!s�\��� �'�]�k*^��8oO���0.�E	�uκ��s�<�vy�y[e�Gw���|b�l�q+X���Ю�������q��Sn�/�<�F�)������W1y��8��0� &�.����`ꓠ��n]e�Dft8���� �����m�y�W����*�_6��a�c�M�p���bL�-A�@�-IE. �ҽ����Hb���I���w(�co�����H_	�Fh~�ۨ�rm% �����)�� ���=(.��w#|\�﹔�(Sz�a�E���Ĝ���5�C�t����a�H`�B�/�����?��f/�R�q�Y�$�Ƞ����(H��?��Z� 6Q\ �1⃚��~A�I;�~�B_��>�OD�&��M�ć�J���Ӡ�d^�-$D��]ßB�1Il��ɣ�K)1�z��{��S�y��ad<�M_y����\��������C����,�L�(1��-�א.�?��M8T�:ܘ�|�5'��о�e>F�^Y�&��u7�wkA�'�^
����;�/�E�ܻދ-R���*;���Xط�p�џ�=�\\�ܢ`�o��748&�I��L�|Ѻә�����$���<@Gd��������������&1YmYX��!5U+�GQ��Ƒ�;�v�7���V�Bq�{fž;��*>٥�-�:0:x=}ZTZZ1�zK. ��	~5���&̎����U�ҩ�q��3��ʙn�0�d����[buς],U�-� 	�jb��8xX������JӺ(���T����!�œ
�~s]Q�B�Ī���DQ���@��Ȥ��#�'� V�V�=��My7ʚ{\�p+`�c��2BKy�D߇�hA�@�2^��p���/����V�u�%� 0��]	jM�E�Wa��.Xr�G�T�0���&��I�����L��I����g� ~�Ӻ�G*���CL�ަoߺF���sz �`Ql�� G�+�d��x��|DC=����X��zG�I�� �ܝ�\q=� �-��vf	:�U��4�@"'d)D�!�3�plWY�C�Gwe�)�>=�n���p�X,}j��u:�Ѹ����2�M�ڭt��
������>��� (�9�/K�  ��&��=�����i���ߵ�`#�'��E>������5n�8A�Z�Jw���I6��y�a�s5L�������?hm_H��f.Tw�
���kS}�'����0V؜�N6t�!2�\\��l��Ui����T|vi�@H���j�T�c�Ū�G�?ܞ�=�L+��-�Uq/]�Þ̱/�Ǳ�R���B���(=׊-�ո�Zl���a���+y�8����������#[?\��)`c�=�>�:�x��� k}�%�3#iL�H(���\�?h3b��]�+�'kx�W��$Av\�F����	MF7��n��O�|j�����uo_��Ns�mMlUfg��K�f<�x�����u�o
���f������USz_=>�L��G�;5��u-�Jp�O@����5�J$*�O��	.�T?�w7#yV�[�����#�2�^�&OăӪ���H�%6�o�D�.K��jC�N!��O�S݊*攠�
��q���|k{W�#*گN+Y{��g���X�jC1MK�8�H�u#A������I�Cu3��5	ˆ�����!��8���S��N0K���g�����W*Ń�>3qy�Pa&���cz�q(<��s��B�8�/��`�L�\��;��\e��+썘���烄��7�ss�O
�+,~9bŃ�5���؜�\�,Qb�&�Q�c��@��2._�t��}]va���sz��2�ql�D!�f�����~��(0lKS��q�)d�ڕa���Ǭ�t�k���m"rF驑<�"���З5�\��;���t����X��şy�g��{�Y�FUZz�=���(!�^0q�Z�#H=N��ҟ�r�a�لo�{�s]),��.&�N�6��C�Tw6�/F��Q�H@1�J�}�C
�\0��j���6�p��9�~��|}��0���	�g��e#�ly ���W�6�Qxg�l��w�o�!���D�"`;z+�����r�2;j�[�K��s(8�b��t�{���Xo�����^)b�}��	�X�K��U�Y�5�5d�e�P��m�ϻ"FI��wv+_��*�87&X���C寄���u�
.�^� zǦ�2ݿv
��a,���.w�F3��7.�]�E��*Vu��`�ο�g�gAIi]Ė=�9`���*���9�9>���6�u���*���u!�'��)N���jeS؈��,�^�c,��o�r*�W7�P�W���qy�V�?���F����4Pwr_�g$T�9f�-Ki0��Pt�	�������K����v�#��̚��)�������5��c�����F�M�54қ�D����l�s�� �B��\������u�*��������U���ue*e��t~;q�0��쎪ѱ�^TLt�R��h�.�}k�-����I��)VW|���#F9��"0P��EGй����"`�y)�u��:�D�u�`4B��^Γ�)f6�6Z�B/�|Vլ�o�a��S*,(j�Y��kTo�a}�~����j3�Y|��m_<�B�OCT��+ppI䬚�(K��������Rh5���rϔ`lj0|*Y_Nv����8���>et��d���< 2����#���p:drffW�`z�y	"�')�"oz��iy4��mqo3Q
���}Hy��2B�.u9ބL���~�L��q��n���$�tc
�Z,G䱕b�Z�h�|�C��s�������e��&�1`�?yk��5��
�!�z�
Z��2);�ǐrQ�3W�Q���p�
9HB*�@Bt,(~B�v١�;�E����K�
uٷ��Sk-m�[�0!�ؚ�h�DL=Z��a�o��M\D�o���� 鸀��~l��X�O-����94��%��r����/�.V��]%,P��
����C=��S�" ��[%j����$3�8d>�M�C�,\f,��q0`��E�I�+�6β6����,�_?�k֏s����w�W+E\)IYF�+@���=pp���<͎�(���J�R藫{�Y�ݵ޷��Q|�����0=
:pTջ�N�'(`	=ax���]�At|š�!���F�YI����xS��Pd��Ѭ
u\�Q҆���U���K#uOs8&zukM�2��>����̣!��|���cg�߁�7�U�ʸc|�����~f�o���M����{U?/*bI�|tѬ�R�M�ގ3�� 0�F���W����>�4�Q�z�S����y���Ӽ`�:��>9F�u�&�aR��(���ԁ���㔼�H��9K@�<��<뉇��m�~�z'������)$��|0�ߖ�U��C�dgrS'J����C�0�1��)�Y����z���ߪ���;#zv�x?1� ��H��q�2�b��4��P�~/�X�Y�V�m�����D�Ȼ)U�g:JRTM�|�HQ �V��b�z�x� ���T.I#�l|�d��0��h$�������G�{s����ҵ+<��^z/:q���d���I�dn$�{~� {W�Z{��� y�,v|u�]\�ScA}ͣG/���5{�k �+fb\	8}A:&����7����s!M�K�X�7�{nЪM0E�����t	[�x�v߬��N��h�7�`�E����ؼ{\e1D�ڴ�X����XaB�	F��=��K�o�����8�h��'�
�=>��6���p��Lwޛ��tY�T�l�2���0eUD�v�4�u�_[��vv� ���^�N�Ш�i��{A��8_<)rn�M�2�����\͸���M�s>}�ч��^���Y"^H1I��'�3���\ix"�jk������M�jN^Ȣ�c��0�Kd�S׷�_�Vx�k��E\t�Ш���)�m����C���![��u��X�`B��)� ��ەa��t��^F9���!��^�8F����S�
�&���W��t�J�Yc�@�h���ܦ5 ��d������m��\2y�����ʇ
lݠ۞`e�~�rb	4��@E+�L�U�n������!sZyZ�'��J��@��^�Fכ�Ċ���w!��lP-w�`D�b?η���'��:������x�1���Q���߮��`�����|Z�k��F�)���i�oj0S�:��Rډ�զpE���I��swu~%�u�d��:��'��D�_:зlw ��Թ��-�p����R'�PD1�$��I�K��R��0!>7*] ��ci**	x)��\��A8&[ng��j����-k���N�\W���~A�TI��Z�[k�Y�z�q��%��s�.�uN�5�ĀY?���V�n�) ���C�K;�����*7� ��ԭ1�|�6g��h_�EA��p�j5G�&B��cBS�Z��s�m;�&�U��$P��K�o?`��ʰ� Ų`P�5���t����S�H�}34"�R���w	�D�bgt�i^UdS��"�=� $��`N�"758�4��7!��]F�pDC�];�ɦ�,�����*1���~�,��wg��;Pu������?����9LUX��9d�Y�/���pl%((�Wk@B�n�Ŕ�9Pr����1�`{�,�����.�� �ɥ8�O� ��c!�o>H���57�A��/�c�W�r��J=B�U-��=��G��0���Q�#��z��x�A C4�lzx뗢Ed�����I���F�A�HNO(��I}Zv���q���s ?�e��v����f.8+\ah7�HԍM��:��OK&Gk�7W�䔓�`:�T;�H�c�/��:�=�{?4�*�V�A�y��Vg�6���,�r�9���ç] ����R\V�)K�Ja�R�V������&E�K�����*U��ݳR�w���c��)t��s�3�4]�{a�#���$�#�A�[h�L�ȅf8��.�Q��G�a�D�ߋ��2��WJ5n�����Yl4�����ܸ;��r���	��o�&�>�p
pZ���y�.l�}	̠�����������܁~�)y�i�S�6���\!q�eIUy�uL���(P%��IR���;�b�IށSږy�(YPW�OJ�0�����2(��@�1�zj�	�p�TK����J�yd��#w|�3u[6�f��5�4 �*�E�B�����V[U'&�(LIan�N w�z�� 虏�J�]���9{��M�{���&�D�?��Iy��5_Y�-�m��1-�r�J�Z5^A�j�Z�ս#�W�1�!�
5���v+�G�2�l�5p_���d�gRT��9��Χ$�����!�W_��|��JQ�ߙl�� 2zc��X��/Ȃ��xl�"�߿6������}�>�iW9ہo���"����Jխ2>*Tp�/�h�0;�R��d�dR �j�lV��u�0��}t��N �qd�Tl���XB���F�
����s+�U}�5(�N�έ���Za���yHBOi��A]��1��[�X0�h5ig|�eY�Gk𧦎�}��:u0���u{a��r�$x��b�J������F�Z�X��]н�Y�M�H�6Y0VO��8�I&��tb�h����>����߇�XW������#�INt���1���� 6��7��Յw�e����+��F�ߞ�5P:@��*-�����c��ձ'�	�1����#���Hk�s#�p���fo�Y8��/������.�u�U"���^�E�@�x�� ��K�z^h��ϵUΔ����ޯ����ij�?n)u�u�V�4[�ɬ������h��Y4�+�<��rL���B�/5v� ��+���P���D��5�y�@��s�CLY�O�TO����6�������ϰ�b��`(s�L�Ĵm�z9㘇���oaA���b�k*~�[Q�۩�7�7TBD
���A
ڙΨ�i��I&��~3��+��TN����4�˿P���_�����I�@(�#dO��	Co�����i�8�1�g�u�1n~G���^��/_�P��ԪL�[<��]?��&���4�@��J�2h��e����X*":�onh��o��4���k\,a2�l�8(��`�xi����:�Ni�D��ٰ���1$[�"�GК�6(B��Yu�q�0�ӈ��i�dx}��~2羖F��e��Ln*�\	y0������i�
�������@o�
��黶Y=I�:�J�
�O�A�J�t���˨�b��r�<�RG]�1Va�f�d
�P�P��N���H%{?�{�d��C�IDV��և�\�/�zE7_$�eE�fO��ԶY�v@OP6��T.p$�B�(��	�)P��d��.����Z�Q=l����Ҩ�����JQOs}:}�,[U�h�s�O~��$3Ⱥ��-o�"�_�SH����(�Q�p0��\�Cx���Y��������/�`�5���@��=>�BD�kn�U%~ ���b$�	Ϧ.��A�u��T���2X~� �֠�Y�ł���1Vf����k��s�4+:��l�^P�gR�;�]�����T��A-twF��ӯ���{p[N`�z�T��w��H�k��>�flp0�M��Q �ˣ����~�L����.�;r}��G%��>b��x�`fCsL��㫴�C��ݯ��z�*�3(�����Dm��7���.X
"{�E �\
]
_��]6�|w�#0y2���̩iH�ޗ�6�VHV�C-w�k��i㮅v��i�#���E��+9�mi��A��o�{u{
��c�[�&k#��1�E���|ec	!b|�kBq�tM�w�)B>q���8E_��8����+}Z��kH�v���iK��3�ym������<3����A��տ06hy5�F2�n3�ȞF�f)�>�m# WB��T��'6-�����3�������X:Ć���Jci��j��כ�u�8��#��?z.���I��LG�7R<V'��k�~�}}~MJg��x�6�:�����ѷ+�pL�q4�'�m�H��Rڃ6�T����u�1a3�3�ԭ3#b#O�4��)�p����p���Z����B����� �y<���;Dr P�f�dz��%Ɛ�&����,�8��y�3�j�1��$�)��>��_YL$o)������^d����Q��t�����c���y�S��*�PuMs�����*��(!��1;׿��w�V�S�����g`�<�!M�l	��/-W��L&���9�"+�S�����,��K�H��i�_}<��X/o `�6�/��%G;~���GJ�G�;�ف�75�N.������u�� �/+lж�JpEe�8�����8�@:w*�a�:|>���2�3((�\�y%
G�>զ��׸�9�����i:�ШZ��%mhD�ka�ٛ$lXv%ՎQ��t��&��_z�$�i�8��9聫 ���5�����<K��x�C^�y��Ր	)���;���LG@����Y��d��Mlԧ����a��y.����Z�t&�Ñ`��Q'g�nۖQ��>2vz;_��	a�jI��7��B��w� ���'�,aM�X�XK��|����_,S�84a
]�|���v����.;�����b�?�eM=4D�>s*�]!�x��|�9�b'���xB�o,����?��?}�s/��/b7̝�)E��t�E�Ƀ�����Qp]���;�6���QVJh�ە:vFHu�{�Ď7�#(�~u�J�D�H�XT�^Ȑ���Էh�=��I�4,2�g�.D��0"����*Z~+�Ztǳ��Yߔ�a�[�A%��g��d����ടQ�^���̝��Od-,qaP_�P�H��U��&���m�Y=>��VǙJ�0�?��B��ď��ٟ~��:�<<�L�����c�lf�*|��uȦfj���[e��XX��C��N��	����E.�1�/�s��{:I��m��M�ҵ<��>�l�rVW��$tzB�_)n��ڻ}�C��c�w�]���3����� ��~z�)�������ܕ�2�)ĥ_�,�0]y���%��3�1���
�aW,���f7}c`95�/7h�y��9�~9�$�".n��r	Ρ��tPF:=>tى��W��X {�AO��(��U&z�ᙦF���E�[ci|�w�.��� =��݉�ܰ��SAɨPז<�хOEƿ��&�D:R��%����@?�=bM�;C,%�X��aٖ/����h/���S8��1Lب��4U�2��-��钽��n�A�z���":�D�8�c��46��]wj��p��$��(gQ=%r�3z<B����8ŗ��tI�k��㸿a�����a�&�*��n�w��
ruU�u�LHv!��N��N�Uų6��cmv��e���m]H8L�xb8_�I�Xv�fD`�ᕌ����!����|)B����2"�3k��OY=�+���(w,5��y^�T~�l���$�.X��c����s�-�y���Q�����A�Ar�� 1�4�hCG�}h�̰���t�,����Xz6h��b���B�w�*�f�	�p�l�ӖM$�#�j5�+'��!��oK ��`��w6�^�7��i�s���s���]��TH�d`J�����%
�z�{߄}#O+0nq�I9�|F���vh��Ue�|�	NA2�N	���c�/N �j�n��>+�ێ�<�X�;MƏ��&FK���,�_�nM>�u(B?�wF�9�{�3
�x7
�ϰ^k)"&��e�t��2Mjʻr����n��,6�����S��pj���W��oh�=��.��*�!ǃ�$L��-̈́5
�zuP�#�vA
�Kt[�8���kT�Ro
= ľ� 0 J=4�68Lx���0����r�.�2k��?nRR4��^���'{)�m�b�Nps�� �5R5���S�svQR��  �v�J�5]"A٭�쀄C��?l�O�j< 7sx�-Eo�
��K��Q��|��r�/j�1��n����x�P��g���L��C��V�qF}N��5Mz�0�2�sс,��.�T��7�;c_����5j�cODL��v!�uK��������&�$���rR#o�/���'yWӻtu
�#,��	�_�gc����@�_�4��SE�d�!��5.�fJ>��B�i���������+�h%��7�~�LO��MQM�j"���<j��PM���xq�ڞ��=�R������DzH_��1YX���;��`�[ƶ��X`M��j�kiD0�v���1�BْOy�F�J����h}n��E启ቯZo\�@!��y"���IqR[7�+FӸ���� ̘�R��3"�ߺ~xg���� �Y4O占@k��Ɵ�e��	q���2�(�(A�'�ox
��u�H�DQ�tc���oZ�7�b��c�bKd�!$�U	�㵛J���c��3����B���Ct���ܡ]��43-�xPS����")`����3Ʒ����>Gm�a�T�4���I������G%�����F�W78�8H����uJ,���/D�R.B/O���/��ڰ-�5�X�י��b�Xgw���19OFAM���֑ӭ�ΦuGnߎ�S*`٨��
�y�wěܸt�{�����B"��C���Ux�c:�7g��C�zr���\Z�m�/����T���$W�$���u������q�a�����3Av�#zs�ҟgT��T��ͮ��O����P�[�B�h���8^��@����or���_~�̒m�� VaC`�;��ǿ��1�b����]��}�GuaWY�����6�Fx�+�P`/A�{X�.F4Z�Y��+R�K<����D�a׀/��4�bׅ߰}g�&:ɱ��~��SQ����U�E��Y8a�tdkg?����s��M����B$��h�Da0�ь��9� �º%X�K�Q�l!���]�!\�ָ�����u�`P���O'����lЄ��U���׃�_Շq�䯞v���[_ވ�[��)��ҋ��P��A�B3�xya*:V��c�3�؈�U)$T��Blj��H��X�~���}�$
��2ˀ��	z+V) ������1|�6-�%~���Vԃzd���ۑc��:6�♷�N��w'p��?�E������Ik���2�.�Zj�KR �ub_wR����&�3�el��J:�\�a_Q�L��%̚�̵(�Ǵ�Ra���<=���)qZ��E�糄8�ǌ������k�<�r���t�lV4C<C�L6��k�n��2
 I���Cϛ'i���aR�_��eK���:Y���H��ɃEؖdoJ@�d���=3p2 ���5xL���^�@�*naDF9��Q���"���f�e��Z"��==C���0C�39���%�U����2NtM���=$
�p݅�j�����0FKk�`5��f�g�bU�_^�d[7I�Т�s��a-�r���蔋e�o���	]C��1�{��b�,�w�~��V�p�� '�?�L�]i����}� V�.1���!m�Z2_��SM�W�}�SnzA�^j��YJWV�p��Z����UJ��s`@���*|�,\#�F��F
�ցԥ���tDg�=��I����d��T� ��6l�|�|X�?`-�H�$�׀h�:nq���)ƃ�:sq�Jrg�0>��b�N�Y*B��G�V�О����@�=� s0�J�\}������-���`��O%ti֌F��!���F���&N��ęNg@�x�>X���ᕾ�/��(�ަ���DB����E�jQlW`��6"�W�b��7�5�:/H�$�9��__�J)���-�2�f�!�(����D
W�S��6^��]C�$�W�C��W��fY?�z�R?�����\��W½W ���p9�	XQ��{�Tsm��)���v�C���u�Şw^�K�*M�7K75>�����h����L�<�O{љ���ǖvp�v���B�,QƁwF���{���[(,L8������w�A�@�8bR��1���K�7�)!�*���5�H>�����1�0A{��j�d^�
Ź�VS�!���Թe�����V�5jr"U<�g�4.Z��r{���5��ٯ���]t��R�aQI0��BS�P�:��I]dWB4�;2}��ʵ�!�lJF�Fq��Xë�c�o�1H����-������� ��yo����>���FM�R��P�_!?E��Q!,ݚPjP�%d�~b�|�
�&�~]����]��g���k��}rk�Ը���}�U}2�I�8�M��/$��L�-�qc��E���Ix{����
����-�%��y��V��,%�P�`��*�z�偌�]��n���'���2��uR3�o�TQ��S���ڔ��Th�%�.L�����d�Ǜw��+
��H��n�2A�"�]_�e�:�)���d� ���GL�P���թ-���4�j�����$�����`�=�x�9$R�n����xf�y�s�SQ#I�c��br>�!���B�[�􊃂�S��amx��hn�����j��(����[֜`�^��kG<���r���l��+s�b��u�~���8@s���1<4Ѵ۪Z����Ae���z���a�$�+B]���iQ��k� �Ea����1����"=��Gʼá�����u�1"C9�4�q��+�z_a�B�������*�D���<X��Prjn�@�t��N�I�A:GP��|7���ۅ7XU7�������+^�x��N���-��=o�\_�_	iE�0��^���z> ��-�PU�4gpJ�<OhXl�z��:���WwN�&�0N"Bǵ�&@a�AM��[>�ڌ�����~�-�2O�`X�8��N4���H�����gDyy�^C_�N6�(����V�X=��#�$�M�<�/�N�!�	^o\/�4S��h<��a��>ֱ�=6�ۦϖ�JG,���쓰p{N�K֞�`��� ��� �:�qDbYi�}�Y(��s�c�g�S�0��e�D��Ǻ�B��Y����-s ��	�b�������v��%�_�A���� ����5����\��X��Տ~GᧆF��i������r�%���v`3�Q�>��6x�o����}Dr�JGR�@��̿�<�>Mݦt���5Qͨ��b�.0I^!�Tl{VfE�okf���D�i;�Rܟ ���ޣV�,缈�ɿ[�;��T�����������ȝ��%��_��LN:npd�{�NL��E�>IQHDT����;����ƴ�c��/��M���O8�b�Ԡp�6+���ͦ]	���d���eETl~�ok��M��	Q�=��(��J�8��i��M�����e�j�1�wA�ڡ���O����s5�k��Ο��V��������Vig��$�����1K��g)������H��S�>&Q���<���`��	��[��Y_���pK�EnZ @��C�yC��M��~Z�����:顎�Qc��z�>߫ٽ�E�ަ��S���5�-)-���l���27hiK��<���P�*�k]O�2�R��Xռ�,1`���I��䱠�g�_��a�Rŀz�1���S\���x�E�$�pʺ���_%g���Gt	��'��R~9��PW��������;q�<��vS��"��s#�ך����
v,Խ
��Y,j��^���?���8��@�m(��?���nT%�)�駣s�R@z�袣vs:�qL�� �Ϟ�5e͞�ۜ���k��g@�2g�GA��Y�2·Z%n>4�^�<g"و�,�\�s�$$�.@�lk���c~bUD�ל�*_<��1?$��\?g���xG��wӛm��H���H���>��	�Q_���L �ʝ��1�^3g��}�zd奻Wp�]�C��t_�͐?ȵ���tU"�e�
�E��f� �6m�烯���~4�u5�]揄��a��m��g˽�7����T�"�����AO�VQHc��6]�ڲ{�CgR�%�V��?,I�o$k��q�1-�`����t3�����D���j�����懻~���@��.E�j�q�e��b��l��)��#3@�˚��v�*�d�VS-pZy5�j�e+#s|m��c��00��8�X�DU*`$��Lb�8|+�򜃚 	��MA��m�0�� �b�F�vs��-�&��N�_*��6����S��5WL]���;'u�L��W��`(+�p�W� n�ɭ�����_��/vt/ݹ
a�z��AvrՎxi5Є�C��ؼ�bȎM,�P4^42�/
9�[�'=l�8�I܍���/�����_w�{h[^/T�By��渧M:Ji�>lڠz��|�&��}}�g��م�2�T����<�E�Fx�8���Ї��l�]ܡY�s�Q�]y�@���������,�/w9��s�t���8l�������+`�hFF��㬯H.�}=@>ڝ}M�w��� �QN|H�<%q�<0-r�GLlJW_��Фz�([�S�K���.g�e \;T�@ەؤg`�V��O�s{�z���dgJ���x�C���2�q1]`Bb�uxh��Z��:��u�$|�n}��c�t�"��S�� �T�)(|��b#�ɛ���䁃����m�%���ɚY�L�ަ���-��B&_��X◛er8�z����N��v�F �??��1W�R'r���������C˷a4�=����V(&]N��¦ܗg���W�-�v�B�cQ_��zc��sB�Bb���%�� ��R�j��	�3�\)/0n�%jv/���t�q�f"��ք+��U�)ЪLP�P����s�E(����.��j��%�� YX�T"S3d�m���v����
��-Mo=ϷMQgG�K�.BȞ⳨�;q0vA�E������ݼ��S��;��Lc��hj�� )���̇���B_���@�^�0�'��ӻZ���z�~rB��4��%�ϨQ�:h���'���!(E��t^~+�1���՞B�s�T[F�Í�4z~���M�	<����`:pe�pP��
����pDH>�}�s�H�M��&�����h8��a���M���	_���/}�
��y���[���02εRz�3���t��'������׋�l���X���	8�"�Q ��g�ٙDh��_��Ґ���qR{[e �.p���8r�=O�*��6��lK�>����I��\J �p+ �󏳆����=e��w®���T.�9��)���w���.�������ݭ* ��$�*t���c�vp
��-�Y$Pά�ͅ��7>�'W��I�vZ	6�*U`�f	�	�*��sbau��α�uB_��0���Cw �vLLe�_w��ʎW*����A��ŉWq^������9��m�x(�$zkr�K[q<���86=Nh��`�&