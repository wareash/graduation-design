��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jåا{�\�u�?߷�dn@6�zf��r������;,��o+�[��z� XH���Fe>8d-�s�M�u�y�x�'�#����Ih�u��J�)��B7�$=]�~R\_(�c�c����.K߹�)Y��.B���6��y.�����;_��ʢ]���*�p���Q�w}�:�v*a�%�X�B�����v���o6+N^���"�a(��*ĺ���d3׽��T��Y�����Js������p�=�G<G�CP���Ϗ2��O�dƯF��Flf�C�
�m����L �>�7��==��G���,�*�F�����[�[���Ϧ��#'5�aZ����ט�xU�w�b��'����4�c���bI�H��~�m�p�ߢ\���ߖ7�Pk�a��Bh$�q$R��̪�@�P��OW�M���I���K~;�ȾEpu�����c�@��q
ٓ�:�X@HnfaeCp�̩6YR &&n������ϳ�}�VH�G� <M�P*	�*�B�T�_���_��s-\����������)�)��8��^���l]��7��n��t}����0vd��
F$��ΰT�ȜfO7�5�a���C��;�Vf�i�q'u[�д�p�x�G�#vS���!SY�痞��"�h�>6��[YG?�����w�-Ӿ4�xZ��c�,i*�����z?�����h㼯���$��ϒl��H�z������<�ꧩL�B��Z$�@��	pгG7�­{��7��*�(X?nI��M����.਻���VY���ڶ2�����ň19\L��*x��'��3��i	6��f�U���������6<u|�=Fn:��u��S͑ZQکd#��]fnݐ�����>���)���l��L|��)r0����c��=	, ��%��B�ك�8C�lw���0h;7�+�}l�Ų=j�PJ�����G� -��@}���~�8x�*��}����\R�u���It���Q_�$R4��v��P��mxT�wlS<q_���Dv���շ�Dd#��m?����x��1��d�NGlI����ǧ������fA�_ՆH*D�F������mŐ���QR��W%�<�3.7�G']Z���q������ļxL��c�%���p�}?�:� ��F2��Z��l�.�G�8��4{E7�	�'�uաg7�8�klk��TK�v��R7�S�/`���߻�K��M��k�Z�����O�3ѠL��|�V�����}%�<sύ̯&T>��O����X�rH�|0��y�>��&Js:�C^a~p� .� ����Y������8Ͳ�s�79W����8�5����츱૲�&E���{���>�0�¼ª����f1 D�v��S������2rv	� ���@��*=�5�=>�D�4�?܉H��Nk&B��lt�Jq�?�~W���Z��Ru�| @) �tX4�u�x�q�(�/��z d||��mʗfUM�q��阮��#MZd�,Rt��_�6�y�x?�+�j����wr�29�R1*+�lJǜ�����ɘ��@-ŝAc-���J�3���>�.�����XQ�u��ZJ�i�?��iAI^��/b���d�z��Dt8��o�)0�
�|y�]׳,*r�SC~��?O�ՍNU��g�.�||6�V����.��h� j��\�����;{^Vіn-i���{m�9��@�k7�j�Dk֞�6dQ��3'��q9�s���QVH��h<�xr�|(,=��..f-�&���u���ۓb�|4_ݤ�k,��Jc|��J1�$�C����=�QT�nwt)�/d�e�)��c9?4굉�	Nh�꼮�@�ao�´"wލ��չ���Q�x���s����t�	����4�%�VYF�P�����l�>��|,��G��Y�-��]}�A�����G��'��%ݳ�$�ظ�Q�~/��_�v��z�N����WĘ�������J/��&}�	&�2
�Ͷ�;o��)�	���UZ�3�ژެ�-�_�ɭK������U=͌9=Ϝ֐��b�5C���4�\'Jw�,(�5�1�^�H\j�Lb��7+V���cS�PG/�x�Q�"V�u���Ǭ�֢D%&�9A�m�&i�F%G�"��o1z���B���ӎ󂍦:�O�RuU�j��<�i�p������q�j".�y.�$�?[�m�Ǎ���.O ��f�U�!�-��#�C��E$G4L�Y��aSc�е��?ۊW���2��n�yd��ϯG�6�I�� �^Pg[�z^���f��@����M��!�Y����ĵ��',�M��T�L�	a��Dq��"xޒ�Q����TV��:�7��x��+oI�d�utp�k��'��q�hi�3�/�m�*Y��n�T���$�x S�>*��⎽�-4�9\��I��n��4�'�<�{����M���C��Ps�)�ǚ��]=�$��,�kH8QV��ۇ2RQMY�Zz;�&a�t�Z��ĳ�����X2������YO�]ɮ�=���l%3��ⶺ]L=��I�C��.KXC@3��Z�Sz�7��3�6G��k��Հ����I<�x�%i�_�Ujj6Y]$���5��&;�W�G,�-�i?t��t�y��䃖��-�t�Fۑۥ$@��]BI��]�V,^
�Lh����B� H�Ғ�	�IA��'d{y�W�nS�C�P���}�騕��Ф~�5��+���Ƶ
))�E�k:���(ޑ�B��R=(����q��R��
��1��nYt�v�_!;�R��g\sb���+q�7X���J�c^C��6���Z���X�M�R/���회�sA1㫩���n��HNhV�pxWuy4|������՜f�5���n���s��b�S���s��e��}�4Z��n�p�!a,�	!�ҪQf寕~��X�B�����b}��\/:��X���4d��?����!jF�g*����� 1	�	�ܭ�f�d����=6�c�a([�N?ɦ7���4ӈ6>�;�4�oLo��r��A�M=�?�������G�*�@(�Z�a��̛��*x����#�JZJ���z�N�9�����= �S,�bm�`܌ [�|�,����{!����4/h�z�M��N�k�;�4�,=
J)�7�[�_xY���S��X�j�-5r��x���М'�؋F�u2}H�M��/D6�"�Cj�Lz�e|��XdH�_���5v�s��EH5�|�U���A}G�����6�����r��y��u�p
��$َ@�U0ٞ��� ��6�f���$ܝ��F2`A�� �6�����(v:7L�ˢw������2Nf�0S�����I�����>X_~V�������X����67|��R;��!i�p�nY�GbAv��p���}divC(.��Na�1�߸;����)�"���	�G�T�d%yx��,�XY��	��$�Z
1� p�ƛ�t�"�:1��k)i)+�X@�4$�=z�~1����ͪO>�o��$r��cq����ٟ!�E`xV@�ͅ�%Aң4� ���$�_�E9W�%� pgiG�:ى�n�2���`��cF	�.��q�@�Mž�31g�x��yv�3�����B����6�6�(6~z����)�Xn���#�y-��SC�ΓF�	Ā��I��h(U��<W�:��oGA�ֶ �� ,�Bp����q���W�
� ӊ���#������3�-9�%��hZ�[KQ'8�r�Ԥ��N��;Q�V{*�}�I�D ��gAOn��G������^a�����(�e�v����Ȧ����\�"��^U�\(*h��&�kT���Ӡ ����m$&g7+�Hr�=���ib�O��c��m�E�J�x�
�er��R�<�/�QGe�!@
�Y �4�a����Wذ��$CW�?�%���Ɨ��H��ui!ʃ��PST��+���iw�T ��B�����lT!y�˗��ٞ=/L�h�q�*�(�<gKA�w����$ �ܗ�n��T�%��0�(Ǻ4;���扜-���H$�����L��'d�c��|^l~cO��'��--6���c]G?�����������-��X��R�� �ֲֳפ����[ΰ��q-*��8dt��c=�_R �F���kF}H���[D:~n������%.�W��M�e(�'@�����]�C�OR��k!�5X�f�n�����@[jľ������j��3pZ�q�c�-��
e��Yz؎�1?K���UҋE��;-�p�^5��b��8	��C�����0���7EA#PAD��=)�����B�/�h�<��������d�$��DI�27�*��	�w���hLLG��j븆:���?(��}r�"@H}v"/�yR����5�9_�=!8w�Q��m kH�!�U����U��0RzAc�(0{�C�V�5o3�F���]�j�is*qF�ܙY'���:�W^pL������+���_��qP�L�����:�.N���|�5����-���.A�7h'���@|��;��lM�L���$��W�R���;)A���8��̃��B��VIq��31��W8���޵DG��&��{�T����`��O���:z�!1m�n�zH�g�V 5�q>g6��1�=��,RK5@��쥨�n'C�&Y�2��化���ۅ0aj�����l(�Ir��@_���Z��j����#7KB9�͒D�V��2�c:��2��ޛ��s[]d��
f�.��Z3Zb%`�c�)�R�a����]$�}󙺹�_F�)����^r��㭕���:�i���o������5���u�>���a;Ʌ3l��\l�^��U��q�4Vꞟl�̿t /~d3�ǕX+��#m�Lh5|=l�P"n��ƳN=��Q�x���f�h2l�4���,T���ADp�.�5��L�[v�O`*%�٣�������c�55������␡N��`:?�8�kq T��n��M���,d�u�v�|�+oY��N���@h+����ϓ��.�_=���w����%��&~�:�]�0�&t@���ː��Ao��o0���ڴuX�	'�/7,��6�U��������4�����D�40���4_H��-�����<�I�жy����5qu5�{����M)�:1�A�f�퍏��X"`d��ŜI�q_�"_r#h]�a���7��EV[e$���WW��ui���lq	"*�i�4�,f�&Di鄻4:��9�D���*ӎSz�~�)A���?����'��9�P�s0�0wڔ�c��ϥF#�8������6�-��%�(�Nt{w��ݝ�jvI�!���s�Mۇ��?�tzx�(�,�� ���&mI�M^ۙ��;Xy�3{f�U��*9�������[��u@h}�p�$%*i��>z� �,K�y%_���G�����9��Z��~��P�_ȏ-UB4��L����J!@�=7fě�w�ǩ�ےq����Kl`��e�רD 3L��+?�u����C��3���'�%D9V���7
�O[5�Q����e����?��=�9� ����*���ڸ���Z�d�R� �p��N��'��\u_��Ж�8N�{�?���qȐ��%�{�vdцӵ���vU���ٸ�Nо������Za3��ͼ?��D1���<7�w���
i�����(2�RIp���JW�#ֽ�y5fa�3�~%&�o�k����M���##cl��b?ʠ �0�i�jT�,�~�7�X��7H��oe�����Z�bC��Hd��],(yJe�J1�����אX�MǴ��؝���^ k�1��!��zZ�V<���Yߛa~�F5v[;��R�m5�)�ɱ�����m,N����Ѫ��JR�#�H�}8�QǗ'��i��OX�
�]���y�Gj����Ѝ���($0�`����
���-�d�2*a>�s��\ωHA��3����kD� ��K,
Z#<�.�[פ�3�St����I�,�u.�ǹkx��5��&2��$J5�� ����:��\��6�$��j���
f���)A�Þ��1�����v�����Ty�Y��Q�Â�	�^f���b[N�AQ��M�w��`�.i���QŞJ�_��U�1{��E�x?�Ɯ�8����o��6?�I��A��o�XBw������ɭl�^P��f�0I����U�4*��"vD����?�5^��.�������EW�n.�Z���@�6�/^i �(�Q��kJ X����@ӎrw撃�wH��0�D���@��bD�$?��7KQm*��K[i���4�e`E%]~1΁�a�J��Lv/��d��T͔��4���:hds��_yJk�l��I�m�%� F�9k�<n성E�M`�dN���a�	n��;�ōt2x��&���(������ǁ�?��,wUN�X�0K`XlJ�
�q�"@�A�n��)eG$��\��2K�CA%{�:�,��h��9�&�+�b��]� �=aL&[gr�z6%�������)q-�hlE.ʶyF�J��:�^4�]���9��u��y��%��gߡ���	Ws����9ȦN@��{�K
���M�/? �L�;��yH�����V'[���ӳ�4MXjE�f<�
�:؄e
��'|��Vr��N���Ѿ��*�������,`�-�چ���F/eﱺ�#[$lw`|~3-`��<��Os��P��R��3�nrŜ0��MW�9��.��LI8��"�i��e�E&@�(L�X&ԏMW_�lʖ�p_^{����:���L����'����Z^�۷p��v��� X�x-(�9��y��]�} n�9[y��?1鈝����.�R*��U(�䎇��ܣ$��HUԖ�Jm!o�?�sZ��e���R:t�pd-�_�n��FK���ݼ�M3�;��e��tY�B�Y����w13� KQ�R�|��ʾ�J �DAIV�ϕ?�P�Q��PsW_�/'{{ :(�M<Lj2ω|�F��4`�n�/i���~�����)l�G��E��0�ըKj�hC���&RU��M�,��C��Gs����l�A��܋��wl>�	�e�ͩf�v�ʌיek�];�O�����'#�Iv;mk$ Ī�N]�vՃ:��t�����F����O�ٮ-�I�5��. N�_.�Y�Yw���#���d�(rZ�!N�w9�����v��+��	^ |�=y�2'�.��'��<@K���P{oM��:�ҍ�����R���p:D�E���Q�H��]0�(]�{�� ��|W(��k���W�)d�g����Ŗ�?E�j���0����D�C{֤���K_�w�m��k��aN�jlY�m��E�׮l!��W�k�2���25��#u���A$�L�q�e�w�j�[Fw;�M�P'E)�5�&�}�1#��{P ��z$[TJ�,h�r�_�s�#�xi1ōn~i�[���K���Y� ��Z�c~Bް ����	z�+b��������a�<{���80U�e�QX�C�Y:�T���w�T}� ���)���zSY��<�f's��L*�IZ���ҵ�O���ࢁ��^~L)�p�t垂x�d��D��:�SM��/\sBg�i���㗼c5X��r�Ds��z�T;U�";M��h�*��P_����+K3D�|4m�i�,\�4�H��W��B�?�il��	n���"3�2z�R����LФ����S|���4��gp��ߧ,�����Yy���/m�^7���`*:����q=��!�Rа��m�����=�~s �SJ�g��)�Έy��~:�|֐v���B�e��-� l��^����?���c���e��������dUFW
9���&��x����jX�.�El5�-pzp�e��D�
)�{B:C��r�{�8,/�����y�ܾ>�����,(n��G���>���\b�O[2h��}W���mr( 4�V�'��ɼ߰�*:37���5��z��LW����T��(C��/�)��gB:�L|�qpw��덐y�ǢvV1�Y+��*J׍�`��NE��o��qn�?�9���`�	��-d� |��{a�Ҳ���k^�Z�:y�0���ż���r/�7N���.&C$�;
���xs^t�9=���|�OOB���QP�� ��<
�ƌ:��pksF��qH��h��w����~�	,ʱ^Z
��n��ƚ�*�;����UY�z���F����U"O���kk��.���KK������80"�S/�d?ǅ�z�+񷺒6�:�lQ�E�����3��f5���n٦Q��z}+��������)�:I��6M�1+��Y��ki��Cllv\�M�uK/1C��{���ݟ=t��H5+N|[��[$�ǁ�ɜҜ�mDk	�B�O�z}e���\#F�H��@�v�ۂdC�W�Z�����%=���,B�s�+j�ES thd�r�Fk8�B���&��7�+T���[��ps6�_2+]�,���A��	:�f �èfׇ4���k~�6��H�n�L:8��K�SQ{l�e�[	�$�֯�֧�c�>���/���>�{�m�[f��E7�ߪl�t�����M�~�:
��dI\
��!: +�Г*� ?Lb,�p
 F-�v�����q��6!��7O��6��� �X�I�8�����}k�*g�1�鉼���ɘ3x�S3�4�񃤜�j��X�H���:�p�/g5[�)�� �_�W����IB��}.���Hy+�O?d����8�m�w��ag���$���*o�^����&ySk��v�W_V��܉7.R z��yυK�^���'�P6�M �R6�~Yܧܢ�0�@�F��o��$�Ez�n�=��=�f��p�mf��y���5�'{�eA1

����ubn����h�:�|�t��.����O�,��cP�