��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�P�;�{��3�OT����n/\�@���V�F�	G�V��]� z�`t���y[q����a2�,a��rK�&ί�8������s�zW{=��s'^��p��)��d_�y�m�g+L,��l����f	�3v�nҷ�ˊ�a:�?a��D��խ�%��~)c�Ϲ�	����*�IQ�����,U�,M��st8��E�߽>�"�A�V>;2!ٵ��f���<{�x"=�Ce�<�&C}�=�����ݔ��0����Y��y����ΐ��ؙ��U�	ǣ���rQ����
�'v�@���DN���W/�ضW֪9��6ĸ��3��(���[��`�_̠�����6��_���`]�D5�ֵ
8�u�Pp��D�G�&~+- ���������9��Z������$��[��?;����tk¡�[p��#��!�7�0��k{�U�s��E�h �V�������>3BlA<7�\k����`VA�%�Adk`�E�QSa]2��Z�&uO+���PO��i�b��<s�)�2h�!yA�^F�F��Q��\eIV�����"��@��l�Q���b'I0���d�/�V�3O���H\A���g��ޚ˻���2�I}Ԛrlvw�&~����~�{� ����׳�hGU�WX�~�݄��`�����^S
���:e�>8A����'� ��pܽ���߲D�#�˭�����Q���-�K�A�����B��S�'�����zӦ�3�=H��p.�/��)P*ch�P�,�X6+ﳸ%�aO��Sa��ܘ=hr⡍���2��瑲{-+и\��ӄ�|)�<�RK1����(|��K�5���E?>���ζ�/KI^�ˌ�N�	 �ӫ�܌p���D���X&����	Clر�b��r��y���̔4��}�R��;>z�g����K5%x�Z�jBͱ_μ������u���}��f�����O�o�T������v���Z�q�_�au{�*̎�[���eS�pu����n]0�GecmW@̹�wh��5N&�
��4���@aM�y��CZN��ʍD<6׿ҳ"�6�<PP� �_=ow�,l"B&���v;I��GH�Ϛ�T8��Ry�/��M��
�oe:k�<k��A|}�	��g|	ۓ�`�����)8_��&VF6���n��z��ה�\��I��J]q�%d7�(�V�]����s�w6�v'������]��d��*�<z���E���V�N�'�����q�J$3��W[�RAs�v\8������u�I��F^�W�Ņ}0A�'�UaP�*������Hl�G�!��U�Mɨ�d,��m�"V��A����Pe&~xq�EQ�Ӱ�N��n�Ā�u�Z&��̀��Z~�5܄Ҡ0��U�#��X���z�܃����b]���]G��縠|.I�DgBQ�h��r��<�Z�ph%� ��nO�D�Oz��tu�4t#2O�x< �%B��m�wU����3��@p�ʼ/��G<Xʉ��0����PIX ��)����z�%m!�Ծ<,ߍ�S����(��A���R[�ܺʤ�׳�d�\Dp����]���ei��!V�WteK��%g/��sF/ S�&�W\�t,b�������3��i���O������N5.�4)���+��4�-w����|S��P<⏔;�~��=AE���aV�g�{�����C���(�/:g�C�Y��.JOw��Io2�R<D�).��|��a���S���� \�$��(� �c���~�e��)m��g�Q~���~'�8k��v�r�EP�%�!&CVX�,l�� ����`����{�p���JQl��PD3.�2:j!�r�Qd��j	_�� E1�f�����4�ئ[/.���!w�H���$Z.P��kʿ�ܞ�2;����y�O�%����J5$*<�qL5�S��d��_4u	��l����������hКzL��U
�qU����Z�D1���N< Ny�V ��q�2�i�Nv�����p�c�q��F�~~G(1�X3�A�u���oX��ʾ����9Y�Dx&�}�����]���*(��3Pe��l`n�4xE%�6�ߐe����xw:.]7�g����&7��h��VO���Xh��һS�+<Gj<��S>�
����"��5��CgCr����A)�:���`"]~�0MW
���@�g_,�"�p�D��s��q��k�/�JÂP��q��F�+�D �S��}�V�zkP�5�ئ!�SK�Kh� ާY[��J@��u�U�$��O���gw�f�ډ��Mt��Q���ƇH�r{͏#*�E (�,���#>
On/�U�=���)��q�44�:hk�*�a^�Y���㚆��[�غ�L�w��c]��u��aj{�|k_�O� ��X��
��{�q���(W�?�g�$BTtdN�-����z~h�Y�"߱.Q~_T�?��)Q���J>��L�����}9{e���e�d����A��>�$|��s������S�M;�թq��z������t5g3��v�r[meޅ��W_�:	A����$r��C_��߃�ܢ2���ω���p���׏�.�V�e.���y\�,4��⷏�}�gW�S��i^��M��\�Yu�G�̳��L(Z��fZ�Ԗj �>��Bg%�T�G�-WtX�-hJZ@KrX�∭�'[�&��Y��	v���,a[�R��Y���K^-ąS���-�&y�e|싀�'��+JVf*9/�WzT�Ǯ�d�a=�O�x��,F�5�,����"�+�2EI�l��{C��ki��c�%��YT����sL����֠=��4E#�#I��+��&BW��sg�h�cNc;|�B�=���qX����P�hDQ�x�����wZ�7'�J�� �i^?�>5���������N��~��P����s��e��=WW(x��j=|AD)B�O��(��<^7w�)^:/%�@��`��e]n��qU��`
Z�왼Ĥ���Gs��
j�VT�=AE}}�a�x�"��CYI{��w��Ύ�@[	�v�N�R	$;]����'�`,;X�$�Q|t��s��
���o��=H�"�q��0�+�ܼ���c�G�4t�����bԀ�jݹ�7�jޮ�^�M��`��"]w�ԵI�eA�C���qe�nn\�6aQ���0���	�<j��ވ�G�6�yE`0c�}��&(;*��\�]�	��IN�z��i��yP��u? �D�G���-������u�Zn3��xS]�U��5�;P��[����H��YW��k���;7'Zh�
���p������]��U�X�)�N��b��( ���a��ɬz�aP�l�a��eڅ�֦�D��x+�
,�ʂn���@�=�o�-��N�'G6�G���F�MZ������_���i3�i���`�z����>�����9z����d=���*���)6� Vj����̧�qa' p�>����S�:��'�,˱t1��5n�I�F,���+�̟U�K,��/Qp�� ��Wy�wF��x�����.^9��+�O�sn#�a��ɂ��rŤB�䡎i�%�O�y�*��ˤDŰ��|H[���{O.a�\�q@.!k~.N��J�c�����E�z����Md&V����Ӧ.!Wp���'���Z��{����D�;u�}�^�W_�=�`��Mò� ٯ���o��^7F�31�*��_�L{ \��	��x�lK@韞�o�Q��C��>bk��\�%ʻqe�
��s��!boȎ�T=�⟞i��JC���EWE"�G��9"3��c�p��ܥ"��~��돺��3��>�����_��Q�����MԄz���h�����*#��K����t� �k}��J�l�5����s ��|@�p� ��r��,��Y���؄�No�@�0Ѐ�C���	����m ��<��]��9�Ⱥ����P�W�h8��R*`�TƜ�*��"�D�W7�_̿�!���:NE�N�<m}�������H�I�����odD�����e���VƦ�2H�� ��P\}� �i���'���*������W��3m�eO.jmj�?Ȗ+�G�à@!�z���6�E�cR<��A�T�2�1�N��+�t4��'��[J�5�MS�iIP8޴��.�M�:ZqWш3����6@���]��˫m�\��i���Ց[��k�$��k�����hEf9`�(Tp�r��K}���Qs�yìM��Ʌ*���Ʒ�M�re�v����Y:�gz֨j��Pl2��F���<�{��0�D�o��V���1�ߊ?�Ь90f��=S�����#]6�A�֩^n�U]b��� ���m-c�[F��6�+�Z�>����D*�pf^��L}?%:��`(MT��Q������j�7;Z ���-$�+��se��kR��٪y�!(9���D���ml��N�jT�H'�"d�a��i�q��\[X���h�:�}���ЇZ?�Y*�y��᷄���'�A�p���1@�7��D�8(��3؏�(w?�6W�l�oB7�㱗��Y�����81p���/����9��/�B���)��Vq�(z`������CbB���B.3=Z+�̇������5���)AӢ!�R�����?�^��j@�r
��Պms�.!5����>���.+=�2_���w��JE��������U��"�*���M�~C9��6������M%�2�a)�`�$x�5�X�*�#�[�-\�K��e4�?LV�'���I�i��Μ�$�1��2V�w���� �R�Gmh�\�]ˋOl,u������&s��J�qe��m���D�{k�%�ꨘq�G�ᡋ�5rV�8��\j�H��Կ��&��+u�h�v�ž% 3��0U�����	�S>k[�vƺq�.2�˧{k,6�j������yU��K�Gt��k3ݯ�Vʾ��<�*�n��9��ZÛJ�G�rB�����g��W� f�s��@E	�&��o��Y�y�Y�R���U)&t����ܬ.��֛?h�R@C1o�./vf��3�^]�l��9�ӥ~�^q�SE�w�1Q��8�3��r�hت�L�D�zy=V�ݙ7dqp�~�ֵI��)A�hI����v�!�^�mZ�����f�"Ď��ab�Z}��NE��u��?X��Vx[�G�M�a�}��(�����P�Cb��|ޘ��JN��������2�Bx�ă��()z�J�O�D-Z���x8-��}���JhO!�h���}WF��n�����℧��]�����e�(��&&�?_��t�8���T��Mߪ	E/1�[{v���"�w��[<nb5lapN��n�߰�<��g�	��c���X|g�}՘��O���V�b�ߕ]Z/��k4,Z#kd��'p�;= �W�pB�DL��Vf��nGnS�̺X��>�_˞��brL��%�%�Ƶ�_��ܱ���րP=��d�O6�l�+��@��cn�Ѯ���sN5rN�-��@�P���A.W��heV�:a($E�9��������_���8�M!��an$��!`����i!	�����=�{�O1]���׹`��Y����gT���4y �[_S`�$�N;�Q�nTB�|g�Z@:U�\$��	�^�����0""�б���'�@�n�y�����ٗ[-O6W���%AUJ���w�/��CE2̐J/���.��*��v�u��C؍6������`���s�- UW��K����S��N��yۜƬ1*�F���qU�ꅓ�\�9Q�j�1SE�d&�V��U�Ø�����`�7�n�%ȆC��T�6*�tl�˻�mV�/@V�_�;�PGl`��D��m���i&���Ԣfm_����%��{��ܩ�.)�h���q�YWJf�"��"v�u����~w��� �N{�؞|�ߋ-&�an�  Hp�@�}7��>�/<�D5vߑ��ӵ҅����h1��7�@��ᅯa/����lö~5�U��Z�PA�;|U�{���u���0w6��/�Xsᅰ��&v#���tȸ�b�s��z���{��b�Vo=�9��m&U]�\�>�
Wdf�����#U�i7?�>I��8�q�8��fw�0�X��4��W=Wɓ��6�z[�\`H +2n�����S��Ϥ���t�,����m�s��9ٛ/��i0�����&�)^���0آ<��Id/�?O�W�1J����9q��W�j�e����r���~}�l倢��z��T�तz�	`H�x&�u*`U=��	4H�"��j����l���ޥnu���An�t0�o���+�䒧a[�,���Z*<A���퍸�w�(:�������Ϻ7}�}����ů;��ǎGȫ�"��9��X��;e�����&�%�W`d]�<�/����f���p^gm����^G��_�o� Ʊ)�ۛN)˽�-������/�i��]+��[@���-xh��;�����B>z��g��#��rT�|�����H�\q_�Ɛ+�����FBH��`I2���$�Ű�2�6RR����yzKeQD�D �w��J�~J6[�h�{����!���h%���n�0�#l�gߙR�(/�����{#Mb��_���d�����'i~g�1d?g~���^Ҩ�r��MM{ ��&��vn}~l��RWW��).���t��,�V���]o��T�g��Ǚ�N6p�fBb=:OQQ�ׂG�э<�}.[ ��~6><���x���4�ـ�H���@{b�����������%)�l۸��u�7|�c�,�o�m�f/�F
IǸ.5�Z�+Cd�8�(�T��K=����)6s�,���w���܇���ie�����r��.y��]D�3y[q������n���
����3k��������Px��h; n�W[���^�4*/j�*eQy�v�3m0��zA���v���&l��)*������u�خ[T���wF��d>R-�\����L�A񌆃,� K��"u�"	�,c���}�~�ե&�i�x�9K�@�]N�Z���՗�2��}U����#�$�-0�`I�՚��(��>��̈́��*��K���5���0��
Ɲ{x����ܚ�D��2�nh�4`���ssFj�Y�`���_Q��1�^�j:�`kٗ����1�ڔ�[�'��14.HOr/��ނ�n��s=x��'�T&&�3������RA�������'�eu�{�q+�yT��i��v*�IL��1Z��_-`�K��*�r	��Y���P�������=��KOoj���E��Q!ey��N�/5�"G���P@!ްv
S<�|�޴)1�؀eI��Đ��>]�ؚw�
|WЀ�ൌin2[l (=����Q�ӛ�x�[HT{�t��A��H�����l�8�s�ӵ9T⨻m�.�6D)�����lt��rKb�o*X�]���ӆ6A�Bp#ǂ]&�c�8��̖:����Bθзv	�C�����7�0 a��g�L)�z6� mR�]��'�AQؑ�So�^&�R
�A�J��p =>�#���zI|�caI���CϦ�_�P�oc�\|��l\&; ̐@V�Q�*��B�Þ�w���ޱ�ݍ��Z�b��(r>VҖ�M#IH�`&[E�	����J)�Oܾ\Gh�ZE\����掾�y��Y��P��67�+tj�K�b��dl@p�'���y�g�H��.��̊�[y��ƙ�ؿ_|BI,r]��?`O�[X��QM:��M1!|�	�W��c��9{�C'�no�ɼ�o_�1c.1ӄ���ww [�uP��Q0���;]�Eߙ��Td�y�)���hg�Mi��
� ��D��xnV�@ʩ `����d{=d� �������Sfw�)���q4�uG�t�b맮w�3��y*K���(�����WEw%j�D�N���~��� ����������m�HmC�^g2$X��"V7徕��tO��!�0Cn��A��׽*0�P�J���UӇ��Ϊ�f������^�jY�^�PQ�I޽��5����ѿ���^���3�nC��^��(*��_h���_���ZLϏC�0�a���b�������.�ĸ�W�6�><�:�BY@��3k�7(n�Y��w& #�w���&`[RdÜ�mIpޞ ���|�
����ntYq9%����8�J�����b+o�RLrWW�U��G��Y�� 4��&d��&#�,�I���/�N�7�a�eNX���m؇|�J?�PM�u(��ɚk����g	3�ބ�d1���U�0�V[�T,�R�	���`���\-���/kb�0�tm��Pg�E&�t-F,�5�o ���$�M:��6�:�������-1Do�(�����FKZ���Й�[C�l!ᇒ!�u�f{��'���P�%��1�3�4b���V�b�k���f�Wك�jhcy���x`AQY�W9��	��i��o"S�K~sA�^���7J�����+[���E�Ef�p^"��~�|N�����PD�z��������K�J���W��ӽg+c�fr�~mD����'�K��{#��c8������hm��K@~�c7��Y�Pn�BX��"І2G#��#�z��-X������f/�I��Y��h�8�G�"v�g��1zR�=��w��W����	��kԍ�պ.���><��ޫ%l��ɀ�����m{�����>A{གྷQ� ��%M�L5��0%�Ɔ�a�1w�*�RM]���@����3(HI�;4��0���_����K.�����n�3��41���9c�C��K��ͱM!�w\A�z�ޒ�D�:�6*�&�o��K\e�6�sQ�(\ʵ���������ł~��K8��iS�?��t>	Z�!��G�}��U1�$��?�X� �����3_�p��b�ᡙ��;�jA���Fu�ʁ�`VmMH���EY�ԉ��2��;����y���4�e9�Q.�/��g��&c�q�t�gIX-�񌼶�x����;N����x3ȫ���������ńg�j���r6�H����C�`��F[p�G�,�X =�T�1m�1��cէ���R�?'���=�o;sא�g4yY:�v��W=�4������.�S����2)&�oR�`�f7
��ZC�CL�:��h`���[�ǃCU�T�{4�û��͓�d�?!y��i�X� ;�.S/��|Q�H�u'b�_�w{�$�o\�;���B8P&B�~�slL *�3�J�Ik)w�?ن�ӆ�8Tѡ��̣��'����QGq}�3�#�;4�9�/xK�6�3TZ�w��#?Z�c� �!e��G˚C,YĞ��%�z�,������E5O/E'{���+t��1�+L1�Ʋ?�#��k�n��ջ�ҥް�� rL�2�tj$������4�\f��Б�;��� G���3~�3	]z?�����׭z�#B�;�W�Xi�A`��$���)��sh�v
�4�=0�O�g�-E��z�z�ByDJ1�J��"�h��8���ٔ�ˌ���7��
����E�y�Ov��3�d�*��t�y��1X��^]��G��u����2ü3���HtT0��O���Z�8�M��	Z����3�K{s>Sm�U�:�@O�x���Ba ؚ>�#�#�	�=t����x$�rCW�OZ��6�ĦK�6F7ݴLW6��mn� ������2�����3?c��������4h�xc����~��>b*���G���(��iO}�h�W�I���o%�I�
c$��@I��iή���1�A�t�|�qKqE4���,��!��L�o�G]N͟y�]ZT�f���	2�f� (E�zZ<��_�+D���w���o>�C�t�l:��nA�qA�2�(��.$QL�*H��K��P�-�9�Ny��	]�r�Y�=m��	�M��Un��2w@7ل����O>��5��m֘-ۛJz�����\}ǴtF�%��6q��qF5���CZ������^�ܙ�'��f'1""��XɳH@%Ձ�h��X7&ej%e��"ݰN�����Rr<��,��t��OɇY��5U�&�j�p�X��M�y�?�DI&��&�x��D6�Lmzƃ��sQvMZ��r XM�B����^D�4���Y"�����t�����&Q�*�\�d�(Gw�#-���y�{{�Y!c͋�2��ܯ 
�y\KR�ۦ��^��ܹ�"��B�k갌d1~)̧�A�e�Wq��ƥ��]%����}ȫ�V�8�l:j�Q���Ѭ��k�ZO^��\��L�G
�B�@����B�c��RD��=���[��׮�]�y����#�-��G7\l����)��2����s+A֢���z�QK6O�C7H(�#@6)(��QH^�9��_�kl'i�n��qyC�ߣU�W��ٍ����T}���n`]̾�I������A�����ܤ�mj���+ϼ���O����0#�KESq�./��v�Y���+ ���Խ.8����4�z�ycs�I�om
�w�wX�K�9��m��Z�"�c�$q`�x�es/k��N�z��6u�B�5�Hq�K��u�h�<�'vn�HV v�y�'#�^���A�i�$6WTz6e�~k��6�
-�-h�ې�9�.+���
z�$k� D�����Da$M ��V��R~��2�Py�K�M㔺�n�ir�ՂZ���LͿ�Z���B�'t� ���C^�6��t�߹��EՁ��3*j���i�ź�M��������ԯ�E�p��K3a���{ߞt<B�T[�����
]�� ȓ�8th�t<��V���B���T�)R�ר]�ƻ �b2���]��GVY�y��Ľ��
yޏ!�����������6Z���u��O��vՂ�A���H+O�����\NK�9�%|(9��ȗ�\�4�O�O�P��v���fd�#�?r}�x�ɭ?ӗ�!5�ˍ�@X+�<�%U�����<Jկ�P��fZ	>�a�Wo����u�T�_�	��<)g�R
��_SEƪ�WХz>���Cկ-���� ����M�<>���;ǐu+pq=�z�9��e:8i4�{Z9��"Q
�P�B�VC{N��NC�V�������5ܴjQoZ�e��sr�H��73���V�[����-ͳg�tL�5��h�z�Y^*��B�����I�������{��
����U�=��v�э mù'�V܃
��b0-~t��!<����n���c	yt��!���"�ZSлc�r-�����L����|5Վ�h���/WL��"`���O�'��3��������?j���oa�2#ɜN�)�F}�5���-�P��Ǧc�E��f�|��70��/�]=Z��)�aĹ��@��J�M��)��B6�Ѵ�u9�[ܫ]f��v�^ u^�)�|8��O���5�_�����pw
J?P5�u��âr;i�����X8<:�Z�S��cQً����"���Y�ѣ E�$�0>,��kV�Bx��7jŎTޣ��j�_ڱ!�����t8�y���
ևN�O���,�g�\;����V;ș@��rfc�%(��
�	}�~�=a�|0��OB�"��C@���6Y;��[z8��O@2�}a�fWӂE�k�1^�[��ګ�}Q&fq�k丨��<	}��h'��m�)��^�L�M5��i�Dl�Mj,lӍr�E��T���Q��g����LE-s�[�ڨ���9�1IQ!��'�wY�e�c�%���t�О,
�[�G����͋f7s�z���*[��t��f�e��v�z��,��a��o%c�O�M-#�2pD))�?g�֓��֗���	�r��z'V����$�X�Ӧ�!�SO������~A݄
v�z�1:m-���~��3���؀q��}Fp���o��ס������z�i��1��cld�~�!G֥!��C������QurߞtQ���?�y�׸�r�e�#QgU}Κ��M��>���L+	�-X5���|�7H��#c�>W�a�\��]�{�n�U�$�k�&�B&���GoN�C֚���O�my���*~��;<a�DhH�擮U.uxC���^as�N��S W�pu�I��@�U���@�.���o2_�%�+v��j8����{i~-�L`ح��II]]����Bq}w3��_36���Z��@�[��x��x�]ě?ⓔW��d+�#a3������.�T�r[i
]��ն	�jR]w���j$.���Ӽ�~���$V��c�e91Wl�5U��sfJg�!�D���)��=B�7V�r�qc���.>4�M�1�����w�'��Rx�$�<�y�h3IöP���+eq�^�g%���M��4�4��nn�������Yl�-I�ƼH��\*�ù����N
�^y�s�~�~�v�e�Zֹ�<5�kR�Z�O�j���냭'º�q[;����e1X�[B�W� �r�4	�\c[V��Z����;�TBj�QΦ��;U��}��x�=�MC�S�؂�x��"[C��|e$��>wa5�S��
�{~;��/���#m'�^Ơ?��:daj�S2��j�
�x�$,��a	���e�Syk�
��p�Ōr���]<gpc��eJ��c���m�O��b_��0,���G4��x "Z3#g�\�:۬f�N�����7�����\7�j��J���-�)��K��^w�δ/b(Q�Rs9;�w"����}`���iN��R,��)����Kz���
�N��h.�W����y%�%���w ��Vx��yG����R�Τ��2�eqV��"B�FۭIs��0+�">�VR�Y�P���̷��n|SZ�'�� �>r�3>
���_�"]�Hg��}��RkH���\��I}D�>_@�[��Ӗ���5�0��
��1����=�������&5����I�_�7����)���\�I���۵���\x�dſ�`�$V���{���1���Ŵ��~��S/�!k2��!��x.��_Hod�B���ŧH�H��xL��&��<�������G��<�I�y:G�*�m��p
#RǍ�ᇤ֔�j��`�;���k<�R����8��q������Jri�T�D�e��c�!<��Ԡ�����D�)>o}���?}�@�S��q]�/a�b��z&W>���"Kf�s�f�$����b1ݶH��|o�#��ij2RƔ�$z�=�$�L��%f��S:dIex��6ry^}?�C7�!ikG�6�m���͎*z�2���I��=Ap.����޹L�>v��>b5��z�T��}�d�*�\��J���-_�=9E�U:��0����������[�"��U��v��1����!)"�J���A#8p�'��?0~n���FA#Ɖ-��l�e��߽�C�GR���5������%�=�8>(G�t�:���ض�ܨ�z�*�K�׋)���E�Y�3��O���w�bb���R+�nl�k��M�@����*���K��Ĩ��4��ˢ�(�00�4#ܿ��f� C8fb�x� ���R������^GnB�'c�B�X.��헗�{�H7��yB�l�����pކ��tL�T�k�:4p��� �^K��i;�;-f���UQk��$N�7_���jV�/��LQ]�����U�:����-><�r�_�ScQ�u�<K?��I��Z;Gi��U�A�~Т��yq�F0��@2a���V��c*|z����+��ڞE@^�A~A9.
ɉ��2D�.��Y����Fv-w��>�-t��T��#����K[�D�0���ͮSfkGy��li��[W����(�<�����|;��WdERݺ��`BKm,�� �h���L�y��#/��f'�i��	�|�k	�ɑ���}�͍���Cn�9���1e��[&�&��4�8x7�˧�|�k��DB;8��Ѫߦ�2Q��6h�6�ߣ�:��m���F-	�����E�|�lڲ�؇�T+����Ln�:7'�M�1�[����	�s��|sy��NwW���#�'�t��º`lJK�����# ���9CH9yұ�.h #m1�v(��ҩЬ�o�/_W��:A����.Y�)����O&GTy@,�.�p�����t���g���óY��8;7i�8o��:�Kdg^|;���|&0��� ��3a(ݨ�a RL�Y .Ъ��w�K˃d�jBX��;-��lzx�ǜ9e���2k1G�Ģ�{�>?�����0�sٶ���$�D�h�Z�R���a��.�}H��K��]���GCPn �M�L*y�#�)�?�-ܸgğ��PU{��9k�M��]����A�PÓ��:2�g��S�%�����G��)Y���ح8_��s�E��j����E/�X$~�}��-���mM���р;�#7�\!9̣�|.e�N(���U�@��x��}�?/L��'�ha�,>�{f@��dT+ë�m�p	(-�Ì��&�"�W9����a� �g���p���k�Y|�c�!�2V�/RJ*�++��L�eE]\SZNV�������$�(�9c�@�m-����ѿ%����(vO�u�v�M�"�=�o�g9}���M�,�a�[f'�0*�BSlGH]�8C3�[��p��]���TkQ���{�.7+zؔߒҁ��V���i��Nu5 ˜�d�M���퍰=�Yw�4,DV�S~���7S����h�p�jz(E���k^`K�M����?0Cv��&�����9K7Jӣ�ʗ�/��2z$r�z�]��ڷ+���J�ç�g�{(��U��&�[5��HC嗫EQ�~����謂b��H�����\4���2ei���� �t����1�̬5*��\���4ʳ'�Lh���l�v.�wNJy� ���-�d3�'�9B��Vy���Ś��������ojAT�8�BY޲&I�n���O�#p�1[����] ~;{�F��m |�����E!?<���F��N�2�R��IFAf;Z-9΀���ۏ�taQȥd�#�Ee���BS1������D�0L�ۄ�t�ԝ'|.u�#�U�K���;%�H�w�5?[)�
3�!\�x�]{�P�e��ex>X��=K�2TY�yh�h�Uyl�\&!L��}���6��}oP�Z����Et�+ůH+�A����j��B�W�Hн~l6��ո"H2Y�0�Rb���ɍT!�x�N_�'>a�����I8�儸J}���b����6T5�ER��՚{E����V�
����Ժ�D�Cا���&..��o�U��9Sb�̩�%���z a�g�߇�<6�}�ZƧ�8�Zڨ��b���L������:��S��?����CٔU��qb� ��+��cUޗo'�Wg��e�!��`�p�Kʐf�0ӻ��A����g�δ��7���@��v�ٗ���'iݦ��~Y��^�i�A�7�����H�P��E�ǃ,7���d������+8x�@��7��Ċ9��D0�����e��A��d��<ӵ������TG����]$*b
 Z�/�W�0���?�+!��sE,�֟	ᛉ���މ���!��9y�y��w��)���Qgߝ��A:El���*#i
'~([���z1q�i�y8{�w���nvL�u���'c����@8(!��m�@�G����ՙ��:���������m��$V+7
t1�Z���!Yl	��p=��ƿC�T�o�^�U>Y���������,u�l49uK���Ж�����z$��5�ڸ�T�P�\/x"(�mg'��Y��o�+���i:��ߒ����W<��I@�#q�@�``�h���w]+�X�Kͮ������I�J޼�4����%�	{w���M9Y>;�XJz'#Ӥ��+{�-��uy�SЫj�Ѫ��?��ڴ+�S���4�N�c��Q�lq�4��p��yɂ'0O�Y�i
�Y�QV�(���Ϟ��#�*<t|FG��C�6�j�2 ��J�7�9P�<Qi?IXK/$�l�~:�W��zCo���%�J�����7��ܷ
�v�6�r�ɝ���[��-+ˍa'%bRb���	�6�K�2�[�����D���ť��2���OS�5�Dh�KG��0�f'�ի"Ktl�q�}u��0$[��[��n&���:!�?�k_�-�Q�<���#r���e7��␹ր���3�;��&p��#�F���Π�_�<(��@�T�_� 5$�����y�[g�)q�bs�S�cK�y��Ϧ`
��"I��ȵ�;��Sr�!�u�Ν�o�3S+޸��C��~�O���Zϗõ�%.��T��~�I���6Ό3ݶh��1yp!����n��n{���9��?�>C�ز�ΚU<eFLP,>��G�.d�-e�]<�K�NW*����|��������]�H`	(KAy��(2�:�UB��Z��#�����c�d�dDOa���$"�^&���a����ݟ��PEگ}l�I���{-&��&f�>���8|~�T�/w�R�b$��4��g���ѹ@���yr��r�ڷ��j�E�S��q.�����i̛Z������ͳ��ճ���܈�}bpi=�ō�е��j���� 7�<�\�ƘĨ��k_lerV@=D�{����.���2_���	�).�#*� S}�ty�eʮ��NO�
��}�-4��$n�C;�F�)<��������r��:qǺ�e�~�+�|@C�x�{�7�̑�I�X�46�i3X��zvӮ���`�ձ�Z�'�F3��ꦃs�^!�8B⼚�3�Xޟ}�i��:�>�`91%I��5jDl��;
������n;�\t�w?�L
)��j��#l�1�������{;dO���h&9���՜o��J�����Xwlf~a��tGEŷ���^����-��.��pIH�P���,T�Upt�)�{���GZVP������~X�!�Z�ԭ=4���	2��Rr��G���0(������*�p�u����U��+�+�ZN���	��7��)��3G�[��7�����J�c'���|��*�������F��B�.�.�pu�0
�8�$���{2�򩃕4a���M\xE�4�ݐr��B�4�1��lb�6�H�KK+������'�~B������W���]E��~N�����U��g��,�Ƹ>�xq�l�(�sGї`߹�<�N�]H�E��X��+��/���|e�v0H�Z[�.��dS2�:^��<Ug]�4������kE�d������<0��<�3	�!;�|��S� v���G�g�aD�=���EM��^�WFU�V����J�	v�59hHv�S�Q�K�j�_�r��o�,� �j�5��jڳ��p�ɭ;��@�Ȳ��d���!]�& ���;�d=�9���ޥ��(��#芃a������+p��JL_寖�!K��i�fR}�9*�G+C��������>qX�vpj	/�O�eK"m:�S_=�|P�2}<8DXgau��	���C5�qR�K�����{h��ː@t��\�IXx.=�"I4�W~���sb�5��/W4r���;��r��ì��d(��[|��pg�y��=z�w���l$���`�dmV8�Z_���a�9�X�@��=m9c��L��=��mxCa�5�,4��>Ʌ��ѵ+�-6��S�\�0�^b��&��k(�r�܁��]�_�(�} 5q�*��f۾
�ZyT
B�/~�1�ؽ���-9�7\���N�g�� �P�g��/|m)��HG�XVr+���׬)��T�<;~��QGꢤ`��iԴe
e&�&���&�!JF0�Ƕ�4�؋��&�UH�k� �  �Ì2�ƐD�^��C|(0�97�i	L�N �lԏ���� �Q�N�A~����1�}F������^��&]��0f�`2��#����^�SglR�ir1��ޑ�4��M<����8]R:w؆�_��UEc$h�0�>���P��DSb)�R���mPjw��0#WTfo�Ӌ�jj��(v������WW}r����Ŧ��u9�˅z��،�׻݁�[&ixMH�����}
*����L}�����6���s��f��}�D�70:�cQ\%�@�%��5���R��Uf�cqMᗂx��9L�FM	��E�����3��X�ͦ���9�ۤ���3���X��C�l��j[๫ +̀���պD�Zs��?�
in��SB.��� �]%��w5xb�����RP�>�M[UѭB�	9��H�{���9��`��,Q����悳����肆�"�遂� (��D��˘s'K���9����s�*E�eC� ?��n��f���hNd��X�~�^�"7�#d��2rB�.�����L\�eR��S5�������c�|L�Ä��M�Y
�k�{a������Z��]����Pr$��ڠ<Q��w I���V�QI���G�߁·���1�S/H�f�\�:�F����B�bcIņ�{�.��0���A㶬���o+�sO����3�%��J��f�ԪQ;G1��#�J̒v��փ�KW-�����ȋ�L��u�P��W�%��4j(.�R���/�PB�xO�,�wuP��:E5d���+�H�_w.q*QO�Ax"���HU����7%�/��7��X�]��H��
 Z�R���]�Sl�E���[����v��d,�l�� ��?"�0������?�_�KcTcϳP�6�wU����x�����GF����"��6�ҏ^�Orz�I��A�^�=n+�U�u=
1����̆���pY��[��5x���CDԺν�u�}ZTʐ�Y�YR���3®"u�ث�ǠC�:M�?+;�٘���$�㺓�DJ.��d��аTyt�(l��-ߘ=G�r�����%������:��f�AT>;N���qBw�~�2��L������M��~�ڜt�ks���'�q��M�ނ���n�O%H������#1��\s.�o���&a�h��"|�i��$<�jQ5`��Fe�1}�.�cL�Zc�"\n���� opg(��+���k&�^ΗQ��'%4��_�Q�tl��$��W��ʥ�Qዾ��J��ꗸ~\V\C�����RD��<���~�Cj�	�?��.A �NA.j�
5�bu�S�݌�{ޣ���qRN\��i�R)m�� .�J *����8��^H�l.�'����l�� b���I���eI�#{*X[�v5B�A~�B�@ŰWB��mw��v	t����9zC)�w��ڊ��B��	y�K��G�>s9���+©��YH�г�ɶyhg�W�����QJ���
� ���\p���܁�F����E���'�9e�8��E����l$
�����=��84�@��,	c=P��bE� M��0��p!ֆB�V�U�\I�W�H..���2���č ���t���z�����[QScB���5�+�ܟ�(��cBt��z&U �5Xx�o�����z����,n~�h Uq�D]	^��!N�g��s�Ӄl���J
�
�ڒ�!L�-Ih�VO6�[�W���Ú�����@?�`��h�u��Jd� >�)���[�_D�K¶���E��e������$�Jc��e�°"�%	���h�������l
Z;��F�1��Yu������c�,{s�ZF=BwT�/���l�4�X�@�4	��#�#5�m��e��BQ�N9�BXҔ�5��Tt�"�C��-Q���8�$�RS�8�&�X޼d	NV�N����(�P5����y#_�Q�����y�hpnD��nԡ;���b�z0��6������5�_�Z OKT���݊]Du�����NI��+�C.u�W���fwP��!kCy^�����>f��H�֩}C�pX��1�r�^qf�8�f��Ӊ�eᏀ�®���J߬�<LbP�)�
HH>v�g��lu��ʗCZGP���<�W��U��#�ܸlmZ�g���W_o�4%=�K�>�E�E��1^3���]%^)ɪ��V.��9l�o�9�A��{��?�������@+p�� �R"�&�8�@gE����ƫ������1���!���0c
�?��TuF_4��p�#)"�O��e<Y����a�0\�ғ+M=U��4"�X|�A��1q���6<�MН���-#]{Ǯ�)��HU��Z"���=A[-"�t���H����F����y.�Y��WAZ�I�ʉ� 5��e����*�*f�9�X�Tߓ}ߡj�q��o�H�?ӣR�[�B9LKz)�%^��iC��v�}�Us�"���A�A7AȜL��Lf�f!���7�k[��^݄e�F,���&�?��7mbh�鍿T�Ѿw�I����=�W��";�p.+�I��-�Ei�B��Ҟ������l��3��A�]/�%i�)�Js������'�S{��2�����R<����5>�����?@N:~��;�;�_�$�n�q#��8{��]kω�Z�٦�%r���j�8��d��j����2V�9Ba?qI|��'S�&+siW\�	k) �׉+"@b�I�)	��u�M?�{�#b�p��� Up=e�1O�� �[�@%A��'����7E����U��G;'N�Ɨ�>vWU���h�UNA��z��a6(��i�UT<�|����Y�l��<�����_��)P���0�2+�eICxv�mt�~p2ާIV�i�����ГYv�Py9X�����N�A�<�t���4���m�2mC��!,��h&b4t6]S�l�AE���,oR�NZ,��V-NV����������xK��-��>I#�s�`7���婖�z6��zuk��FEK��m��zor����%���pD����7S��w��a�C#���!w��@�_PT� @�Ѽ7�l�l<�x�7D���R������4���"ɾ��y�-\�7�VI-���Έ^�&{�P��4cTTEw�$~�(�<w�m�KU����D�M��
��ih�i�1�h7��f���c���k�8zK��Ey�81�еB�����I�����Hy�ju�N�@돱�I�Kf�Qn�ۏ܊�Ko�]^y���l'KP]��	�D�{�-b�=���e�>���J�f1t���1����
��4}S%��1V��8>�-�-yo�z(��%��^�ע+F�f���1��OCD��� �����Ay{�D��4���Z_}��:�����ԕP�N7g�dϰjQ	�l��V�Y@�T�w��Q��rt�?����q9�E�D���vn��Xkݹ��"_9���vۯ�[)U%z�Y�е_�ڎm�a��KÓ;}��"oZ��:���Z ~�yUv����@����=�iŋj�b���2q�vƠ�����AW����,*�������m�UJ!�HT� B#�$�[>�ʐ;�k�ZL�"U�8�K
���2x��,�C�R� :����Y?����5J���|��������^3r�_}���P��ǽ?Ky{W��9 �^��Dh��~�	��>k���'���_Z/�>��]��T5�<Uz����M�����Q=M&�3�j��,�k�J�̡ظ�ͦ`P@9Lj��%R�C���v�M��ț�$?�~󳋘Erd����)�[5�<`�bCMA3���[�ax�:���Rׇ�2>�GE���J$d{�3�����2)�u!8;�X��Q�OT�d�B����C��CT�ƅ�	����|�ܞ��W���2<M8��i�.����\LI��@�§h�b��f�\�B~�!�mv���`��G�i��)��:D`򣕔�_�yI�E�I�Ќ�Y���GO^�h�;F�N0��m�\:�~�w`�D,�����9��GS�{]��\���J�sA��k���+�/���θv
tSۏ�Ej�-�[�K�}Wam��;k�9p�2BG=V_%Eb�Pҋ(w��ȝ��@�/j����J����@�@����YT�4�@�XkaWЊ@M�1�t�_/b���2�U�PKW��g��?m2y���a���!N�"��9�՛h��X�E�NӋ^�SA�т���:t�σ{{0��j�y��iQ6�G�t�F��2�{Y��:�~��U@ֱed5̤t,�6���A,��A���/�p&�sɼ�B�"N�̉��N�nL'\��l&/�*4��{�P���z8�`K@��"�*O��d2y��4C�0���?�I^�=����|��{WƁ�nF��M�YF��$���#���A>P[�L�1��+s�,Nti��C�&��.�o"��ǆ���y�p~�5Ȟ9m�s�:d�}�@�p[S�V)@���+t)a���0yԉ�B0�Á~� D�~v��q��}b��Zϒ�TH	��7�q�����l
7�<]r>�5� ���bɟ=���j�3)���~�qj�*	R�l�iC�?���L$4���\�d
��;Uj�cp�t�mܸ���3�!o�wk���5��������G�)I @ a:��r<sy_�)��}%���?)Q��!�َ�s�r�j7N�PǓ�Wq��g9(���u[{����B�+d��[rOrj���-ӝFWX���NS�b]Z���<<1e$4C{�y�=�.��dS����cKؖ�2٢mk������ 5)��F�Q�	LmЄ3�g
Z��L�T���d�%O8$�r�^��a(\�ǌ����%�%ѐj�=���y@�|�Q?׊��!5۹���T?o�V�t��t��=3�L���xX�K=S���?+v���&�؇�!W����P��$=�h�M��	��4'��H��gp�B�=f����Y5Cg��d�(���@Vn�KR��練W�<���U��%P?�ѯO>����{ޫU�@��T۪_�sw���}{K��v����v͐^���	Q1��x$&�Զ�F����5樲��o#MP
D�;���X(3D��i0���fK��Wخ����}-{ �t�l�x�����C�v�0�+&��X�H��Δ0q"�2I�e��������ͩӯf!@��v�aP���P����3e�@|��^JU� �H�Ӫq�J�	%�q��s<��A��Ƙ�X��)�.���K�X�)�ڼ��m�u�ĞM�a��	Cfe�js�r��F
I� �w*W��D��)�4�K~�3��d{�\�����W���Y���d"x`
��|�@�n���щ�TPefN	ѳ�p3�zw��	%ҡ��;V����v�cQ0[���)����H4K���$�JW�����!�D>���
���'B�H�ܵV�v�����Rk�UD���!�v����/��_;�k�Nc���1�����7�+�ϙ�H��<�k��h�{�+�0�=��$ٸ�%���X���뱓�5�~��+@7׼�Xat��X�R�r���%���:�dך��M"��<ZX��m�
���O����X���V<j*���_��T��_y_�S����u�I���ӫ�'����VUÓ����(-�xS�&�kp�'S��R���^��0���1 �ORslZ����]��"�7�:����u�O����gg�й����t�x�f �w����<��?X��f�Al3;�&�;��Nb�q��X����4vX/9)I!/pCk������jЄX�s�$�(�c
:�A��d��}��p�Ѻ�CŜt��K0y���X���@o���~��L��!2��V� %���V�N�@`K9䡒���K۟� tD-
g���h��+��d]��
Z�8�L>����&�{����G$��?�S� �g�0$$.G�����A�@f��"*�Y��^�߰���h���I/��.7L�b�pCͶ|�s=�VɛN�\Y�H��R�!���P<E�l�&3E�S���3�9��א�t���<^����|teF��/I�%�r���lj� ����T�l�.=�� w����C0��ʧ!��֔Sb��dUE%���6�A��k̯Y�²?I���$�#Z�)���h��X�f�m7x#�&!,�7j q�����uڄ�kqi =��F�vt��r$k����L�IJ�Rg:^�4/�%t{��&����O��k�.��"e0��U���nw��QXE*�J�$E�.L���dp�h|*��C�).���(��銓�U��YGQG6�5� a�T�$��E���Vp�]$3��}r �;���9@�f~��XĶ���u��S�D��1UJ�v%Yͷ�4�s�A��Lы>avt��z{z�:�� c�T�)+�<X4kdn�g�sS3-�k�DJ��B�������SO�/L�q�Ge7�@I������1�Y�@ՠ�fj�7�.�t�4�K�����8ߨub@ ���!�c�=`����n7�ہ�I\���ؙ����HyŰ��7�p�v���Q��ר�)�0��,��l�8`a�"-��5��2����q9�_��>�܍�wj8���4��O��a�XnC2�(��b�MC�dU�^��y�Q�dΆj�3`���Bk���Y�a�&�1OOD���Vw?7�;�i=��p�󥼋N�H/!�}���߇�L�S;�I�đN��}��-�׊�+��|����ȆMw_	�wd��=�����zw���_�JYc���lc�R|1�X$7���(���!Xt^`��A����D04��o�n&' /i�#ih'�&ϰB�ص� ��᜼����-�YN"��to��r�`8*Wm����������DH�Y�)8��hR����(q$!0��_����rqtXZ�{�깭�Ɵf�����ܽ�N'�e���_�� ��O�4�᳢Ҵ�8휄�k���!t%?�N� 7r&�CGݓw�`�i��e�c�u�@@��4Q�#|�|��t��},1!���c�O(h6����������TTzO�'U��x����e�����R *������pW.Q��3vV k�V A��e�);�
�?��n0߷*ҹyͨmIK��L���p8��/U�i�V;�O_D��V�fǗzM�&�_OV'hr�c%s�l]k�ǁ`s�=2>Y�:��Y�p���VLAַUÕ=ASY�:J�(�̲&��/�v�JL��=��>ѡ�u^��	������/H85f��%/�j�-�P�W>w�5�ٔ��=�#c�5F�l� �9'��%�>(η���|b��r�'�������r�%���f��o��\H�:`8sy����/H~H%�[���R Z�e��8s�ꦹ��cf^�b@I��?3���i��Qs��Y�n��׶ѿ�\���
�Ы���|Q��:�~���zm��u`�{$�JcY[�^9�����Ƿyd�Yf�l��Q+�l[A���CF�˒ֵ�q��HRn)�:��~?#D,,�� �N51�ۨ_��*���b}���eť�pM�<�K�D@h�dD�|�N�/I'��@]�q	"��bN*�I/�v��*�5p��>�!��RX����v<F�`��V0X��dHV�>ҷ�>��k��G\_&܊��/+��5��<Wb�K67z�5�@z�Z����:����#,3�{X���	��L���[�4Ԙ�^fFh�oU�r���6��Ρ;���Q�b��x�x�8�}��@x�D!����ӽ0��˻�<�0o�Σ_��	i��D�4��j�/=�8ˏ=�QsD�%�)�.9���ܚ?���3���a6�d]����N0��S����0#C�y١vwU9 :"� O-�׃nL�u�L�y���s��?�|6I�\FX碽��"���xA&ͬ�,�t&��b#�@���DѨ�0������)�{m-��s�P��k�Mr�R���m��|���9y_K}��/��xA�8�qղ�U	8�].(K5��^����-��w 2Ń�)��]���*h����"����\�&�	����n�m=b��5��$��5;�a*�yҰ�1\�5�o�0�C$E�2Ն�Ęs��M�	���]jF>sk����"Rx�i`ms&�c�Վ��\Sd�5��ʾ0{��s��*M,d���ת�x��.�^��#���q���9�6���M���,�|�Y`��:Ro��y-��І��O�,�T��̡��/h�����z��v�����%.;�w7�rd�q���*���>V��(��)=��H��1`M��S������S��A�
��7	��sB�,�n C��H�8S�R�GY�3�ݿ�wWb�CQ��ś$�?�[�/���^���K�N�x�rIC�I�����~a��Dȷ��޲��n��6v�JL+8���Pd2���%e*��L���x����jp��.���w���#�n�`������	�*�:l����n]YzSi-4	n,$��øWP�!�Ji~�XG�i���>o��N18�����܅ϐLL0ITA��\B�T��6I��4\l�5��|�dy��X�(�J��Hϭ��&�S��E�L
E���$�D��!y[�(�-2yk�6A�J`z��z%ɝ�yI�t�̻ݙ�} ěe }�[L��y�!�3J���(�㒱�Y�"�K��p�<��^���{��D���iA��c�j2���
e
U'�{!ſ~���#S�w�w�=_��/\����K������e�2��I��ǹ��;�^+`^@b����H�J���:���D��T�4Mk�1cG��ѥI��w���f������͛]��Jc��?sE'����7�v9���}	�Wh(�x '��a��e��'cWa�:������-~��2�(�v���n��	0l���_���÷m�5�IR�ӡ�ţD���P|SB�� �r$��O1�Gh��/X��M�.����Afu�F"R@����SmK#���c"`�Z]�xhJ�d��ܤ�"1�R�����\n���oS��z�'��� W�VJD�fN�Ҭ�Ȟ�F�m�I5�F��H���ϳ�xD �����ê��UD8UCc�R^�y�]�f�w��9#�p���� RF-3B����5��ͷGR�v?�X���39�����߀Vl���镪&���`=\u_�6��β�������RI��il�=э�b�<uz?��_i�H	�Z\����BƎ%�2f}Ɖ���*�q?�[ãh@!S�Q�rdx�J��qL�j�wr{� �Rw�?iK����2�%�z0eT�#���A,�Q��׻x�Ł��{kO����^��}���ȃS��c��WD݅��O�͵49,/`�q0FF���*�.�MNB-F�ܬPhf0w������h�5��*%�'l���
n���\�ӂ����J%��尨��f�B��c[��ݤgo&9�������d�?[��$Jo7:�t���W0~��Omu�f��e5����-���&o�B�s�7�pr�)��"�ߡ�4y�^��\�G{h��P�5>�
(f!q����Bcj��@@-�$��2�j���8�g!~�<�lMj��.�l���)Qx���ɻ��S��p�����z�M)�ֈx�x��]��_<t�s�w�(�ɞ�N��1o��.�^�+��' �"��:h�]� ���_�y}ͨO��U���i\+� q���t��dTu�c<#�����WJ�W�c:�uh]�ྖ��n;�tC_�QՓ���F��%Ўɤځ�0�R 6�b�A"X���6�ȩ1K�}
�s��%�Z^�܏n��keƊ�1��ـ �����+���� C����X��K»���Wq���g$�Y�:�|U�c�4n�����*q�$���}�T��
��t@D|�,��go��=�m��G&���`X� ��NoX^�gulhd@{(�(�e�6QoT�©����W.]M΀ӯT�ELC}�{Β�T�0�N���]A&J��yCB-��-x��z��rK���SEh+��� ����{�{�h�$�SAVW���~����E�F/7��d��B��t�`=����#�4\ٹ�;�q�s�%o�ea����!�m�2�+�l;�\�w�TA#vL:�����/�t�R!�k^�]r�=C\=���������+�H�n"a8!��*��_�
���@�m�o�c{ϸni���*�~*~�	�vG��֐$M׵1�nF]RkQU��j���]�>��ؤ	q��tް��ְC�Ǿ2� 9�ʆ��)W�h�Ip..���랩�,B+����@yO,(S�y�Bԅ]�R�m��Z�Ơ ��)���j��͚�'zyi�1�?�q% ��җ'GLկw���l!{� К;\U��o@���o���0�N��+E9�hǒ����?��#�P,��}�떖�͸�o���^�N&v����\���j��3�O��fᤸ�<�n����x��p���ܽ���ʿp�n���q�Z�k+��+��8�N�������i��/R����F�
k�5ٴ[�^V�3b4kF�����<N�e��"�� �7��x��A�?d0���A��y���mw`
���q,���&�k��2:KbT�������ZP�lQ����(�8�͈�FN���ܸ��NV�灑ɝd��&��q8dMyR0s�>O*� 5�bxxX�B_�; 5^N�X��`� :��"�:��P��9����4	,�;��J��z����2ef�ǀЈ�3�E�wG�?�E4���H���TڽZ�ۊ����i14S�z���e�+�c��Z#*���`"�I�{1�S<��SP���U�3��rϡ���w=�d����^�iس]h+Z�/��������L��~���§����b�cXY��m�7;�5�S J4v�H
B1Dh:X�
8�4�ϼ�b�o`*V!�|�~l�X���m�,gPC���6>ٝA<�_;�g$��x��Q�!Qd���N�B_K�)�]K1�qg�w�Q`���,��G?�#�� ��86@��/�!&�_�� �u`q��`rǈ���[�\����i����+��A�U�w��E���'K46��tԊ��E MF]�Oj�u.Ii�_�B��i*{y]���l�G@����)kn(��|�v�g:��+�;�HQ����-��Nlg}�*[M�o��ё��x��$��/ǫ
���2��6��ϖ������,^ڰ�����V
D��;�}ġ]!�
ƢrΙa��OLr�g�aem�7A+�iA2������:\�|e�����rG�*+�p��GR�T*>�;�s�.�E ,�V��sE�Ñ5'$�4Ϻ��8<�R/�l����M~�î��+��ǩ*��m�F|%��=���m�4�: ��Qd��_����Y1n}H���i0���b �7Ҷ�,�:�*�J���3�	��zTp�B�T�#�YF��L|�3��ٰ�+J�n�̕j��04kG��e�{�^D�n�47����5���Thry\zR�	>��� R5QUA09���I���?Q�/�߇+p%U٦�KYJ�q��`�*�?�H#(�|�15��o�_:���
j� �1h��1v[$�"!) 9MB$F;H�j�DWź�3i's&�c�kt:̉�i���1�Q\���Ft�H
sB��#�u�ܴ��v#�,B�2�bN5���!\��H��u�XF#��{��Q^��̛M���HY�ݴ�'\FBc#F��o�ȩ9 ����Ю�����¨��9���� 2�#��&�n�+$(vK%�Gأ���\�iϕ����`*G�!���2�|����J�}O�*��+����D�t1�'C�����%P�Æ֎qC~�E5������>,t������=�^�xJ�ZB�ĥ�!�ڀ�$��&�B���k�D�I"lG��� D�m��7<f_�������k4,bK	u��V{	#̈́�I�!��;<^.M�gk�����۔���c� ED�m����yڃ��1TV�5�<��n'`ׅ��C�����O#a3n��&y?��p/__E�#<b�p섕�/]�	2s����0���L��m}���*l,�� ŗ��W�+W�۬�H$��%�?���&���Y��%�M��!l44x�/`�"m;�֞~0cE�/�0�E�7K<Z>�ɨ ����G���f���Ģ0u���*�»�+j$��k�_c@OXN�/O�q�������c��8k'�.u�#�����uV>�(&T�{��H#c2��_~�la7=�I>��2�f������j�����>�L#�E�T�f ��a�zJ������/n�5{>h�Jlw�xަy�օ����8�+��Ä\�ogB;4�!�9`��>�=!�Fw��s�7��/Q��e��
�EЃʡ�)'vUyR�C/y�ǡ��~%�Щ���;J��l���0��:f�RZɆ($߀%�;e��k�k��"��� '�Å�-ɩ�ۧ ���>	D�,3#��E'I�!����S�����W�v����W�n�)�/�.9��g�I"(n}w���k�!ZI�c��I>�� }b�����sPyܰ}��Cb%��n��i���+�"g�1��[��-�;
j`1��TVN��)���>�WHML�n��m�'�sF���1L}�Q�{����m������$�+�`r^��o��m�!i�y$:1�[rh��r�I;�D�V�����V�������t����R`VCU����y����=`;SWC����4��W�к�Cr���^���5�3sp|�$-���w���R8�I��C���zY����q�`���s?ߐD�YwT�ǔ��uJ(�/��4'7i�,�E��+�Y��k��t$��UOɻ�h�cɎ��y���>��F�s�j&��1g`��w�K�Ĵ/ Nmn��t�jA 7���A�qWt�����<�J�i���e2{�0Ll������3P���|HM��n��e)��Ο�/ih��"���#o�����RTq��N�� ��̝.Nz[o��h�<�6�M� �r)�柶���NK����i"j��m��1��S����ʡ?hŻ�^�3Q�F}������>�w7b�� ��k5����w�В8Ag���-_��m"�ɶB^^� $��=����A�m��2�`�=���aM� �{��H�Dlm"���|�����G�:{�7�k��s�����qם8<�p�k~[���U�+m��6�*>b��҉j[��� e2C�K8�K�'�9��7�/{��s�_��yQuD2��[���=�;
�Ÿ����3��y������M�ڗ�X�i����e��K*�Oe��7Z=�(%��>��7��g��<Tp���ꀅ	��Bփ��86�-KTUI��UAJ���_��/�t��p��X��9 �}�N��v^�B���;���*��K��8BKG�?j8%��&-�Y�5��wD�S��D��14c��G���֔b��1�ۑ�E�yT^+�-/'���6L�Z�`)��[^ߗ����k�]�j�=�Ow2?쁃W�S�h���$D�`@R�Cp�[ͼ��(nו �t�$�	#�@�+ksj9���*�����]c�Ŏ�� �.�2ǔ}����
v�$�C&i�����+ф�VE!q0��Q
}��>�$��!.�3��6�/�X�S�Vv]��DBWmɵB}d���a�	���ؑ��g���$cP�|�lD�5,��ٕF&�u��jA�^7��w�7����y5�4�n�a��� ���Ҝ�L�/�����tc	��S�x�=��ի-��a�ɑ�4Ԟ(�i�������+r�z��q׏���]�"|��`*�է�Jp��n�S�������5��$���29�R,�� �8�q�yn���ҧ�K�!��d��>�A�ZM$����ڳ8�z�ڴzx��/q⭨-����.qX^%�4�k����ad{b���٢8�?�Ԡ��"T潹�.���֖gg\w��	 ���!��h�=gr�@�D ���k�&J�',Y��;�
:��C4k�rx�c$PZ�d���e��Y��uK猅�^�s��p��a	بj��6c��A��%~M/����[
m�w.�T1�Q��.��i�����W0#h¢杶e����	S{�q˒���Q6�ȡ��Dt/�$�!���d����9Ėhv�8f�}0B]�X���b:����q)Sz��T�O�6�������j;��E0r�iCM��i��.NXV�+<����������/�GI��B����\x5�]I�fήvO<�֘/Fb���l��
�)E�1���$�"a�����"BA������=-!x�����X�l��m��؀�v뢕{ߑ�,��입��߂h���=u/���ta�Y��ŕ�/V��?@���}�>��8	$hI���+�(���N�VY)hjz�"�N���R	��`�:U�f�09���gvCf�)�׻1g@��Ӗ ��s52�������m���Uofr/jZ%_bs6�c�~��2����߽��<_v%+�˿��*wWn�D�m[�'LM.숳�B䁾-��y\�3�f�=��:#�7&yb�ӆ�ڤ��~�4E�������컸|���"Ml�iov��7�[�d��9S3'��FF/�շD�l<� i�)9���C��+�>̝�h%�˫�?��i�SJ0�蘿&/Afm�;Sŷ�FkI�)H�K=�V^�g�l�5j��2*R��#'��=uޚ����/��Z1�@c�%BS�5���h�x��:�E�IO�Պ_���z��v���Fq�$��i���kf��~��Q�[? ��T�&Hu�K��p�NM?�(ޑ�d������)��kTS�&鷎c��#��ȿD�H�z$ER<�$���>�����bߏ4g[}�]}6Z�Q/$ηZ<1���3��	��*�}M����6[A]w�ۖ�nm�z�!I�.J��ru���OC�9	��@��-�w�Lj3�W$xϙ��wKYO	&�K�|5j�Xõ�#Q� ٴq����K�h����|���>�S��!�*���j��B}ˡk+�!���8>8�P��U"ޥҶ@Xܖ��:�D[k|:;eU��Zmˋ3
Lȭ���ЛW�@���>�O�=�`U�QCU8�om�60�e1s��� r��#�m�//#��/
�R�/
�*�jу&;�{�������(��x���$�����Ȥc����5X*�t�v}����T��x��$��p*в0��o�hͤ���y���g��2D}�(h���,�{������A�^f�U;����vX���� �+�`�g{yxƴ�(ZS"g	�roW��˺vd����݀�H���S�S��F�4)�jX8���#iux�V@f��U4��"7�l`�T�G��y��2�&�N>�K�4�F�狲i�}�݄@2��\��C���р�Pu`�D�Myv��_X���'��2p>5�4��1q(W���r^��k���җ"[���9�=lć�ڴ���
��׳�nr��A-l\;;��lk��M�Wx%��g��39��R��y�=xA)8Q�ز��Qk�O�i�G�e��9�N��d�+��es%��װ�=�5X��3�0��21ijA�����G��"O����;j��XF�P�"��k9T�Fvħ8R�y������nպ��,���ʲ'Jг咼�)S�C��U�í2]���*S~��g;�K�$��-cÌ �e��zE�� �����<�X�c3�V���Ƀ��S�!ڛI���	6��չ>��P$���1�!�:vtϱ��YČ�c��{c`��c�=��(!9,��#�C�ʑu����r-�Jc⒑W�Kv<z�Q��l�� ẃ��-��pwz�O� �[��)<��Li�ŖǢ�aL�'E�v�=�F7�QWܶ7ޑ���5��9S6������[S���T̲�:T6��?Y�Q�뜑	�%yTBZͣb+ V��܅���w��߿�G	+,$��r��˨O�&����p-F��B�b��Rc[����6�hNJ�{y�Ax��� �r���FO���Z�ݚLn�6,W�C k.�(�`e�zQ�3�Q���6�/d[B�r�Ū���#x�,����x�gg	�Z�,�p��K���~wFk��q
�57�ۡ�r�@m�����$KDqȏ��Dݹ��k�@&��Hޅ��`|`M8@\���|���ﾦ�}��)�7a�<`�K��Q���u���c"o�� �kփ������٥��	:�yBm��Qۘ\���;����X����}Sk�na�=C�RfXL��>$�5ݖ�E����zD�|��Kؿ�� �RWk�o��t~P��VX'b#Z'��dt�f��oC8ۈB�Ɍ����&�5�����_i���,;�ٰ���_�
3�e�^;ةh��E|&U��8u�?#��hq>�%m?Ӕo���k�~��ѓj�ᙛ�d��<�5��P!�BK��,��@7ޏs��R�:��Vᅣ�
����.�M�k��_0:��#�/�<��( �9)x�����!N<�Wr7�-��2B�)���Y�=S��O��ҳ�v�uQ�1-� �����AW��P?*5��� �\*o,���C�B�`��+'��	�* ������[�v����e�ra&��0dmd����E����@h���
��H&y��\)/��J�#�q���<����P��A� οUp
11"iK��8`�'�1�
��z<($��m^���8����IP�0��x�'S���}m=yw���%[i�0�kJJ�B�̈����1H>Kee�$S^;����=���@Xͱ<��Z��sg���r�2����@�(��b1S�S�� ��i@��V(�f-u���mV!����9�����'�BR:A�;��GR���	5D�i~pgj>	���|!�L���i��v5����1�]�&��@YQ+Aݏ4�?$������_���^��QQ�� ?t����?F�#e�����0��i�e�S8�=�u{an��k�حa��d���K��� Z!δ�C��3�)e{��U-0�J�t*|P�������TZ���*./������Kr�'e�^X6���xz�����V�fϖ�ŷ�40�A�f�Ȥ� }$~%�/1�����E�.����#���g������L]~̠D�j�'�_d��}r����`�zH�51�;ܱp?Y�Ôp�0����V+�y�����.̮��9Շ ����̻��7�����1L�gS�k�;��<c&oiҘxד�)~����k��m"n�ul��F��m���e��tk�7�66")JVz�{ZF�G�n7�$�Δ�R.�n�z��M�4�$���g:������<�1��] ׌��е�Px�'�������U�im&��&�e�p����(�b�ڌ8�p-��l���9���I|�A�p�"¡�pd������~V���8K\�������S������;���<��m��J|��;�[/�T�6�+�� �֋o>񧙖�����uZ�;�س�t�Z�����TPs�Y�i`�^�t>.�X��UQ���!�n���^oFZ,�Ȗ���a��G�����u_=B}X{��AJ-���+Q����Xm��� 挋�����S,�d�bД�;}������Q8^�)���X^�@_^�7K��k�n3I��$�ů�YԂ]��Ν���P���5�LVM���d������5OI��b,OBV/>7��ވ
��J6<�2��f���SN��R^��l�.Ǉ�SMn���E�������F�����ĩ�����t�lv�� {;Nu-Q��B�e�	��=���~<v; �0N�;=`[�9W�-=9�zV$�ᓨL[�T�٫���z�l��A{�[�v�5�>@3�h�3�f�}����|�<
��x��I�<�AD˄��w�rvN,
�Mp���(��5�:���P4'�Q&����Y�����(|�F�I�����;̹�����_�&@�̗mD� ��S���|p��f�k������E���x���8���i�2��={�X&E-�;o���[B�eI�w�ӟޮ��^n+�x}ڸ� ˪���ƥv���JCq�`u�\
����6Ws�<��!�(=s"�ӯ�0�s�r�-f����|f����%@�#��D��5H|+�717�Ԙa0�}��S2`����X�Ja��5��?�`����T�h;wm-g�ht�Ze`L-F��@$x�!Ӧ��?�Z&�L�#�~��V�qg�w�YUE�!�tv9����j(�ij����9nV�"�qa�9�f��?vս�j���8�! A��u��I8`/o�|Z �W[��5�nZO�@�G���^㽫���'�f�iTբ5X���HC���Ә���`i>����#i�+��?c Ä�n߸.1���#�?_�p�UO!����l\�b֬2d�h\+�7_�RsTV��x@���.�}�t��K���+�y������ MW�~9;8��z���?��K����_�_��jRn�������<���Y��H�O�BP ��Sd{�wIq����5�����ã=�5�y�5����=	�%��з "/Fb��$S��w�^hc��X�8���0z�e�����9J�W�4u�pcq���+"�m�c=E2��7E4��r�f$�qp͊�*R$*3L���"J!�N��kK��1�d����J�.\r� Y��f�<]��*!��!,h�e���$-P����Sl<!R�����gV���'F�Z7�A2V��jߧ�u��|��<F	�2�n�ޞ�|by=n<I��g�H�Wg�\n��ZKyBe`k�D�D�38��и���?|��$�V"{.����B$���S$<F�S��I��*:?�APq|�E�����5e��Xɫ��<� 5��m>�R9MF-���ݐ,l"��%͵l�#H��9���d��8���:Q~\��Q2�p��j9T_^����'�Y_�'c��M\z*s ��!,�@/�����+��Kx�t�����j�ޞ�VX�h.�l�o0�� /�3�S�%*2��s	锚@i�Q&M��GY�,Fc�B���ԟ>�W��-[t^/ �D��$�ھs�a�q���p81 D\m)��H�C��i�8�5ۚ�v��S��vG��mv�Ҍ���;5��Ղ���6�����~���P@�RB���Euϳ��b�a�!F��c�TR��+6浳/\~V�o��*��ܹc��ѩ�u3׼`�׽1L������Vz!1�Mݚ���܁��TȨ��|Au��.����(�~Щ$��^�S���Ej�6���
R�쳃I��l�B�Y�L8@F�A�)竛]z����oA8 v��������]�KRbL�]��Gy���o�p�/�1_�u��9�hH��5VoV,�2T�q� ����ׁ��B��{k�?����2=Kg��Q��?��5�|���$�y7�b������[��W�4t��7�k��NNw�KO�X�yb���L��>��>�V0�d�]B �~�)��i7Xٲ�Ǜ|
�#N���,�x����)�}s�Y#R��=��]��ـ�X��D���,��AY�/yoIt��Ы�=�y���sA��b ��(`��9�S!�3o!w��ުa����M.[�36�<�k��m��x��xjnԆU��b*��v<;I��I@`D-8�� i|�:���Q����3��m
��'x��r�&.n��I<4��{_ܬ��Y	;/����w�2�X]<�^�_Sq�&�N���w/)������!Ϛ�9�)	o�}���v}=}�Q, gX��w :�@9<9lv��
����@<<���J��_��odTLj�u9Vh�5řN��!����[/�`�r���>_�g���o��9rӸ:=���a�O�)��.!_"����% <C� ��֋T�v�p�����[��R�n��'�����S/w�7���H<ǇT�}J.��jO'���ݔm��0.G:��|M<�c�%O����!�"8߯|;k,����+@8�c���]���j�/��ư_�p A.�DcE����DϬQ���ÜK�A(�CT	P��cA�)1`��	f�H�WO/�����w�<��4Y��QnX#i|>?:��q��M�˛S+����8t$���N���|�a��4v(T�E��K	��m��RC�vTna0-�I �x�F5�!�u�S�/���g�ò1�I�J$��d�����K�,��漧��]KU���'�]ʩ�~���	~�aULt8t� �~���e��7�i�`7qY��(@$2 ��z����8����G�Pe|���Hq9.L�;Aǒ��kM�[�=+g3!�N��$Ѧzf~�jX���Y���c���7q�Dj¶WY��CDgm�3���t�����d;_����/���=�Ѭ�􎶕���V-d���e�Ҭ�i����G�?�:5r[�#�*��S���S����<cp��y��%=!Vgfs ,��|LI��ff��`�F�4^ ې:F�u���/eܝ��a=��Q2��@�;]x�脩ғ�]�dHR<�1狗�ūy;d��$yt��e	`=9ﹽb�d�����;!����F� �հpI{���R�J���MmD���?���S~z����K�G����ڴ�¡�ş&���&Ŕi���)T`�=�ъ2��M�G`���p�{f�υ��T7�R���R�MP�n�F������$9���L� �1���!�$��>&�OFq'Ħ�i��>s��L�"IӨ�W�F<'��"��3g�n�Z~���X�{3HÊL�<�����P��Vūx��s̴�J��&�9��n-���}CsX���<��o"3����ˇ����c�F��>�٬�ˊD�ƶ#����R֨��"�elm��i���;6�1���B?�P�7��;�&�f����x������*ة��ϼ��('ޅ��_;K	�������JP��a����pE��Q?XWh9k2n4�,�)�EtE�i�0����ێc۫f��@*w��a�;8�)�)�|�xn�������!@��ѷ���
�]?w��VJ�!8�Y��󭴉�����x'��E�{�DJ�k���6��i�t�fJ�3�7Z}_;�CT�MT;:DԺ��ߦ��z/�����ڼ�
>R��3���صD��dyZ�s�-$�B��o�Q����b��\�����}�E�*-ZE��q�ޏ�_�e�χ�E�iG��.}Q����ڭ��*hŰ?ɲ�Z�(p
,ޓQ�+60Ѹ`�"^U���W�w�>g���Z����R��nk=٘�nh��֔�������sjPT8ʃ�⬮
C޵�GC)&�����������v�����no��@e�K�֡�⪻�SŽ����|��~hy�N��a�����T8��}[7�n�
ʗ�c5��=�5G~�����Z�e6a�pd�7>x=���K���.�tF#<S=�fFc�C��nt؊���� ؍�b���r���A��a�;��|e�qiqX�\��{��Hs�p��`���������ެ��&�N��:v���}pwOሸ==m~w�����S�F��ݺ�T��f�bk��oc�Gv>A����8DC�����o�6��_�9f�%%�1QK�+�AM�*#G3��1yf�:<�������������x(0��!�Iя��j�Gi��&�VL�qG��;������XH2ˡ��L�Wii<9�����Rp��h��dP#*��>Yo�n�*�O����1��-�Z����vG,P������P�P��=j�
����z���ɂ�P����S��)�i2C�C	J��3�%W!��9l�@H���w��ԏt6O�f�KwD/�;Du���L�o���P�P�mt�n��wȦz��吔����m
�-��p`0���^3TB��Bah�+fݱ���,x�� ��E��W=�ØSo�7��%�[���[%�HyvWj�N��W{���+����*�!�[���4o'���η���-��.��,X�w�oa��SY�3�0��5��,�}t'J��&b����k73�ˁ�-:*�<��h����&�<�͜M�R�zOY�P����vT�E��__}C���j-� �U]�s�=+u��qAе0I.��^�*���� �o�[���6��;�)R�nԑGEJaIfϼ��3u�K�Z�g>E���$}��;����X�˷u8%č?���^3�C"�ǺG��K� ������)3�������K(X]8�/���y����D�|؈���'��_�����������>ٔd�xzQR@��^LR��ϯV�^~�/�@80�tZ���_���$����d)R����[g�?���*b��^
�D
���	9���ԇ�z�sqQ�Ԃ�SS<=X�d⫂\�	ۈQ\�o.!p݅	G�C͸���ԥ��1l���6��[���_W%0
����Qձ�N�a^�[\�׷\�w,%����ir҆��B���r��Qx�A��{�B�^�$[�z�J;n����N�ڣM��\�Wrc�j���$��}�Y�
�e�q�
�b� {&�	sN!��]ı��Lg4t�6����]S���!�=|�.��X��$�f�r�k����jp�-��0� ��7#������A�q .�+��Z�r��7��F�W?��a