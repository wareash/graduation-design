��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�k�۸�m�i(b[�{�㇌�]�i�5'�`;Etg
<������H�W޵α��wԊ�6�a�3� G��λ�:~7 !�v sh��~��P�'|#��x�C�[�~���{-چ��!�:���)�#aE�C�;� ���&�'��c�w|�:�)��$��Sއ�Y�K��N�4uFLN��6n���)G�Kh\��V���IC�"Ჟ�w�߻0w8B��[�vIO�#1IxS[�n���s�h)"��
žgAB �0��wp�L%>�
��ւ#>�4P����6�l⥊�q�ዌ��V1)����yN"��:m%�/&(���`�UcT�XۃUn;xی�
��(uh��=46{eF�ȭplc�qʅԑ߾uo�n$�k��CghI��w�Ĩ9A�,Ub���gBy!ƛ�e����kԇ�$�4�aP��??�N�{V��Iy���#bguګ���</��ɏ�1�3��}�~�Q�*n��p��'�t�6�+ �����a�mo�X���D���|r8S�!;'
�<�w��!d!y�ߑ��#���[�����+�algr_2'����K���j4m]&t���18�q9��'kT�@�9��RR#~�+[��Y��.�����o�,���o`v�zK� ���%��m�M�uN�v�C��Rp��f������D:�[�7M��ETy3܉�z�T���9vT��@([��:����Q���ʱy=����%��(�a�hl��Z��vj�I��%~�:��	�/
���o1�e�����k�5&ꁻ�q���� �Փϳ�Ѱ�2�����E�}U�����`�*}�dVح>����qTL���8,)>��vk�"	�K���
)�}^ࣜ�a������)�Ã��앙�٠����6�Jr%^Ay=�@�L��Jx�����]�v�����c������4��?�^�:D�y <�4`@��zU[�fu>w=Yx��}L��ā�4��k��������r���ٞK�����C��%��F��i������x�*g�^�z�g�7M᧫�X����>�q�t�rt���"�~z��)ш�bmn �g9 �A��cM�9�~x͚�{��ډ%����sxAr�%Bpx���`i�;m��[��o���b�H�]̏�c�d�l�V���G!���=Q�<��o�,�c�{ִ��I)"pd��}�Gv%��[�fyһ����Iۀ��	n�ͣ�d���n��zB��uO��s_��H�;��u��c-��+��S��|�����D%�yzG�r��@��%��:��&�Q��N�i���q�cڜ�8�y��K�k{=4<��Q(	�T�?5��輇,8�C�h�av�.P�lo�e&9��9�����9�O;�LPt��u!7wY>�]�ٙǠ�r���h�矏8ĉ,U2��۫�f����^���!��.u�������^K�P��U �E9be��yJ���id���	ɂ/�R��yy��"��O^�XQ*x���$��Sq~,�;�e\��E�1�S���"���qys+�n��/����`R�C�Li��QpTW���2|u���F�i×
>6E�K�ah��"�hG�AA�ZO$��<}�,�]Ρdy�_ϦR�6��g;�b��%�]B��l�I_�����b��&�q��&9@N���!�i�ˌ��Bs{Rз�k�k�����D%��?�~+���3t�I���Mh_o�ۺ�*��Y�r���2�D�!�/Sۯ�
p{U2�d�R�[d�w���#;#�VQ���}89�\ڬ�D��CC-G]�I�ʧ�i<�h�|J�J���0����î�C�MW������lc3[� ^s޻/�SG�,�r�e�-b�gRU��d�+4Rnn1-�
���<��d|Jb V\L��5ÌH�SƼ�t��Y.�6�*'E����'�w	8PU��N�	$ �P%�7+�=#�a�S|�o�eM�:���4v�q��\U�X��#�zI��$ź�^��'�BS��_{�	��Z*13D4�f"��	�q`�y��1r]�^,�})���T�=��M��<�X�G%#	�[��d���MT7������	H�`m�>�S���������Kb�.-g��G��}�*���0D�"�z|��|0�g"� �d��o\�©I*ޯ���{�t������B>�oss91���sw�FC��_�B��#���Q9E?�3��g���&�'YH[=Hd��
�"[���k���R�~Pݝ�W��w��M�k�L8j[H��ZdS���� �O�G�<[��c�x��̺8]�7�%�������i�����h��Ϯ����(@b�՝iLv����f�����ߘ����R�1������h$���5���K��>�}�I�-S���ts��r�h�0�\R�Y/#H�N��D��p�L����� ������O�NzH����S����<<���M�RƺF0��,{������w�1��c�r����x"�!��Fѳ4D�c� ����p%(㎈Ɖ�.�I����A�����g�q̧M�����z��~k��6��B0�Ɍ��i:H'��͒�c�Qg$g��!����P.��r#�m|� �T�@�f��6�S���+�� �s%!IBe(�Ic����$!viS�(�q��c.�T�~Y���P��݊�n�+BM|W��/{L?�y#���䅣� D��.[,
�2,�Q%e{���	օ�%q��Q�Dk/�#,��WX�$��wBһp��.TE�ݞ��ߢ�TR��d,�
v��'�O���
XWI���c�ě.��Nb�s�f�����Շ`�A	D�Z�7��Y5d2��⠚�;�:�]Q��~XWz�U[�%,&�a6�����Hq����H#E�p΁�ᙙ`P�h�CI����s�J�J��8ڱ�H��T�*����l�k�l}Ĩع/�⣨��[v�}^�zh=٤�.|n�X����6��f���;�8�ڦ�F��2C ��>6<�dO|I��!��4Ϙ�T␄/e.gZ�Wu���G1��F�J[AL�qHg�a�u"��ڝ�6^
w}[ӓw�Кzs��gmQٻa1�]%�Ԍ/N���CK����~��p��sy���j_�f�� ��E�Q���%z�.