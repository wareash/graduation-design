��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�x�W��$�oC�Lw�S
�,h�eԀ)�CQ�_���o�E�'+��l�����qz%�[LըMū��ş��Yz�g�#Vz���E���_�����/��'�w|g>ѐ�=dC6����	NwJ!�
�PΙq����F�<hŚx��#��aT��R��`v����*>wEb�3�4��	ηto��b���RQX_�?+��M���C�ӛ��/�7X�FՃ���W�"�Wa�'_ ���0��a�ߛ߈"�|J�0�g�w���r�~����"0-̦_DoU �0�,���-f��!3�!
\/��M�;�P�[ni�s� R F|�h�[��UtNi�qDۏ����F�N��Q+�9����f&D�����Ш�q�v�.x�a󖷮�]g$�3��|�jWu�m�lB8nB)
�
:�$�y]��Uhֿa�dfp ��:��b��Y�ٻo���i1߾x�B�i��F�"�<0A7l$&������y�Vk����1 F���C�l(*�]}Ԓ�*H��*PPm�>�Z;8~[���Z��{H���^��-���؅��ʫ9di�����K�vk�E�:�3^t3Q1F"�K����>@�H#����]է��檹J���7
W���Z��c��<?��_�[d{�ч��Ϩ�lB�����A�捳�pf4{T\K�:j��.~�����l)��r�^��y�u���s�:$Hh>���	��'xN9��yEySSKҐ*���L+C�4�]j���*�ŒqK�KYeU ��	���X�Y�C�v����]!'XK��q4"�cE>��q9�����2įP����?(�"�{�����,l�{�?l�7�`�@k3L'�����2u[�*R�����V�YN� g��}&U��KG5��[![�@��bH�<	�� "����ޡ)8��0>u�$�U ��F�Zd6��E<b� &S�|�� ��c���i�ڑ�A�h�'��vS��y��+,a�OG7M�ܪ��̮2��x��y:]�/���>5t(m绶Q��
NqC�M����a3�@IHb�).[T�|���L�ʻ@��rk�6��˨�S.xU��x�	��uo��Bf^�-�;��J;���@^��I� L_N���̀v,�Дm����+v�3��s��\�]�(�O��c�6ې���)6y	�8PBSC��HUU=&H�W��cg��P���N$[0�����{h���y:�_���u>��
Ի��<�ɞ����%��[2��zތ�Åh�𓩕}n�3S�i�;�ۙ�RzqO�ADl����ʷ��іO@�ĺ�A
a��w�?fR7������n��cUy���?vԵ\|1�7֩WjM9
��5x�Y6��HZ��.ڤ�<p�pzg�"B��_~\z�c�jA��%gPJ�mC��B�r�=����>��\�~���i��ܼКj���R�9�fx%��b�- �����aV�}��B��Q�w�ˍ'#�ޖퟑb+���9��$@0�������%��AQ�̘���4*X�l��i,�e�>�����f3"Ef�V��n�7��R`� G��\-uvC���M��	��>3���p�X�.�{��G�<?�g	8��c�
)��e�{��cwg�xm`,�)ўR��%���o��LN%��}�f������ĕ?!��y�uD�>;��6~�4�N4�M���V�O[�ݜcm,Ga�*��L/½g]-`�C��镦��rB��M��yޱЌ4�Q3�s�]c,�~F���/
�q�̨w�?��On�x�6���#�;L�D�@�
ܰ.h�Gv�e�;!�>�Ah��CG�@�sq���_���N�ļo�2C��7+e�~�yk��r<��7��"H6l�Ub(�7��W�n�f�Fꋳ���҂d�5��(d���Z�j�����k=��O�%=�q7�A���;9Ưd���ev�x[�5���4��3��,���Y1��E�Bˆ��{6�P�^n����o�����o]X�1G��IB����"���$��������:�$LS��w��{!�{�;h�9A�a��侽I�/*v}��va���V��5�9@~���:��?p����$�Ҹ��>�����`-�mGVH���%�t;gR|�d�e1q��m풑�̬���3�M����m�O�AB�8pM�/��I���0�"�XEH#��N`�?댭
�	�	I���&�vM�����w+���	K��I�P��m��'��F-j������g�[E�Wr/�͓*C��*�vB�z
'��Ղ*v�W�!���
-$�f_>���+u�D�LL�D��"G�Mh|p�EB�4���F�z[�[��2���UQ����f��IB�V��%)ۆC�L�Mw2��$ND��[�[�B�hп�PH���h,�p|��h���T|��w'M\_�>}�uT�ƣh]`g���@]-�O W�عhX*�.Z�t@_N��e\�Ś�ө1�B��(���آ1��G������oBR�������+O"i^h�i�9���W�3u����`�n@�9n~�T���/�b�2`W �Ɠ�\"R��a2O6њ+�Qְ��A����t�]�L{`�h��?�}�F1���"����;y_I��(��Z3^�edd"��@l ��$_n#}໅O����3��S��AŠ � ���er�S;r���I�~1�ȋ�������|R�Zy�4����PM8.uh0pi�G��}̮D�����D�EL@���4�}����ea�AC�6�������Ć��)�Ab��M6��U�&�O05�z�����\����{�W�5A&�Q_�����c�&;����I��^���j�fh�.}��bώU��w��>7�ً�c?�=�g �y���]?;*�|�%�4/����ҝ�XZ6 �@����|�"�B+��c;��:�����dm�,��n�#͓�� ʐmo����v�]��NK<�M2n�Mt!�@���X	ޢXX�����?y��N���4��T�޴Tt�J=��oy�T�l�����a��ɹ��s5�_��A�މ$��._�ʸɖ+#3.��7%V՗�j/����gReࡔ�X������H�/�w~���țFH�1� ��f�V�_)�s��aË�1Y�z�C�u���E<�j��YwUt�]Y%���KicH�IEeZn��Bm�	�=\
���SK��8X��!��Σy�w@�u��+h�ʎ(�:8ȕ݁AV�w���o��Y�e��t����hy@Bh�D�Ls���`H��zt�G��:W����⇐�3%���@��/�a�;�o�2A�O���&�Fl���q�E���"GBvlOm��Y_Qm��6G�r��t�����vH~Ë�E�1�g��nР;d��.�k\�	���ҥXHK��+
\���0BK��R�ܒD�!Rux=�W�q�G�H�_���*�$�lpj0�0�Qᰂ� �40%�V�䢝q���Ujډ��S��or�vn�_�� ��sE�D[��*)3���Z��;�u��}�;��KEv9�������M�2���� c9U��\St�V�U��հ�S3""  �	e�/�d	�+��+�g]��+��#F���wnw5|�Z��f-�rݯ���v�φ�i��1k�j�RS%�.	��I���/��؆Sd�B�.âpu���lhrƪl���CG�ݡ�tt���e�E'���MJ����0���
Ӵ�n����I�F7R&�T���78�Uĺ&}��E}f7c����6_ծJ�n���F����9��6�q�����⇘���%í��*�-���;b�>'��U�@9x��{���X��cu&�.�1�.(�� B� ����r�H�\'V�����a�Qj����n����쎇bAo�uk+T(Jq�-��x���6�-
;\��͐�)L�Xu5���]&(�a���ȫv{�]J95ObY9l1�r���IuL�B�K�����b}��L��&�yΪ��N*Mk�5�D�.���M�&���������52��Y�ޮn�� }��}<����Y�o��X�8�C�>���wE-�j���bɻp��_��%�]���d�$���X��?�L�l|��7��0l}8��yN=�#���N�/D��?�kt ��(_����(LK�V�Vd�����w����j`��f��P{n�x����u��FI�$?gg���<����z�kjkB�z�
Op���KQA��� ���)Ż��@?x���
� &�r7wٜ���D�
4D��A�٨�b�*^q[�����#�BX�R�bn3C��o[��c!�T�Ƕ�P�'�aysӕ1����мG�z$�o�z�aW���t�@'a.��a]9���`���k������O|��o�w ���Vn�X,z��nɬ�����sl˨�����:�*Bܹ��[D�v��Ǘz�����^��?#��׉Bg.f� R��^�f���=�;��EJ�����O��@�T���a��+���q�B�.����su	�g���,�W$�EE���2R����o�� ��~GX҃I3B���P��x�Ri�N���W��Z��Ly���	�Ť�e���v$�Ds戂�J���3
��L
��չ-�����,�����)	>��|C���H��Iܗ���O�qTɲ�&�vqqo���W\L����]��<'�*�
Q��;	E���CL���4!���De+�g��VEf�J|:.�LMB�����k��>�tH���jE����8�_7�7$N]��˖�s�@,ҽ����5�'�A�U�ⅻK�"-̆'#e�/MP�1N{���ϾۑS�N�e�9pkpD1,�����-���qA��i8O�Ղ��B7j M� O�|�uW/���ʪq
%�>]�R�M]�Ri\�o��t��6@+�-B�hmH^r���dW=��|�=Z���Ja�H2C���Q��x`[��G���������ݰuX?	k��EJe��o�p3�z��	�5�Rq�Y������