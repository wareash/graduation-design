��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jåا{�\�u�?߷�dn@6�zf��r������;$VF�w��Tq�����Ʀ��@f�AޭX�tQ�������Wk5)�T����%�h��H���!���|�)���`u�u��X�')�8����!1'����g:1G���H�k}����ˎڀ�e������ O�A�C�����EܛF��g:��*����Ǔ�g��O0F��#g�PL�Q��g����L�K� )�����i�����=�NR�Ͳ]4N���	�)X�uîINA��>m�w��b7��D^�D��:B�N_.��d��U2X���	PtZ��]d��D$cV_"űY՘%<h���@Cj�N�ѮtyO=�)��E���!�Ct�$����k!�y�����j�N�P��`�O9]	��Q�>@x(����x^��%�=F��>w�%���m-��hs�W���f�^y�cS�>N}+�&�)B[8��ͦ1|�DI��hJ-�D�c��l�i���[AK��)`95S/K7=����}��m�̻ח{hU���!m|���l�E\��n��>��� ��{��:��7%W8��C��N�k�3��O/�f�c�׫����R������ ٺ�{Л6ۍj�_�L�4�y�>Ӯ�"h�3�JB���7(���apN_K��lo 8�.�|�mb��wk��� �Q�၈�6��04LϠ�p�M���r�����Eξq�L;�&|��a����ی��|���v��*O"���\7X��B�HRT�����q�� �������H����(���Ec�"��=��s$N�cM�&S�ᓝ�a3� ՝q��}��&��0�+�J/���0|5$ݪ�����5���G��a$�Z��B� �Tr�-F��8�[5iW��&�բ3�-�Գ�W?݈:��d8�㑿}?ue�:�9Q"�B��$+�`�d\#�wS��~+�]&B�)>��2�ށ��h�v�#��}�?E��|7Aྋ:��>�/:;�.���� ����g�K<��vd�t�/��K8�^����=���jfҴ�Z3p�;42{Q��J*j�M,����4eM tb��ՙ[p.�jŜ���v==v۟� KSU�B�f�n|Jj�̺YQ3{����N�2̮&Jy�8���v�����J-�E����o#N�=�ٯ�[�~�Q)}�����=�kqޮ�����2��ƨ)
�+ðɅ_�qP����d՚+Kdi{Z��ʯ5T��	�$PnS��'BQ�u쪪]"0y�<�2��Ŵm�ľ�u�ڪ�D�_B$&�$A�<�
]�\���%��/�Ӟ|���)��V��|	��C���l���Wj�Ŝ����sA?Y^�yZ�Y�F�3F�s7��o�t]��x= �I�4��<�Sv!/6B�����<B�K�����U~�TN@[;.7���(�"��t��T�Н��jU5*:��d�X�US*ƚ���+�w�U���<i�{k����k'��\j�E����ȁ]xl��A��msJT���6�w��Wh[�>|����c�=���@��x�*�;�$'�j��ܾ&�"�.�dcAMO� ���Vf��q'�Z�y�K��䭑�5s�Ւ*�z[_�ڨ�OF�t���^�)ޞpj�����'�u���:��b|�:�zzp�Pf��F3[��a\�ʤ5���H��V<m�b��m�7� tG��|�B߫i�=���"��2�u4赊O���Y��-�z �J���kk�2p�Ȃ)�M��7�7�Z�U��G��;\nO&V"Kr��Z��EA�j��G�B[Hvf=�cl�P�qa����ś/J��]���Eo�����Zԡ�6"���o\B��npm�u����a���'2Y�ٍP�e�O:� ��
*( �!�L�9�6+�*�u�S������u�Q��U��!��f�[d���L!#о �[f�][s�: