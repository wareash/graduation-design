��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|����z=+���v������~hP7�aZ+W���'��T�/��ȣ��<�ǵo<�gX�Ȉ׀B���,�E�Ƶ�,#	h��}4]��>ePVo&�{eA��/*��i6������ߟ�g0����?\����<c"�Et �@r�u$��������b+��f���@����b߮$l�&� �'�"��!�.����k~�S��Q-&�M��ǭØ��1��G �.�<��|�+_��ب���Ւ�m��SJ�m��0�)�K�f���
�8�;��m��_,�a�hB�V�n�a���b��ë�+/�f�;��:�~�����vk��"�iw��w���N����E��z:��IKWR1s��1��zcMY�s�D��z�I|��?���.`7U� �t�Z��׿��"U��>��93���Dm�!J=�U'���"�Ϯ��
9��<[�ar�ҋ6�o��Ja�2�[�3�t�)4;<����H5�SӒ�D�0X�/�f����ՙ�-d�5�����!���zamw�+dF�����	�rR��,��^dի�q�v�����بGҨެ��L�;����H��gC?�((��s�0cD�$�����ϩ\��tD�`/�}K�Y[�� ws*)A����h5�%��!�f�ըPw�PGwb��7Q� ����A-<�k�_�:��� �H��.�e�a���k
�h��К}�N�<�Z�F�`�-`�e�  �Z���;�-�RH(� �`*W$<��M/Ҁ؍�F�Ez}i�J���� ��ux�v8씸T�{��� ���w�$�4iSE6�wC6/#^����S�i�z��D>+�V������G�_ܫ,)��1MA"�]�󞤏�8[��ٿ_�J��d��K����-���9ׯq��Q�B-�F7uXL��8NB�~�Կ�Gw譊�)�����t?(E�2���#ոVAը��'N+�$`��P9��{���3������G���ڤpu���.�x�w�9�,�$q.ò����r0�MbaO2\	�<��F��R��uu����)not#L���<�+OF�_:@s��e�[<�X��^�-��x+؉�����}V=�'f_M(G8���k���2��$Wj	j�Y�;o�a~�����eI����1�Md�3��v��,�GzL�����w����M�lM ���006ۗ)�Gi�^ce{�1�3�8l�$�pf=NN@5"n2|���н���W#Ԇ>�|���M��m���о��+��T��ܬ��\ӭH�xoL�P����3W�$RګӰ�Y�	T�N*ec�/Z���
�.�X����c�V_�W/S���0���\���W7��������WVy+�?�Ma�ܸ�c��e�����AR�|���\�����R�w�ɞa�ǴI�/��2�E���(4��K �ϫo�6��lTHVi�@��'hm6�Yi��zӪ������T������Y�RCf��~�|嫢���Jcư�[	
!VS�3"�[26�]���:"���Cǣ� 5��Ml�3_����L��t��o�*���������ٖ᪩���w�Avp9a���0 {�!1FGvȐ7�ͨ3��N�v(���y��0Ѣ�D�/G��!���) ��u�-��LO
-����6���:��o��byz1��۱K[���^�����ˣj���%��N�25aپ�vy��j�:s/��q7u�B��&�q@"7��i�S!PF�� ��K+*@�\�mPyU��	�������*�Ӄ�����p;0��y��3q��6;�0[*�x�u�3�NH�b̂�
>h��h���3e�[��ob���	0��.I�d�{G}hm�>�A"׵_WX����Es�x���=Yʳ�D�<s}�	9��P�����WoPFv��r�R��ȋ�p��)v�~P���4�;fƋN���J(�7�y��u� 5hY' ��.�u �C�m�ת���=3�_f�� ֔�.%�V�W���)�jxm@M*��zș�h̊�s������ ��p@Q���bNP��uk��UڢC���mJ�-7���g�x���"Ri`�{�566��z��wwEiU���y�j�I��i{�\��WD�mz���̄�����"AJ�1�����9�[=ӿ�=�?{�H.JZ{�`�O���?q�{���S0�;"ޚSJ6��c�b�5�P�@up��呇��s��ӎ5�!���Y�~��5
����b�$���|�O�����K_�5,�.�J�y��m@���s�?�i�Ї%n1G7C����X/������'~|�^+?�i�m��[���`|�b����s����h*�,�CUP���)
I�C�N�����k��5D!���QEޣ��O�]w��r�i�^�F�Yu�ˊ���XO��_��U��D6�z�Mí�[��_-'�C���A�mm� d�ʌF�^�Ag"��i�1�Z�N� v��-g��2���wR�D0Fq|?����5Vf�E3��bq����&����f�:�T��+���ʜ����� 8>��b�d�nX�"�)�Y���aX�G�3wF�A���s)�a���_��=��?Q̉7@�gy�݄��%uB��!:�іTe�?�p���P������s��$�n�t�*��IpC�v��R�b�9[��h��m�M��w��Ԟ*)�䥯b<O���7���z$	_6�&|\��O���5a�����#Bv������jB�׌�UW~�e%�u���"Ҧ�v0�}�g2>�F>fޮg/W ��ʋqB���'�x�i��pU���H���\(}^	�5؄M���r� �#6DBS�LM-��<6�h����A"�aH�B[�;�͆B�&D��x�A�s�=����\g���'�"���oC��p�"��8Xѧ��>��x\]ݳ��)oW�� �͠{j�A��p+]#��/�$9E��hW��k�=2�rd`J�t� � Kװ����Z��v]cQs�<ɵ �ZF�p)� ٺ�|V��1+w�셻�|�G͐K��$���+�17�s��Fݸ�}�8t�$���˸�V騟� �b聡�\�}�*Z�2�0Է��X�k�l�jC$�X�����}t6�Z������8�g�U�\B��Kn�C�8{�=��VD:ֈ��?@����L��%�/�O�x�eݿ�CZ�/{��������r����L2H���,�-��/�Ɉ��ȼ��p��7"��yR���D;ktP���v�/��'�Mqy�'����~���&�<�Z�3��P�	v�3�.�@�DF�j:Z�WX�;�gOA��������|�o�I"����l�ld�6L8�%��`O�KYgDѬb< �$��A����Y�
�P$�@ԐT�?����`�"��D�-�y��BR�������u�@_���3l2�U�pnJ���¦�,�R�𯚇 3�b\j����%t�����p2#��-f0�:C�<�ӵ5 �d �b�i� ��4[��]������z��O��o���
�?\�w��c�����л��q������ XoLj���^
��è�V��2ԏ�(9��0�9�R�*]����