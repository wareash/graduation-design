��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jåا{�\�u�?߷�dn@6�zf��r������;I��BJv2�]�l���n�Pu�оx�&n��?YP&����Ż9�.�+��۳Y<=�q�cބ���%�Z�t�5dz��9�5iN%��k��E��L�
�"��-G�NI�*꥿)3Vn�L���F�����2.�ꮈ��/9a� Ł`��} ڎ�3ג�d�+�ii��'��8a�'�u^'�5ߟ� �-no[�Z�U�\�i�}ʎy�pԦ�{��卾[���WZ#�����3v<�Fl2��1�I�i�d�lǡL��>�W2���mh�헽u�Ɛ�Y+q�j��B��Ҵv0��+(<��N��0��u���$ݾ��RT�VP���q��ʯV�8#�����XY*r�TГ#��Zb�p���.qᑕ���g}��q�崸܃W�SLh��d�3@
R�Z����!o��do�4��?h4wY f��N��7QV�?�Ɛ׻�T��]&��陘%����[p�ꡧ�y����*�DG�9�`��9��?�s����]�|����8���A3��e5B\n��0Cu�M@w�I�O<3˙WcVTf@��/Au�Ç�Ⱥo�P5!G���xG�鄩���]()\�/��J�%�=;���=>RIk��=l�zOWf�Y�ɝ��=�`�M��Y�7�Y*� Cu� ���T��z�<�Ў��Q^�5\�d�����%	 ()�32�X"A��x ��E�X�hH�lZ�� ��+�>����	�F�rQ�,j�S<Vrϰ���8����MU�&L��6���\�����E��"��?��xM�:Ɽ^<TI����H�#��N�����-�'��ͩ0���	�s���E�R��h7H<`��G�[�#߲W���ITtz
Yi+��6�R�nT���ɪ#�Q�C�Z��P�l"u�ZA_w����ȉLQ��% l��{`U�=���V�RV�;�&:�F������� ��ދ�W��a���:�R#pLcG��]m����>ܯإ����8𽹝�l����Ld��'��+G�B����:?�z(�">��K'GO�$�	p$-������$2a.hsߍ���{�{:��}�l�ރ�����&���7���O�����Dc����z۴�퇈.3`!����y�?� 6f�nZ,fUn�  ~�e�O�}�Q�J��W��qO
�;� K�&���/8\��\��b��t"��JLR�븎f�e������d���71��Dܐ���AW���gv�̺XMk�3dh�F�;e�t�W��u� ��#�8��It���q��#�2u���1��@y,�Ȋh���k$�;�S���g~�K������{����{A��^b��D�ΩoF��f�G�S]�fP�h���Ҍ��jZ�	�'�g�t�ޓ�2�s
�RL2�J�I��������V1.������pt�\x9^�vp�p&=?V%̞�e*���`���hG� P��\�|$.��c�u|��׻Űqy︢�����O��(ԍw-�,j	�<3z]�p�@|/��9�Y1q�LO�u�Ż�X�J�-�,F�KZA�F���٤��3Ѝ%&,z�J�')��t{J��Z]M1X,bg`��dΆpE��@N�IY	�r|b���$���^}�ySN����~��@0���	�=IZ�^((<d�U�|�W
W�#J�;�&����}�S���Y��Ijb|#Y�ݯ]q׮��w���p?1�$i`Hsl��.���;�H]�笌��oY������u܉�Bb���^��?O�Ņz43��UcQ�e��Ҫ���
��}[��mϦ�@l@�����r�)f20g�y:���&l��v� 3�ɪ��覕�*��q��YR3h�Hi�TV���7$K��E�}ɨ�P�G~��njP��<	D���͇@?�o
�c��H���!��v�"P�5bP6_��=��y��Ѩȼd�;�ӱ�1>]��w���b;-oi�Г���D��Оz��*�� r&��}[?�bJS��P���!��l��p�}�B�J�o� ��!��y)eu�VK*lv�K!ͫI�i������~P��=v��~����\|������l��|�3�7�k#�\�Z؉���-���
��3��Un���}��n	Z9�1I���h"��o-@"���i�d"�Q�|�� iK�����U�#8JE/��L|xL�تz��zڗ~�B��-*���.��v�M��c��b��?�HK�JQ����b��ni�vި�-ح��1-H����5��d���4 A�{��P�K�C�=�o�A�E�U��բI\K��?���W1w �w\��D}�Ă�Xz�a)��{Jϐ-���<���誆�Z���p�+�8���'c���
8du��"B�˙��	AI�k�>V�R�s�h��l_���Թ�N䤸���8/��SܯX�9��L�-�)����3�j�:�L�l�*9VS����Wj���M&Y�ޢ�������x�!"|���X��T4�_�)+��W�X��w��}���G����H��@�s~�Os���*��i�g|�]R+�
�w��j�s���w�U�WG(0nw<��K?���������q'��a��#c�ԝ u�m��X�{�Mvs��Uk3���u��}��l���q��0�`;EӍf�O�k���Z�+Z"�o�9.]�w��"w4�h"4F̍��Z-C�ٯx��� �R�{3�?=��R��/�C��bBW̾�J���t�V���	��>�Oy� �^Q��,�8@�g��B;�a[�����b0rG�ZM�[��̧�XK����Xk� ��,_�1�|�����pE��H���h�k|ƟG��9�ڱs�e.�,�
U�Z�04�NS��⮢��[na�EJm�Q( ��F�drmE�.�+ߖ�1�]�(&1�>�f/%�g���SK�;�
<P��q	;��	�R��]@7�����=��V��E���7{a�ym��]	�op��:�؏6���g�����f��8�̜@�()�\�ZH.�K�	ًA)�.�w��<��V�=�\"�F�ؖO/y*��\V��(�*Gy�HuLԌ������ �;(n
İ�0͈���@5�33�[;�`���&X"��3m���C� W�9
8t��38 h8��1 ��Z���Q&��[������_TR����GR8�-��� ���i�XGH��y<t�?+L߲P���^�%-�%�������V����xd�d1l�x/Iq\QF�:����G�@�O�Υ���������Ԛ'�vV�zF���
��2��A�&n�����g�R�́��Kj�k����O�H��4Wq�.�9�:U���-�Sb��,O ��"�'��j�C�Dr�^5Ck��g[�����c�p�Na%f;�^Hm.Z��m+T �� ���U�����r>�9r�X�r�n��(����a��������ƫ�^�{���=�3!-u
<Qk`�ry �C�zuz"$�W�Q*Jx�I(B��FJ�ӈ��#���s�y¥��
�����?�f��D $�9������Sd= 퍱g�������l�D:Y�>0�4Ƭ6����{��O�I�#��W��5"H��;������1J�P�I[U�nr\�I#�c@FUCǛmeUI�d �!|B(V9�ٙ� �6���jװ}���a`>W �5Ja��kP�X=�#F�u�J䖳z\��/���@*ޥ�С��K�EG�vL�U�����=�|=K�<v�50��/��k�)�J��PS�~0)�X0h���NG妟�� g�c���iT��s�A��N�{��X-��w�� ;`j��nΕ��(:�#�vmS���f����Y�,��%8� 0"�Ze���Ï5�s$[�0]C�����G+��_�iGm�跮�#IR2˖D�KP)��iud��	��) l ���I��I�E�� ��ֳ���rƹu��ǹ\1arE�e��ArBZ�_j�15тE���Yo���x�u�;�"��䎙d<掠`h����k��W������^{~Y-��u�s�7p.5p�+�H���jލ[�D��Q ���xL+d6�9�lQ�io�tˢ�9�0�z$w�M+�Nz������ T>��rP��Q|�	i��V�#��E�-[����4i�X�2�˾6 n��A�9+�m��t����`��w��̕��<4Ȃ���uK���r/��|TIoɊ,�"E5� ����/��sN�+߮Yg%
t��������(�/n<^���a_k������6h�i�|�}*�!̃;��J��c���
�]�"�f��?���dh��3+]T��)*O�D���
��<����9�G�G.��T����b07���ya�~.�C(�&��̓o no�����~�h0��dUt͜M���;�(���MM���~3gX.��Bx�ֺ�@y������ٖ���kua�h�ɔT��I#\�gQY�ׁm�t���r��	����ҭ	���77�1�Z���/�Uv6.���nb��$	�Ɠu�k�p#5�a����@�N|�*p�@�OD��o>~��A�;�╵*3AG��Q	��ԝG���I��e'Owݢe��s�e��.�Dۤ���|��\>ų�Nݘ$op8�����)�	G{oK�r��T��	2���4a��3��E}�O#5�)Ƚ�;we`uR�K�
}�EMLہ�{�DZ�}nG��t���341Y +�x}����ZP�_>K�޹�ѿ��P �\Kok��KU1K����P�0�Ck����Zr��s��iwo��
zA1��z[�ۈ1F�3��$�y�&I×�0'��h��9_ $��S�;��[OU �x3�a��0�&�׷9U(������*�}PD��|-J����i�����#��*~$��o��\�Y@y@.a4HMH_�/��D̻�:��@��ɒwP��e#����O���=>*�<�@/��x'�����s��uт��n�.qwc���i��+��d;&�x#	-������[}�;t����F�"]F gN���8x7r���7"Q���͍��$��8%�v��6j�6���0N*���O���j������>�i�,[�nɌ�cZ��KM�tg<�L�G��+x�R���J�^�a�Y�����j-�7eMMLK8��vG;g��+{bp#��O-�m�W5<��{�:x|{A�C��T(����K�?�B����_JcJu���θ��b�946�D����_���$֏�@�G��}�p4�eR�_�q��E�\�2�O ��|x}�4��\ݵ۝9Cr����:����T�U ?�?w%��r>!����`�9f(���b�-L��Z��M�A�C�&S�F�
�>~Q����`��oy�0���@���Rgn/p�}�# ��<d��G�^=G�(ur��7&�;>��\�l6A�B=w��yH�\�9�I<�;��T�I|f���k�yPQ���8W��o�E������J,�8�8���E�m�2F����k"a#��)��RL�O�4r�h��3"��aўSDAa��Y,��)609BN�⮎'��\�;F��-�eU���Q�ܭ�%�����s���ʍP�w��.ǣ�
&/ :%���϶�j<X-�P./XDJ ���v��0Ѻ��C���J�_`�O�(�$�E��b��2�U4���7Z���qڱNx���X��끆cOH�+q���{�>������D����M�S��VU�����/o�1��T���5�mr��������=�ϻ�e��i=��x�4�G$iۈNJ9I¥V޴��LM�|��f�(�S�9�DV�%�� 3J�A�F���_a#�����Lr��K�)��yL >��&��b��b7e�X�C8}g�����92l���~��dA~|B'�|J7ۘ�<�[�H���^���=Â��g��y�{F9��4W�$���׻!�o�:��r��H�o J�� B銃���y�����]��ݵ����hם�c�y�R
>$��Q,�e�l���H]��w����v��<��G�FHg 6MӨ)ΓZ�\1������pw�K�-H��;��z?��/<��X�:3���=@]��_g[>�o�Q͗@�rT~�����R޶����	�X��Fo���5ˑ������e���M5�J2��a����B�\��?z�<���V����w��VI��M��Yw�i�x�M�R*�@<�[t�]�Uh��KJ�E,�]Ѝ����[8_AwTK�)�m�ė)�s��z��g�;v6��V"v�l�!=��!%Q�h��pr�(/%�+������L�52}K�1`�#��_.q �y�B�	"����3Y�NTȼh���7E��B��P񓓙l�J`
w���޻�}Q8�ꋕ.�vx�ί�ʮ���=�^���=E~���I�S����%��y����\��^�x1����Ύ���S&XЂ�hIT�<��fӸj��E�'�a⽕pr��T�%��Y���j��G2��#YZJ���搗��|�ހ�dհ<��=��I���9��;f�)�����2�)��
w�ƙ�d]�O(��,`����w��X{y?���?�ע�3T�0�.Kq��i<�2]S���5��1���Sp���!\��7&�.��oG�8�<�[KJ���5�����}�$�"h�r�F�_�Nk�/F�Wa��_�;��kt��Y��mՄs�#D�?�c4����nLeAݢG�#_�>�%���K����ap�|"R}�fubG�0�U������ІF���}�0�:O̰�Pռ�͒C�`dqrrًCU�݊Q�-�iѺ�o�_��a�mM-*$�UΛ5L@F
���^>�<��Uw�5T��);L{�G�X%�ˉF/�Y��]�V�[@��6A��h����D=y�5�Z��S���l�'ݾ�`�'"z�:�r���jK����.��5ܓ�S��k2�r�'j�oI�N�5��ڷ2�W��u�
�̹��Buc~�k�/?M K��DT]q��r!+����gY2wT�~�yݺ���
#p��G��J<�~�VlJ�&���I^9������t
W}ø"���}%C>Ț���Sz�Mմ:�qmgb7�����cfu�D�^��.�Q9rĲ�6�5������q>�u�D��$��;�e���aQZ������bg� @-��	�x�k��w´��2��y�eZ�� ̤=���:.�<�SɏA �GBT�������{l��6������?Z�'�����%*`���׮�/ \a�w�����v@���Z9�by-;�z���I�ɗV�H4G
C)����x���ڍ�c'QFZ���uݵ]�'7�);�`�_�'�+���A��kN����(��U������f�4���Ntu��HZou��-�Α�F�/���z_�>Jh����4�V�h�L�8�� ���h�Oɶ+W�B��苓/��6��i�?�w�MI��l��~P��ڥ�xe�����H"l(f��>UweAK�6
�2�X�����������P�8�7�j�FUSG�R�m��}�>�&���BL���|�����|�6:5�{!ռ�}6�K����C��K�H���V��^?&�Ѷ�W8o�Ѯ���6��\Z/���i���j+V{b��7�Ea	�p�0�ᴘQ�0�%Z�Vs�$��z��~���y�'��w��_|��	�1�&�^��8n�So�H6�jυB}�/8�r+a�#r��MY����*�O2������{>qM'�n�G�T�<�,U��+��h�1լ�Mr�7��^A�i�#zӒ#�RQ�[!�%�ތ���+�L��P3�#�Rސ�}9hYbUp��_a|u�I�ȤG���yF`�g���دN@���OJ$2�R�\8�4����T�z��-a�6&���r̙:���(�������J��
���Q �pƠ8L�&��#���>^Z����w��%�5��l���(���JB�͙#��p�����0�RB��9��q�o�gdY=�����g���$� �)({ju�E28VF{
� J�S�� ���sv�����x9/�b��z��HX�Y4�j�0�HY��>N���,���r�<,�2݄P����^����c��X�
�O N��'N-HYS���w�����a~�m9����s\���
��XlT�%W�Թd4Y �Aw�#/9wF��Ƹ`N3C�B� S�)����!CD�!��Ԅ�+Ν�u�:�WjPw�d[��z{�3�}t	�,�3�F�H�O�:�s��w��S�#�������+��x1�똢�F�*x':�Jg�`d\���u��/Yic��&	�)�,��6�A���g�Wa�Ug
K��Ý�(Թ�DvN����{؞A9P+��; �p��\#���ǎ>T��͍uX�x�0{BZI���~��u�Y�(���o�L��o�}C�+��56�`վ������5F�$jŜ�2!)�p�����[�Z�[͝m-���&+���P^�C���\Q��|�5�Ű�Ķ)U����ډ��6j��vS��%fǿ�8f� DՋX�7/*|1܎tISGHp�M-J87G�0�U�����!連���v���E9��w���A�L����5A��!�l��)�.���F~�,� "��wt.�͚r���[��ʡR�9%,��ɭ��L����|��ӥu.�`���2`M*����j�<U>ޖngƵ�mΧ�.�kB���?=_�ZM�����J�/r����)9c�@�f84J�%�2[��B7��CQM�][��s�g��R�m�VJ��S6��L|?F�V\������/{ւ��x^A}�5Z4�����?�e�{�$4��2z����ţ��& ����c�e kN
��_M}�O�p����M�jz3���UN����Ĉ���2�ƤRS�a�0�|]�$�^o�u|9��o�x��$� ��X%<<矆���!�TØ )�Yq�k|��ӌ