��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�]��Xȭ��p�oȡ�;u0ީ�^�)�>vys���2{�L�~|c_Iy�K����-��9!��\�Bi�D��{�Ԣ��r'T��NjH��ဣ]��9��|p���4d��oc���_LG����*k����۾�T>x�/>:��e�=�C5!)f���86�$����ԤE���oZ�&�x���� ]1����V'���Hci������I���-�;����{�gr�HR�l�q����~�n�2�����̴S�c�6�'o����f�?L�2���r�����uq/�Z��a['R�)9"+",��:�l/
����#���U\3�$π��`3��J�,�;K��=.�ʄ1���c��ą�&Y+[&��z{��/j��?|��~:�%��?�!M1�3?ߤ�	d���j"VlVg8��j&84)�|K�\�Y��m���TU-�^V <h�Τ�4XU�/6�����X�_A����W!��i��o��>��B��.��9C��iżׇ�2�%>+o��q�(t�
�%�\����·�*,U��y�oxmX S�`���;�F�S7�
�(���!�e�5�I��Ey·���e�`
&NTv��n�������Րae�m�d�9�<]����kw/��׼3`����ǧ=��ό����d%;�4�����"?E����R�m%���<�:F�Z�䕼jp�j7���P�U����AX�����:;��}1I>�[Z�洽��J�(T��(A���ik�sO����al�	�y�7�Ady�3� Ck�ѐ�9���#O�XM��@ŏ��X@���6�-i�� �*D�ӆZ-sa)K�7�
�3�`8�"\��u������Axw|*�>�y�Z��eDJ��rs�?���P�ι��Q \�f�Q)hQ�&��c�'��n.l�.'I�X	�D)!���s_��@U[%�Q�A���"��L��֢��۾����KJϽ�U ��T�/�f�MYA�����������=��D����e��|E��T��_%�����̸;�[�T�J������i���~��9׾$T�r�j?źR�o��*��C.�������uׇ<V�6�ĳ��Č�z<\�^?�����h�%X7�mp�Y^}Oa�V���_�L��������|fMX���M�T�B>�W�~l|z����o��E�m��9,�?&�����P1����_�"�A@j�6�~���H��7����^aJB��� �y��;l C[�~�c��6���솮ᶓ��S�|������nQ*�eW^5��m3�pP��$�&�A������MF�����:��l?��gݣ��-��͈�5���y8�+�虾w� �؋����M�y���hRr"a|�_�C���������+#<B�y�A�t���b��&�QX���ކ�2%�������6RY9JO!�1�^��nî���!�ܘ�ؠߥ��ՄJ!�e�}>4�/%�qS���P���u��-N��G9��X�c�y����e��	{�|�/�pj�����k�S���'ޫ�D�Hʍ8#b��H�z.��_;$���SК���<u�����"����_�V��U�UF�#η��֟�·9�h��Fڊ��>�֟*H/.�����͛l��A�f���ɔ�4���eh^E9�gĭt�Hݐ�d��7�Z?���4��)]���b�8o̮-}
����)���?Z �\/��l.z���]��ߔ���m1�	�N�e${�2��F��&�-;�����h9��H���) �S�0�+�ă�g����9�:FlpU���%C���6�% -�4�m�&����$�P�7hK�F�+$��E���	iy/��2�J���W�6�!ae�i\��y��d�����b�5{�^V�x��x|1XH��^��W��.H\���HP���t�������Q���6V4I ,�I�Zh$��?�͠�}�]�R��h��*Լhr�5S����O*3�R���_7��+n�s��F��G�U�k_>S�u��%����:ȼ	;��x�IM�70�c��?!U=٘`\Z�L#�$�e��f�Z_��1l����1�^�'�XI���㾵^;�>a'"�d�:���)�N�C���B��� �ȁ��I�N��޽d�d��X��n�Io�؊_� �V�?�wFv��jz��N�~�;#ŪAn��6%�z6ڈ��u�$P����o�؟��Tꇭ�zD���T��`��`"�����
�:� �\$ܕ@{�`���Vz�Ly��=�5%�ܳ}���r~\c=v�K[��s$
��3��]k�(1u$ȴ$EC�W��Z�(���)��w2!p�=P�|�)*������Ub5K�tSK2ȟ��Wp���Γ�]hrt�5��J<�5���C��kK����rGC�"�q��+4y�|��P�u���Y�(�Ր�Sg}�,�+�����a+��`�{�� {51Q�򓪻�q���V�Uy����,�S���0��	z��Gg�RZ�)�Y��1��ٴô	�M��9U]!��E�@C���Q'՛��v��6ͬÙ`�Q�.�@Κ)Q��f��)�H�ls�|Q=�r�0>�J��gy�`��M)R7rgBt񧻊D��9�%%d]e}P{��9�LՉ���eχ���W��Ҕ�:�p�تn����m���CYiw���sr�Q���]��W�� 4j����<�[w��2��BD'ÞE
��1��n���O�f�R����f�c�r�p�ґ&�� �B�����Ƒ�޳A�񌆘E캽����6G�T���	��9o}��Q��I\Ǭ:�8��H����%N�����=?��zܝH�C������5��C���L�m���m�Ǳ�tM�h�ѵ�ӮLXym[:�h|�7H��{�<�F�	�TN�R^�2�}���\�d��6߆�����l�g�2��#0�1���T0pK�S�vre^!���C�)=�o�� ��"�ZQ��&�K���7�����Qq�ּX��J�,@mG.���S�\U�I��	e����Q��q���v�"�08��9��OS��xF�p-��:K�k/{i#�2�����M-�{n����U���cL^#�U���~��w�7l�ؾR�1�k�ac�����t�u��C4`��(�����bx�=t y^}<E�|-���n�H}�K�E�m��Y7�/�$�(�>�f�E��@��zoS��Y�1�7ώ�N>����Z��5[���"!���W�{ļ�5�����~�\0	�d_h�����ſ��Y�#�[�zH��[��V5�� 
�t�]�#�4h�",��i���:ku��S�	i@��3UX�R��E�q;�U��2i�5ҝ/>@Y�� p]��P �'>���w�yRV�^E��q8r��h��;R/�S�h�A�/}�#C�
=c������[��/�=,����]�q��؜�ha�h,T�]��_@��KӐN�s`5�}̯-�����}���L�W����K-6�x ��J&��{��T�����r\`�����v�«�C@�.��EN����R;�����`���R�j^��\~�&���o�X��֌E�ň6�y��}��+�ݪ��`�8#�����<����)Y���� �߱Z��4}��ܾ���3%��{��mx��;#!��L���S�/Ug^�e¤���P0��ױ�vȶD�;���,�P�Pl���ż.�N}�!I�<$�%��,Y���\�Q�\d�<��Z�����(Q<T����_$�9�ψ�,�~a���m��Id�:%�}��C�>f��^����>�C)fAC-!7���щ6��6�oEK��:o�s��7IAP]�4۶���7����14��S�Ю��(n�,�v�lp)V�/>Enֶ"y��.K�7���N'��0�+�%�0D}�� u`��oT�]ih��5�B�9�~TG1�!ۀ��i�<�59y�Nz>�m�yYB�B⎢�W"��_��?rR������K`�n��h.'�\��t*}��;�H�+RkK>�N�P��`�����t�p��U�(��!Hm�@i��}��<7+�{>�k\���Ƴ)��vu�s�{!�#��::�x�=�����3]CI�h�׬�~�U����ez�I��J���n�b�ʒ��)����wȼ���П<��� ?���p��j|��f����+S� ����T�ed,:�z�3���cVR�45A񷁵�5��/yo�p#=�3[
^���M�7���� XM��+�($|�H1+mk��0w�c�,�����u@SC�V�o0e>��u'v&��}�v�$hlh	_뵯������h{����#��Ce �\"���V�^��aS8��%�%t}ө�~<n�%�?�R��bX\G�F�U4�cͶԑqG�yE��Q�lӰ� w>�ogp����&�U�{I_wK��t�)�Mnd4�-�C\��4ڢ���%���U]�4�<��Ѥ�ְv�$](�����)<"v�<ZC.�g���q&H׉�E ��W�C	�_Y%�_�v�ta����[B���~g�pܴ�WC�)�>�|��P�P*�����yw+��)k'#�R��tn��kR�
�P.�˗��|}ĉ{�?�K�W�)O��3�o��b�#�u7�QHT]�����w\/�խ́�=�d`[j^B@-���ޥ���~��a1�S7��ԍ�x�����P�����"S$
�j/���D���d[[�3E"Ԅ�L�2����X<�OX�讎�
g&,���^^�X&lZ>�Iֳx~���MN�o���Ó�����'��o94d�y��P�Aȇ �\�<'���>h^�X�нa"����mlB�N���I}�g�'a����\�M��tq��*�25G|�gE�Pӌ���qk��&�Iz����kV�D>S2�tF�����
�P�M>�(m�9�uN�G��94$6�J�ѵ%-gJp����M��;hT��� Y'���r�ʑ�{���t�6�?����C�����VP����L¯׍ϔ���
�~&QɵZ.�:M��/��o���L�y�<�R�j��B{�%�.1��T��h����K�����Gp�&��6��*�@/��Әkr����>�� #@=#v�
���܄�_;�1m�`pD�8��ep@���.���!��_�a�d�b�8.sY�[A�_R2ʤ�A�Ʒ���Mӱ2����GTTï����ՂA�K4�ptYm���d��a�V>xu
n��lD,Aw�2�C������p��< �koq��8v��u?�%p:#z9~K��:����C��KƲM�.��dD��/g����!����ͤ����|E���Yi���]��;����a=��1���mԑ��Z�z�ťP���+�2ڔn�]4��	��2��2֣'�.�$�S������:y�2+��n�|�߉-3�������WGz�����z�\+��@������RW�i���(�b7�R	l<X��-E�5�8� ��O��L4��Z�moy�~�֧O��^xO�Xf�*�B��,�tjV��L��d�I�O%�t}�%�6{��l^O9�*V�(c��0β�@d���l�X����Ʈ�8#W�O�J nw�Q�]Aa�������0js� �Z��m-,]�����'f��$��Ҕ<��{8b����W{���P܁(��=;^Uh�����]a�u�Ȋ
���)9�&�>Aa���ؚ��8�(���7s¡:�UyM��%d/@�g=Z�45�t�ޛz�H�j�6%'!���hA�1(:���_\�0��Ӌ�U��� ���6q��I��h�:���6���gQ���T�h�.��a(V	V��
���8�;�EP�m����Jة���S����w~.<Y�]�'�Qu�%Y�A,�qmSEU�t
E�6