��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jåا{�\�u�?߷�dn@6�zf��r������;�fyk>�i0C���<^���W�����4���m�8X�!0���8k�~~�� +�,-���x���Rc&�~�H��U�܉�i�5X$"�o2��%��t��넿���:ú���t&¸F�Uo���ও�b@�g��@IqU����D<�r[��9N�
�.eq��g�u6�xG��]�aP#�2g��W�� �Y)�H�5�s�`^ܤ��e�sB�Jؗ���*��s��H=B�B��J̼&�뺾K�q�+_as.��L	���[��;��@\���WU3!eU�+B��:�N�8��#�jS��������;�dF��G��['���ۅ!vU������B���Z�2)d��x��kR娥���V3�?rc�CF����5�՘]'�颁h;����ϝ^x��`tJ�	�M�v�8�+�D,D:I�B��*̑xv��I��i��|*A��lP
���Ez�p}��#��mj?��2=�hw�9���mӀ[������c5����<�7/b�$6ݍ��҂eU�q��%��ׁuǺ�AQn���%�-j��q<��(��
ܴk�X�� �k��T��s��(^��uz8�CB�>VW�m������Am�� Ao��3"��mE$*���˟L/�<���%�����{uծ�xK@�-����ƭ�Җ�3'�֯Rf�:�%T�
4۱��:ɣ��.�ۈPmA�3�7����]�/�^f�q2~�8y�Zd�ӊ�k��UI|���8 �~���z���ߊ�k�	�Fh�G
�ؐڨ�k1[�C���{ϰv�,#��̹�O3m�b�<~Hq�c||s:X����sWx�}�C�hN]�u�9gM�x���)+�Vr�y���_��y#�wlC5x��d��LK�F��y"��W�$��eOA9�E[�U$تHn�=˫q��E�)p���>�{S*�tp����Φ��𼈹,�E<�H�Λ|f�����[���xmZ>
�8c�x�����uB��5��p\ɴ<�B3gq!���>�ȕY}�7�^ñ�ֱ�����K}~���*eS��B�`�uҡcۊ��n�3���?F��URY���{��I�;�.��3���~���iN�3l�&^]1_MO`��L�˭�TT�aMձ��t�s�癆���l2�z��Ove3$.�*4V& ��8�
w�1n��������(`q���>����h�b~d�ݽ�x4��W���\7�9�Λ+��<�� s�C������JykoʶM��q���1ߋ�� �Xh@GS�ӄ���%D�)������<f��=��i&Mx^��xF"/�*~
�����@/Sp�� �Ź���.���SqBYW�p�}Z����֧��#0K���&��u�4=�s�*abVs+ͮ�vm��0j L�.k�bpU������Ks�o��F��������wg�v`p��[O�i��2Z�$�
Ss�g�agCK�b���}�}����H�ESc�P��*|���>�k(jyBT�ˏ_QI��κ�r�q�+)��g$�%�j��(=@��"rc���p��tIE���F�O�}W�U�"hGi�X�T��vB(��P�5�W�W��p7��	�
��6֢�נz�vYjt�7��.-���LQ/@��znZ�H�C���J�{MK�t�ގ���>җ��S�B�����H�����]��o��lY��?�Қ]�"���Ec��E[>^oH��Z�6���Z ��~����Z�c̃'j$�˞g��ۂ�:c�M3+��}��t�����^�L��}*���;b���ď+�Nh���jauWәЬ���G)�k	y��q�$��a4[ 9��� ��K���lAԳU�g6�N�K��>a�;��ѝO��4��i�F��C��������Fu���ףɭv�����a*$i��I���)J�:�)�:�x��xe�N;b(mz�}��̑͟�������4�?ȅ��n�͇>�k��ú/�'; ����P�����Y��d�H�����MҘ��}���s^�ٻM0PW	�j�P��G*���%fE{��8G�1��\���.lG �.�.�2sM�1g:­߯J�}5>���>���3�D���mq�H��V����a3�	�A?�H^���Kާ�K���%�]eKZ�f��5)�"�H��c`��hB���V<-GXi�����J2��v�c���<n���)���zs��_�[L��W��Z�#�׈��9�0�Vc,�|4�j+\�� �K.�h�+����"굡Í�S�w���w�hg��u�Ko�e,�)��Nyrj���D��t�A<VT�+��3�XF>��ɾg�g�9Ae���
Y�f�dx���nkY@k�ܳX0c�u�	�q��l�~$�D��D��Ɋ@��$��&���/:0}s���`�?���8g���3��e��Z���:�3��9<��;^<$�pDH?�:�����W��{L�SE��!�Ax��Kc@@���9��b�[�,�\T�Y`�&y��_aיߧ���_���%C=K�?��R@{E곟	Zu �.-���b�ݦ��gQX��nyB�0��'��EU�{Љi�)�z5t�E�ر2r�=RS%��.S����0�ɔHZe�vυ�q��*Ntr61 YM3���ϽM\�(�5��3`B���S�d�,@��d�T1�Ws^�7�S�6����wvw�Y�2>��x_�݊�ٌ.����XC�|�fQ�-�N��ki3nk{�� u�%K���/�lqy��?P(Nza6xM%�0t
�n(�8]�̭���� �21I	����.�{����Ҵ��"�ܛ�r�6U�Ts�HA!o�h\�L�>8��ݾ��t���G�Gy�D�'e�w&m)�A�-�QՊ��z&�6^�F! �膣�����	Jy�J��nc^�s��V���+AtUz�G?^Ƹ1�2χde$u�ȗN�F���.�]�ˤ � a=�=�L,ܡ�p�b����ڗ�4Uʺ~�����&�i�ÚC"�5���JvZ�ǯ�p�8O����{��8P�$dBI�{6G��r�>ަ��f�r��Z~��,<m�Y�pѓO�ȏȹ�����c������ϒf����(�po���(�pd����-��T��c.�����;�0�.P��j�c��\C���M��������ޜQ��k%V�&�����#Ml���������䩸�wp����%�W�	���bJH0�ƁHS��I��C�Wk��!y?�{�}C��[�'_��˨Ph�5�{��3ִ�`��!���Nw#�u�����}��Y�*+���[>���	�/�s@Hΰ��C* f��i��v�����~��o����q/w�w��I	+����� ^�Le��ClJ�����	k�e �zj���*]�*sa��^:�MXjy�}A�j�oR�Et��b�f!�Q�<Z�)�pe=�[ڃ�'x)8L�N/'����يhr[NM�?�}H»,�
-�A��Fu�������%�PPV�(�%܍�l}��O��FoԈ���+��{[
���Ģ&��R~���eD��_��k`a�9��/�n��K?;V� �����˕���MV�׼���E��Qe�(�9[�2Տ�����"l�U���l�W���[c;�:\%�7"7��W<~'D����Mp���;�� �/#X�8�ai�ɵr�����nQ��[�u�5ps�ʖ�;���v��g�St���t��WV�"��-����Yn�+m�%B���:�W�K��.}��я��^[HJ�K�"��S�h��g4�(t���_Wi�*~�S �J�/�q�A44�u {ݘэ����ˆ���Z�|��>=����+��<�\;�8��2�"����JA��4���Ձ����M�n�Bz��}��
E��Ȅ�W�x^3����B�\�ǘ��	}Y\^�˅���p��C�h����c���M��}tC�k�7jt���0{��N"�������B�EjC� ��B����	��gu���ůP�-醊^�φ�*��w���/ςD;I�H�ZH�E�b��ֲC���w�<�[p(E�4)���Ne�����nl��٤n�2]c��):I���.���鸎�	ɛ�7=�G&	E=��y�{���}�yB�����_�����%�f�d�р���ǔ#?��.�N_>#��c�ڮ�>���W��xcok��ۯ�|�;�}h8�d7l����j�P��ȉ{����
�I���c2�a;�pCc��8�Nɯ9����I�1p��.�S�X"�%7��'�br�W5�Գ=�4.ő�f�r潸��vA��,�E:HI5��� �6�y�eCv�
���##"e�Y��j.�H:&��tԊ�d��4�>a��7���ٻ��GR�i���J�xš���ډWFpg'cǩ_tC%�D�<������HO<| F�z��� [�*|��|d�><1&��v�������'_9�G�X�Ud��վ�N@\.�B�".�N�v����������{�OTw�%=�M<6��P���kr�7�n9T�?��l݋,Y�JrĂS�ϊ��� �T���.Y$o.0��K`&Vq?�
d[\�"C��ܶ���rTf��ن��:���ɶy:�K@�L֣�=����C,���C���x���jF��p���1 +����*|���S�w�Z��ka���HӋ�����b�/3п�¨V}��,�=8�7g��<�eLBs���O+��LSi2���V�?����}�>�� ���]��O��3�>�.f����ٜ�h���Z�4�5��>F2��7���d�����mF���*��La����s�����I[�H�?�[�qpQ".L:T�@��z����J\���eE�*xV��8�L8�R]7 �%�]	@c>�4��j>BbQ*�0�(�܇}����ؒ �'a�U�B�[����.g�kT��ҹN�7�^��V=��"#_���)O��
R9�7"����.�`������~7�ER��tl.?������(�	�=2nDM��E���FJ�~F���Qt���9C���K������$9�D5�~�-+��E)<���wJ��<�AY� eU�42����a��e!/xr[����$��!�WSa/�֔��r�B����]�2Z�k6䲳�$�k��S�=�ǒ`+/���6c��{v��0�?�ZHgvm�*EV�q"��c޺pks�0�&&�}f�e���
Z)�r�F�*rW4�՘�\�dDh�@܋n�@��᪽�P���3�B%!w�@�"�r��d/p����{�`oM�����Њ�_y��`*�M���v�@ϰ��ш��Wۙ.������dQ�ρr8[ �B���m�h������X�w���C�����QњMDd�A4�'���v>�f��Y~�C���j"��)�κ�u[�Km�n�J�����8�	�Y��J���L�� �� �Z�6Y�؋�c�I�Yj�|1i�a�����ZL�� g@@,�h�*�a�Ӓ��|�WȨ�{��Ց��/�Ѳ,ˡLW���XZ������y�K�ǆM4j��7/}��ۈ5q�:�G���N'"1{�o��]�4*�Қ�W�	�1�ݤ!��u����bĉ@oz�\o�}2�!�c���[Q�g�=����(Ug+��(Q�K�kө�s�R����հ�Ej��� ���'A��E��y�۞<kEy0Q}b�����&g"�{alN� \ݼ�uo|B�'�]Q4!	�^Vʎ��-a��'���!�@��GL{��h�3�c5p��x͒b�dNEp���{N�m��,�� ]��ԉ�(Bڤ���Åŷ� ��O0`=�6Q/΁�6pd�l�f�}�8�4��G	v.w s�w�%