��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�P�;�{��3�OT����n/\�@���V�F�	G�V��]� z�`t���y[q����a2�,a��rK�&ί�8������s�zW{=��s'^��p��)��d_�y�m�g+L,��l����f	�3v�nҷ�ˊ�a:�?a��D��խ�%��~)c�Ϲ�	����*�IQ�����,U�,M��st8��E�߽>�"�A�V>;2!ٵ��f���<{�x"=�Ce�<�&C}�=�����ݔ��0����Y��y����ΐ��ؙ��U�	ǣ���rQ����
�'v�@���DN�����2��廀�/���Ӫ�(��y}?'���h��9:ID������V4��*Aa����|��ʗ5�R�s��O��͉U�8oJ��h!茐��G�������`�#U�q�S����R,3ܥ�4X�ކ(n���A�a��'�c����<`���2���?�]���ʻ!�R��r�V���n����^)c���~S. �D����b-s�:�H��2�������`8\��$?w"���h}m�R�у���ڃQ���=�sQ��K����B#oB,�F��A�ժ����݁�i�1�ȥ�g-e�a&��0�gu�xh��p=��\������a���$'�(x��'�j��Ah��z�Xn��Gg�5�b�~�������A�hUݣ�\	�!��#�j�Six�ϖ�l�ơX4��崪J^E;
P�xՅ�����\i
f��4\m?�֛��L��4}��f��a#���#"�t�}�y<�#4K"�:�4-*J�Ui0A~�J�ճ�x��ؽv���^W����<A̝�)P�����ysĻ1ma�����3i�ѝG����������i�2������]N�+�D ����Zщ6��F�~���.L���_C�y���^|2�U3��:i/�>>�6�ni{bF�e���8na;a����c�v ZUӻ����^��#?>�Z�d!�� r�Nڳ3i��ꗓ��{^a�ˆ�/�~hi$�t��X���%op�|�`,�O��"`�^(]��oE�3�ъ�*��(�
Z���Z�6`�#a�:�����;�m�k��`�a������w]�K�s��IV�O�1�ޣ3��d����dåɩ/J��D��i��0����M�N�d�rZA6�"jY�>�oj�k��]4rS:-� $s��������͋9? ��k����e�����0f�[ӣr�XF+��w�}�7���Z%�Ov�]3.�S�c�d[(��A~�Q���$탅\5mb��C��v>�p*Tzv��+��9�48���D?+$�tY��6�.<.�fà������p���b�����V7�f:�' ��Ƿ�EP�����|��MK`��Xk+�Dm�P��Π�bk���=�ٞ��T�T�Y�S��o�fr7"hgn>G6&� ݪi?.���y��s��uO󃕊�?�W�bGN�l�@��n:�b����E+�R"=<H!&ɔ�+�]�q����i�j�ā�r� B�)�.��v��S�T��u��&u���t�Θ�w\���#�Ҷ�~�-)ݰ��JYc$\v|a���0�gN��m_��[#h�����, �C��b�cKC5�d��KT����?��A���?)�?�K�Ht7�s!"��L`X>:���oo+���7>f6���g�w�R���0���8Z35+�K �.t��,ZR�59�
���*�`���!��(��C�KAk�[�:Q.-�/�C���Ya� �Z���#�6�%����}9�{g)�Q���1��׏�q{9�	m�d�&t���?@Or��ֈ�Y�r�%"��K`ǆ*�f�s��*���2�Lߧk��~���0A���D���V���_r�n{�&'�t�o�� �wP���.�*��w��Xn���7V�1��MNY6&��]	�է�
p��f����8�]<^zb�V'u����XJ�67�h��%�g˱��;B�e
K$�Lq�l��7�	��q�S-֜un��t�z������x���/�	�&�A�t����������ԕ$O$��oEc��<("7�^$��<�ƭ���jP��1�4R�@�o݇�c���1x6�:��)��8�����Q�}[��w���)B��`�ݏ��D?�(��uSN�o����.��6eO�*���|��[O�'�Z���ǥqFN��Ӯ"��U?jTG�Q��B}��0�w����H�N��Mtѵ����?�ۚ�.���8.����Hj��c��sʟ�`mTiI8�&�"�SW�����1?df��l�G-�\#h6������7;]�M�Q���t���3��pm�� 
�.�~��C���D��BIfErYx�%���b�䕷��(�rU��Y��E��uA����t�S2EfC�l�b��c3���3�� ��H���zPlW���pk6F3#s�b�HV��ƙs/�FU�4!STD��`	-�iX'��Ǯ������)7��2,g�bk��w��g�҈��l���0i�ҙ	�z���_~��5L�t4�v��SX+c�|^'���S����wF����6�?�2�߮��M�@6�ZVLJ�- ���l�`DH�cْ���l�	o�J�Xe����X�%�c��R��H��7�Y���k}_�p�����k���yF�����^�H�FX���/�C���6"��!Î� ��>SG����<��%N����%�����7�t���5hN1^��L�%(��M65��CM���~���/�Y�T��_���NZ���v`�֯~gt���M'9�P!*KQ��h�; )yCv�$�Z�7=��	:���JV�kZ���By�%r(�֘/0Kv�maS#5	�y6W�$��g~����C}z�Ka����B�T�v�Zą����\z:��G`�������G�5��$�Č�x������ro��7���#�~�-E1��Gg��@��������o���cB$
�{�!�F�6���u\b>���i٦+��Q?:_{f��NC洹篗H��5I�g�P��T�o�)a�ї#��4����t�)��?�%��v#k�am��Q�����T7�W}}�B�{K}A�����J��`��rvv��sE���ۗb�E�>�"�6j��_�!��1y��mH��yA5�>{�ZDٞ��W��1x+��?��'��.���� �^껭eX͛.n���`��rF�Ϲ.vތlmAL��D=�nP{�)!`������yh+�l��bו�K�S�{����Gg��9�&�����e�!��@�Cor�:�br�/ c��ǲ�����Ѫ�Jk���&���1��7Ii3޹�/��]ޥHL�������Q>Qӱ{Ң����Ѕ�����ÙW�HV�7#�F?1�'���l��hCh{{9�[�H+k���3p.g�P�D��т��֑Teb���CPhZ��y�45���x�m�R�F�W����ًEz)�hfv���ux��^�`��<�nӻ2l�����ꂞs>>���Gf�F�Ecg��YT�*~�/]G��|z�IǪs�q���I\���0�Sɺ�5�Y��Y��`����_��WᲊZ�i�3Gw���P�h+��$�7�eR�8֯�,���?qt�&j�4P� M�Wɱ�'@�_r��T�w^*{?;ڤ���V��52qO�{PHҫ��$��-�"�k-���R�_�*��E�-�~> �6L��6�x�"��� �����v�8�p�*��I!�G^խ]�'I1�Ah����3O����J� �1�e7繁ۧ�^��y
|�`-�NIe�(
��A��5�W���C��L�>�ը�mи+�"q��,V]�+�ބ@����+�M����?9�@��/�K�k|�0YD/e�Ύ(���e�X˝e+�Sg�)L�B\�qsY�b~Z/�p�/l�����2:3��,E�㲫�Г|��N�m����p�	ĻФS���s�:.  �fSZ��3JbX`�J])M�T��zK�!dM�7460�O��*�z9��o��c����a��\M8C&���g�-�����:t$�����R`��`���IB��ʭ�b�S������]�()����>�#��vSz�PfiR���s7Y�@��)[L&���/A�3���Ȱ��ǜ
$��6�;3���쯽<j��t&�2����9����IS�&��C�]&"�R�xV�:(;N�V����k����@���� 	�w�L��4�,������9���:47�i�[p�S�/( -�$MCf&�xm#���d��Hy�[r�v]%= |J$eT���_�KJ�����S��:в�,(�&~w ��]ŷpI��S;=�!>�O�'@c _t�(���<���\W��6-�2��C�m<�����;{��y�6�����k�Sφ��Po���7Ҥ�ieq�V+��fr�:���6�{���vz�{K6U0wv§Mw[�y�����
�Pݺ�ضlƆ^b�K����
R����gB�*:��#��ׄF���C~KO��pxmt}]g�_�� �����d�C�m��>��;���q�0 �,�4��V<B�S�?�<Z9ږ���P��hf敄�e���@A�)#~OaN��1Գ-� R�JD�ӱ��b�<"�����B�~���A�"��9Z�ϑ��Ӧ���t��� ȇ�8O�/f��]���V��W�j� �%������|�7;���X<�C=s�}]���q}��l~K��X��O-��� �O�Sc[5)�T6��g}y��bH����  ��tC� ^��}���8j���U�u�����B������\������\Gr.D��D ��)�wsV�i�	�\M$Ðn���Hnjm8��i[���4)I6��t�g�h�&��-���M�w��\��kN/��+ť����@���
{i��Fz)�tvvxf/����$�����~m�˨=W`1��9���������_�?f=)`K�ND�S����|�����\)E���Z�6	�x-�ij��@9�{k{U'5�������ٯG)V��Z�ŧ ��~ߐ���O�(adz�ΰZ��"C�U�x��y��6{��e�VY�א	����i��bQو�����N���Kf����*`;�f��V�p����S|�V�F/Qh��vE�����#�IuM�y�k+(�J�醸y�HΉi�p:���������w����;gC�@D���Jս��B�a�Ɲ,8®���rEO��x�or�Vl	MP��T���ĸf��
I�n}��r��(��>v�t����Y�e��3lZ�g��e�jpvZo5=�<�&�Ov�<.V��+�M�U����)�;,(��0���������u�tr�������)+l�|Ƃ^�u.����zH���7�V��l�w��¶�~�Lr����B���D������!��R�9T��������p�P�Huc��x@���IZ�vab'��;h����8�t�)H��y��-����4n%t�#���(֑؝�r7�	U�w�*��a��xvπJ�yI�	We}k������G����Vt�nE"M���V����@��A�|{�B�������j74-�S*��E�%���↪M������ϘV��C�������ִ��<Ɨ��BG���&>���"ż��p���>c6o�V����-�d¿�Q��J�Ώu��EE6�c�==���+_xQ�y)����Cn� ;Ii����K���t�J1��M�R A�	��7��ȥ[������z�[���eo4�; �O�{0�5���y��C��j���
��J�v�@�B���ڊ��]���,!B��`/���m/s���ӑ@�,�֞��#����#��쑡��	�N7=�6Z�.,�/�6g��@F�	G��8T����et��^n[�#'�ÈG����K�6�Lp������N@���!�~����[���S�
w�������'%�qC[QK�c� ���^&X{_��g��r��DZ^\���}��cYa��K��#hiQ��/^��L��s�z���+p�A���9��l� ,�T-��`��5-2�s���c���k�A�ޭ�� ���)��{��m�!�y���ߠ��2X	���aҲ�R��h�3��9=>R�І��O�7�_�~�/1՟�!�������7�΀�Tb{�"�R�r�˃�q;�t���b�e��u��m=D\@�r<�yB>���0�����P;?�R \�zl(���^O���2���ؼP&����[��:]I�66�9���Z��9ra��RF/6�S��߬�,,k*~�Y�ڎ|���h�ٌ;>J�D?��7pO��	��ӎ��r{AY�?�_I�HZ�~W�:�f?��ElSG��$��/=����6�b��!�+��RZ/_w�p�QU9>reLd��3^��Z��BBt�rH����(�u^ ���N�ʢ���b��}�b��I`Sj����p���9Q��
"�8���Dn��bOE<�f��B���MV���9��hP��bFx#�K�c�n"��Q
���4*�"�����W���w_}ɣ����v���N���b�SqYgI�&�P����=���'�(%��m��Xi{��,w���T����Sf�{��ip�z��D����������
���s>�/�C����H�G{������H��g��\4��䳃�#�R��͗�}�����y56�Dg�Nwv~�����;�Ka�k7\Ԕ��ݚ×�p�U���VE3�e��)uO��~����P��1c<��Ѡ�n5#j�dб�P���#<��`u�>�0`jR��:+���V��� �C�����g7X�D�J�۷r�f/�^�q5&n[ྗ�' �~�lj~���+��@ƾ�|�߬�lh���fO��3���K�� 4����ʪ�5I`{O�T;����:�>^��M����O�jLr�]�
�#��*�ݚy�E9"fd� ����������C�v��j�f�2�/��@��ԗ�y(BĞ����_��-�;��o��v�*��xz�2�o��+Jowat|H�H���vYy~��@Ei���5�jF�4��bB�e��I�G>�8lF�dD���W!��I����Q6�ά�5*'~ca����c��5�B0��J�,��(�7%��ͪy�[r�=#�΀��`t����Ջ.��]��RvmK�1�??X1|J�7����mQΚs[呲��P�����Iǫp� �8�y��t��~	*����Mx�V3�c����k�>�F��-��&R�؆���v�>T��W��J��Q���%R���/��C��-��\�8�:�g6�vØ�T��v��w��z�U�R��o,\�A���d��ZZ<)�Y��{wZʢX	��L��J�𻢼y%:�:�fźg�|�T`p}���3���7gcQ����G\�Դݓ��E��s�>�('`�}��D�Z��p��ܷW�[��.����M+Eav2����)͊<�Pg>�=n�ė�� [�[�Z�RL�檿�}W,;���#��<�6�d�:i��}��h��w�XaEBt�?�ݠ���ů��#��:�}�:�9~�׽u���R�S��&�8�.�N�{�qlY��v���%���՟��T��o���)3�[�m6ԙ�+�g*�/��&I�ӕ�}�&-ò9�p����0{�/б�~���ѵ�WL�����J{�4��G��m��*��.�h��r�.��q��L�+|��k���#���q�3�(tq��:�l�x�2˽=�q�`�"���r���ӈ�����s�t�7��vJ��a&d-"�/�֢��µ������$��x[�GM��X}�����*�����hn����}�4)d��q��iq�ӍCX�
j�
8g����� ʕ�M+pL�	�͠�h��,S��g���9W��À8��5��&a@��[�&أ�US����m�����!1���������b�ܘ�����B�4�t�xе�䷮��WY�s���@�-%�.{�N�u$?Vҧ�|/1Y��H2� ��=��hP�`��������E�{^ws���ǜ��:��oe]ɤCl��q�< \�$)��3��(8Q���Y阵�%���?����t�!���A�
C�Z���X>���"�ڋ�ƕ+�> ����� �	+0r5�R	f$�}���2
b�KG}�o�Ha�~�Bɩz�!g->��|����/>~B���s)�q�/A��eq[����F���zfr��_8ٞ�a�&�m��.u��R6��GA�U���nGQ���J8L:�(Ӓ����r�R����-���ǉ��(�"m��}��{�����2%��mL�w�:�z���(��0��lI�;ŵ��[O���>��t�0{��[Qᠾp1Wcq��:�j�ɣ#b�PH6�Ʋ��᫒�
ZC4ZfhU���7���T;�>��qG�r���a��:���ܙg�t��,Wf�dE���S<�9�U,�/��,]���<�K9�BSƧO8(�E��o�vO�t�]����Pܕ(T���o��D�A�W�@&6m�G솎�"�:ğ��Ys��pؾ��By��^��2=-���:.2F�[_ͻ/@.9�6L��:���oD��nM@i�?F��k�~q�]���L���M��-I�X6�3�j�������_�y9o9��]�!m%�Ft,*J/�&=2������`W�|��b�o�Z?�~*7�b�3�I���#�ȣBXT_� �����ˋ*�]ǝD�����g��0$҃zp�[䐃��O�Բ��P~ �nZ���Ɍ��w�R�Y���Ä�@��p�q��P���!��|G�;\�cG\l��E�8�ζ�������d��HB����7�I^�u4�A���$�����]d%!
.��wƈ+.�T�g#r�@�T!������Δ�T�9��9��PG�0Tviqe���������K��޵����;��)�oL�
�C�����2F@���(����a8����`�\"�H���>��OE�)��-��Ǻ������6������^g��BL�^]�^\�F9�oE�1�+�I�qF.k~��N�m�����k^6� �'�
M�<��{qY닗�ԡ�q�����茳V��j���ПY c��Q�N[��x2劗S����Y�-�J�X1ہ64٬i��ɽ�����G��uׇe֙������� �su�ymd�ۖ�'0���)����x��s�=�D�Y%뀈��l��Z(��0�4@���a8V�����٨N��z�b/�#I�������S���%Pw:N
M7#�N�1w\�H���c]��I��&돓Ypf߮��ʋ�U(���6{}ޅ��-���e�&��)1Rs4��e>�J(f��`��õύ9�-��>lxݴ-{/p���e�{V�� 	j?FC,ߋ�p��#�߂�x.��lH���g̈́y$�}����b�~qE[X�-�Z�8��52Z����P%6 #����B��3�w}�2s���C��>V��-\P���w� )j���;�98�z���R��튴:h�_w� .���u��\ȑEGA���.�M��(��x�ߊ�s���Q��f�J߬L@��JwW��H�r�:*�G�Z��f|��f��,�,I�m�.��[nn~猑޲�]�Jz7���>w��C�w��ROY�[n�_+��~�R1��l��"= ��7��� LP�d�^����`�N~~�c���$��G�sjZ�*v���t�a^��i�3/OFC�3^�W��A�je�� D=���gg8y
b�΢�۲w���b2s�]��� ��ۛ^��I�y%��%�08T4��^��J���i�2�*��"z��0Tĸ���豟�!�����M*�\Cg#Gy5�!�T���P2��B抻���҉�Pz8�V�q"�˫c\��
p����J��B�Z�(�t�1q��:1�ʥ	�l���[���T�H��7����7T����:�����J{ƣK�J^ůy�SC�)���
6ل����Ü���@ع!������B��7��P��	��v���[�-�H�s`��>T����o�mS#W��LG^����	���|i��<��-�4��mQ3x1�^�TD�Nz�au��!�2aT�|�P��W%�!2��yGe�N������hEN!�]���A���*�%�:#�
�p�>*�����J��עNO���czE#2V�р�=���x�q^;��$���)������҂�T�{��?����r���h�Dmn1T����.��O�Zp�(w�s��/J7�/m�0�D0]�s��i'u�S浅_1o�#Q%�4�X�1[b�Xu��{�~u��Ic���i���	��������E}��ʹ��6�QI� �ֲ���ޡ�qfƔ��j�2`�p��d�}�[�Ȋߔ� =�4�^��'n)��x@��#@��ѭÙ�f��9���^�yk.D��s�<:Z��y���L�����&	��d�N�P��)ꆱ�WlA�Tʆ;�I��>P�,A	��>_T��bV���ZC#����:��l�A��S��PJT���P�aq���u�.�St�CH�^��s�d�bH�m��7�XWI$ݥ���F���+ �6&��{��(¨�d*��'=mǹ�?5K�W6�Ќ6���3^]���7�~��n Z�F§/9�s;��7'����BP���_"A��y�~���i�E���k��$!q7%HR��&�`���h8>̣[�N �>���\���� ������PYt�p�OȄ��pp��
�%00�.��"��͹8�x�~�R�y�ˑ�2�l�K|�%7�ob��*�>ח���0	�_n�ȑl0\����
�f��i_���Eu���^�Z�?ǰ��\C����nu��r-���t���Y�`��?�͑�S�?AC�ނ7^�Ipn�C��P����$�Cz
A����pb�m��D2���6���SmwB���.����gj����q3%���,��7�̑8�7l�?iiO./�le%������͍������YQ�n�e���;�>
lh�A _��U�ψw�<5�	?+����C����PhT9r�h���D���粥�������U����c��s<_�0�{
+A��5��]���b�"!h�%�"�;_.�%�Oʡ8�B�-ʹnd�U��A0��!�L�q3��,�=D[Nx�����4���l|��"nX:/Ш�H-,���$ׯ���}V���qn��Jk�]ҶFz�T6�j��헑`�������!�,Q��d�\`�a?�<�M�\OD�(�.�=k[N���Ɩ�b����z�`�.;��w��䣧�ղO��S鶐&���h�T'+������!�#�م�B��$�?�HvR+����F�w=�4]� ��+����� z�����c),AW�r�{�q�[�ٲ�Q�%�;Dᄬ,�^?�Q�����2v�\�g��odu[}��c��ʚ@R��g��%z}K,�v�W��S�zH�'][���Ԧd��I%���v�P��� @�v�B��^Ej���=-;*�@ȣ3J�B�_I:�ܸ�nKo�H�39��[=�z9
-�-��s�(H�e����A����%ʙU}DF��X*���L����A���@�ņ�yѬ�Ŕoj
8J�
�<���boK1�0zl�A	�-I�k�����_�fb�I3�t?�Xȫb��n�T�{!�8���=��Qd/��w|�3��q��� �AL�"q�s8��R.R�SC�#�w�'��Y�~P��3&���;��/T��#ߥ�+�)��%��~�*��f�<������pf��	3r8xۂAe�I,"���"���F��ߜ7-�|h��Q�\($e :\M�f��x�Q������%K���+��ȟ脤�>��C�	�����k�}�$s���a
�2R9c�x�qH\�u;�2���$�y�ڈ�"��@Y�))T?�����0/#�N��^D
�������w�6^�J��Bsp���62��T"�SR��j�$m֋O�o�;�Uɵ��d(_�k�Hܸ����U'��X��EVX���P�R�#=.�Z:9����lGX�|�<=��Erz�Dry��:W��u׎d�Gd\	,i�#�xo���83aL�[��Eh6\"}?Op:�I�HAB�z�c�q�T~H��ä��f�G�U��G��x=D�]�Ǻ�W<]j�+�,};څ��3T;ʺ��9�P%�<Y�j���o��7��|N9�����(O8'x�jn��:�f.������-��f�#˞r�p�Imǰ6G�8s��(vv���)�o���TE(�r���d���lxh�����b�;TXe���M6�A�G���Jp�B�O:j�[����7険l�ŵ�j��O-��A=!&�I4�M-�B��BT�T�L��T�����!f���3:��Z2`r�-.��e�����ߕ����K�Qʏ)��*z<�<-��=I���!�X�Z�j�c+���� �F��+�:���R*��*���#6�Թg4��4"�_Β��������fnZ�6p�-����N����j��<�ɤ�]�%%e�O�v�j��	�������\٫�A�`Y��l� ߻���*�;zz1��Cv�h���g2��>놗��*E(��"=�c^�q�5�����<<����R��n�T��בq!x�M�1n!{ٱB����@�A��M��Cvb�uA�Xt��1I��m�c�������|v?9C�7I1�ݓW\�Dl�C��s_�V.<������@K �~��Fw�S��H�MJO��2�+��<s?�zr��+P�v�'Զ�⃡��
�j�bjR(�ɏ�Z�f�A�Z}��U�)��)�cF�� YM��ax���eD��2j�bHQZ'�@҄g{1w�V��IP�T�N��p�4��T@��);485K������*es� ���b�B�S���G�}[�!�d����524RαI/9���N�d��/��S="L���1z�=��"��&%���3[�	�����%����@�m�XC}�R�6]���xّ�d���$cđ��i����o�ޠ�Cg�tq�-Q@.<�0�S�x&��S�8ƿ2+�Wx�jT�����p��(�����?�&��ߖ�����[�%�)�{��P���7��v�j����C�Z�H�m�Ѧ�W��9!e��f�m{:4�ݻ�"��_b��R��*C)�����*x6w����~ ��#C٢!5�/�"hltm/9�BT��L��X��6>�V�J��	�e1	\�����X|^_4a���?��Sy�2�U�����I'�S�`|�c���$:�o�Õ�<
�m������1��g�ε:��֣��Q�8��>xL.k�y&T�w�U���)����*��oR�뽰Z_�Y/�Y�A�;i-V)�Z�o����R��W\{�,��z㜝�8�q��cO����J��Ck���bt& i�iϥ��w�r���{^oD ���^���Ƚ)*̠��u?R�]����G|�8rXo��m���~ZV9'oFM�E�#�6�������0�*�2'���(:;W�{�
�0BY�*#;��J@;�5d�U�p���ah�V;v'����"��L����A�6�m��������l������	�³G�ƴ�h.ws�j�w�5�2á���������/���q9��n����ޒ���n��`Ʈtq?KP9��^<_���:r?�?�Ѳ>V�s�Mͽ�7�#*{M��J���W@�nw��&�ZF�!-�br!���; ��]v��_�h{��-znK�&> p���u�Bu*�i�C_p�}�e��l�/�'�K��҆i3������P0�����!_�j�*�@;�[q�S���#`��>����\�fo�ش�\4&�yT�q�Q��SJ��^mU�Cm�M�����e�ȗ�R��f��K��29��7���W�hUN:�#��B	�OH�%Dw�S��l�m��M,b�Q5���dfM������T���o,"�ݹuG�֋���0�Ţ	mF�yb���J���Jš�gE����I��0���q�2�X��!R`68�����\LRw��m�
I�P׳��wu���p�"�s�P2x��eN9�e��	ݗp�Hи�fy:���&w�V����ְ)���|�bd�����>�c �����C*D�u���ՁI³6`�.� ���"�1ꞏ)�էw!��b�ƴ,�rc`H��������mT�pJ�N_+���޹|�͵������h�P�j�9��r�"�����_�cb�<�����R �B���� �挒^zjTVʐ���j!��od�Zv ]cr_����ݺs@KUy4���&�����X��նS��cx��rV���vbDZ�e��y���+_�Y�2�mo������E6���Y�QP#�y�D�����¬8Lr������f_�I4�OZ�:H:1�	[�B��Ǔ�Cz�͝BE���H�a��6��ƙ���[ˑ�L� Q�*���fbݷ�6���|��V�Й��e��/��|�:8�įy�o"{M�=����)Rƫ�e��
�**=��bg�W��H�t���N6�ξ2��3)�J�*�rÓ�DG������[�D4��Tz�z��8"�Z���x�K2Vo��|+\Gp\^�[ҪjeD��;W�,0Ko�Z�mϓ�ʥ� [�k���H	�n|�l���T��������I�t�]���m;G�X47�)"��ٜ�1QJw
���� |�9:����{�D���:����נ�@�6{h~�X*�Ei��@@���P|Ց��g�9;��6�b�}�O?���n�4Zd���⢌%�(����{������1�t���j���ew��?�w��k��X$��Y�צۡ�T(J�����+1��8h+���-���AV�9���"ms��/�[�,�4�2�I<폌Ahf;!�K�c6�:\��y(LY���d���|���׌H(�R�-'7������9�R�M�մ����K�<b�;��K���uG+9�����ۂV g��}��ik�@n�F
yq}�O�����1�{2�����m$�P�9��+��:(�"�ʹb<���0���=q�PZ/;%�~"�r���驠�d���e�<�=��Fi�Oi��=8�{����w��d�;Zb�
F0�0�cb��wj}"Ī�H�`�r�	�p��� ��@�M�A������������Jl�O���g�cK�ن�7���%`�v8y1����]c�X��_����Kdl�ν��!��PB|��tp��.Z5-�qn�#��j1`��7��`�xh+.��ڢjb{y~�_ZÍğ��g���2�K^��C���gj@T�	��_Q�P�4Λ���hT�Z�Wj�Y�Tu��!�`�N
XP�앛3����3圤ki���ţ�jQ�!���lˮ�����ܪꔶ�sn��3^��/"������B��/���d���/g�J��e�4Q��h�qq��Ra����Xh"DS��z=�2I�oVR2/�F��.	,�G(>J��Z5�y:F�P����9�kR�#��W�/�J
�s[���eT8x�O��_�D*r���Zz{����r�}�,�z�\f����8�<k�l��&6Ҟ)F7�x8#0jA?E� �(����өTm�U�h��)�0�I�G��k3+ʳIs�\��y����Ɲ]����b�z��H?�wj�H����������}�t��xdM��e�)V����y�+V�ߺ��r�Pb�.[@���{�<��q1k���-���o�����	�0�_n�:�hw��>�����s��R
��sA�z�Q�����L.�J�y��n��r;��(���:]ϲ�!�j��W2��Uv�����.�A��N[��9�)��u�)z�'h1��o������s�/�eB"	�h����_pݰ�'�<��پ�P��q���2��
��3ݕ�ĆK�P��k-_4�CI�!H+'Vx�
j��V"࠷C��!c�_�=�,g���+��n���j��f�n(`����kL�	�#�X��ɫ�8r�f*V��g?�IC��kO5M��}rJ�i 6��O�p4Ø��[u/�)�����ތ�7G.V�6�d�@Vn�))!
o%ž�"���� #B#�Ie�
]�vZ�f=�A�bh�($
����6d���\�-[^.��Q�I]q���Ȃ�~L�Tg%��	��&w��&+09�u(L\`U�t�?��C�֤��k�;@��G���s	���V���mB5p^�Z�q��y3�5*_^�=����iek��T߲W'�{�w��A��8p��U8���G�n{)�Yp	1���O����x�_�6�٤��6�Q�&E-�h��ْ��(���x����O���K�:v�B��{�*j_�(�IZ����m� 4 ޤj�g�U{��'�v�w�.�@i/����4�m�������<��1�I�(6@ۆ�^d�]H��4����.j~<MVUD����{.�#�VlS�T}Iv�%:����քZN�m�!uY�����A;*�k�v��3��(�V?��'˥�����A�t��	��+(E�p
���yW��4�����i�c�y5��'wޝ5ռ�P^��t�Z��>zCa�)��{C�"�B����̑w{�M0"�[j��K��0h�$WV��S�Ŋ��,	�dO
E�s񼍐|�-
��N��~����SQIvuz�a+:�}gm�2 [W�X �8���f?�Z�O%K�����%9��~j�.a�K��yy�M��� �r!���n(T�s*�ezi{i�
y�ia�P����e���J_y>���Zy��A�������k�S.�xu3�j�ݷ���Zb8Ak�T�����)�r���<����Ϝ/?�2��]A�g vDh)r���W�4ҩJ�$@)�3 2���w�GKWֆTb�v.���!��!~2'�)~!�E��R/�`Z�PF���Cm֒���i�Q�N��������Su?=�G��H�d�q�2T��l�}.͡�Ӂ��VPFJ�9�V|���P	�P�5���d���k�&�ە:e���0B�Q�ۧ$�q㲵}��sB����/�kQ�c=m?S����a���j̓���)R�Щ����0�Ψ#\���������D8�o�[z�23�[�j����A�H�����gEa�$̃��� ֳ�K�I�4!��״�t��o��\�Ӕ��gA R�%�O۸fl5�;$�(�6�b��|w�P�xW� �$~=����}1g<7c���j����Ʀ�Hk��sw��8I'�w6��d5�����C�-j�.?����G�t�V�lV8}D��Q�z��<B_?�ŏ�n���@!5rn�Kn�l?�ਕS�|G�o����1��c��(�
�����5/��gs)M�v���,��pvfW5�-��M9�H�c���쯏���]�j-N��+�O��̲�������,��;�gT�+B�Z�c���[�7��NG7s��H��GEhIn���`�q�*�9ko�"\u�ZɚFNj�/��~" I���8Gԡ^��L� 'Zp�F)�ዀ
�?~U�	�����s,��p��F{�i+�骢���p
�;ϦA!�4c0|�;��G,����(�����h��vI+�g�o4kq��d(G�P/SPu�^��ή�<���QŐQ��[e%�ߙ����Ժ���u�x5��(f�&k��A��Px�π��&�=��
�Z��$@cv���#Bt )
j_��9�*#}���{�_1�.�d�Ē�y���g��T����~C���\�ؐ���>$l)� �U�;�.>"���9� 淈O}�%�ݱ�z��.�0�u}��?�
��7���C��(�tuD��tM��n� ̽���ǵi�L�������}��^J�6M�G/U/��[�]T���NQ3zLX�R<�6�>�3�Ͱ����ѩ�1��s���0�����O��P/�=��V[s�5�&�m��J�v�7��p�{��T�'�s%����:m5G\�4�7�K���(�g�Κ�Q�T�k鈤��>r�ܚt��6��ҳ4���6�5��ʰ�Q9β���DM�eDv�E9.�B���.SSP�V()�� ź�5)9�nA��\a<3+�\{�b"B�*[|_��l�$R����pM�F��w�)zSpǒ��ϸcȎs��S�4���dN��j$��)��v<D ��w|�ZN���^��x'�#l��Q��}r��n�C���0���ootI���˸���,\�����;0OF*8�������:�*�1��ee���Gmcb!��6�T�H�4� H�,R����'뒘,���>ׄŞlc����H�e[�keJq�{�߽��?��E��̛�k8����g���T�4��!���=cbV;�L�Qࢩm1�P鐯7?��AOKV�ph�7��#�]���9�0����j�E[�J�ب���$Ÿ|w�
�b����ò�/l;�ʞ�w��"��qNnX6ݝ��V�^���l�}qt�'\mʙ�{�;J� �	F��H�ߤ��D��Fi�E����v��/[�H�hWi���~xk�sq�)�~h��+�:·ˇs�?���koE��h�q�k+Z$�@@~�������\�����
�}�!O��^����V<�Y��k��<{��&Y��s�_n/�
3����o���YQ�x������YA�h���Lc��i+��,�BYJ3���{�$����C��K�~Q�~����K]�(G%�56@i�5}�P&�f��ق�ӟUo >��%���#�q����ٱP�;=�-ł�����&d$��=�0��oG$5��giJ0�a���6k3�V��-iJ$��A��+*����:�j���PN�8A9� �+f83�/E�S��:��K���}�]�5�e���R���	��]*6�V��G4��c�<k����hL�)"qp''A�����#&����*>-�҇��Xj
-�Ϯr�8��_��f1������+my�Z��C�иѷ��2F�����|������e�n��/7�/����w'��LN�蛴�ۣ^u[V�=^Q(%qc�y���m�� o*`p���#ʛ��� 5�y\4�p�P��{N� ���+k)x��ʫ��;~��v��|���8�ׇ����o"~2N��]��Կ�ɯS�p~y �-�n�G'`�,:O�Mᓨ��� �K~ͽ<�L+��-f;޺��Ǔjױ��s[C��@/����U��PFP/Gľ��(��#Te�>ᡉ��l�:�T7s;�Y��E��K���F�\��BP�$��d^���.>c^g��ѽ�E՛HTDo���L��ͧ�\&�Һ=�}�oL�e�2�%�|��b����i:>��(~s9B�W�g�6����8�u:��T�E�]�B4�V��,lyKȻ�%:�H'Pl��m�����(����S��Pԑ�{�`5�1��걈	ѽ�T�Fr]/C�ɗh�ǟ��LEX.-2�p7�/�BbE?&����	�� ����
�׆�ޓ��}S�0e8s`�|��]���W�0�yO7���Ӌ/�8����+7��NH�3��B�S��*�aX�{Gt�jا�