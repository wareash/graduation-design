��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jåا{�\�u�?߷�dn@6�zf��r������;�Ƒ>J�f<@+ڃ��i��H�M�L���\�
z���o���uļN2UXG�G����p��L{h�x�5n�%P��{��0���M����O�"\@��g�=��r ���E-�Ӑ�RB���a*�WBlt�^���B��7M�@(P�N}o�cb]��X��t�44�\�Х���b�U;=o�Z�;K�w����t�t�-e�tPU0��9�(�S�|H�"@+��WV"&�A湽F%�.�#��Z�MQ����O�����.��H1p�ak��̢q��k]��6_�����b[o*2�|h돓u
V��E��uM����^�0n0���k�V��@`~���еb��/Gk�d�mH�)Dg��iTͬ���~kO��}ͩ�P�/r)�U�:p�D�#�@��PG�YuU��(��c�xb�v��Kn�KǤ�M��t��T+<�c.�c�f�:�H�=��G�e����s�22��8E�&q�:_���}�L/�/[䄿k�(�m;ܹM�����夭���F�nc��)����z�w,����|y��U�y��eU�hy�cM��_�=��[J�i�׆Y:�k�g�g6�p"��Su���Y�ϗ�bH�w�PM�
���4קɀ�XA%u@ �B���Lճ�<֠�(� ��>bGz1A� �v�F�+��Q��f�0�U���$WŁs�{�TҮHA�pF���Z���C��[�L/؟R�W��� �Ĭ�+}�VQ�R��.�G�����S[EF�xE}�oAT"R\k��Hh��iH�u�cq���������z+@�'��7�O@$[����/��1*��T}�}��6M�P��s���֭E�W��DE�e"K�h~�Ew�������=a�8ї}�5x�&:���kR@�Y[��t|:_;�~��`����+���F��<�=����<D�:m��=�`�[wُ����ƿ�C2�lch��!k��*�Sk�(��|S���S���LH���W��֊NEV�d�y�z6lq�2TtI ���`��v3�~���N��P�o/Vz�K�9����s�����	d,]NN���#mM��jp�b�;�f��@Cb4c�pA+��j�e/c7m1�s:W�8���Z!����a����Ǜ#D���қ	�4�^�Mt!9=��Y��s�͆#�f�y�"p���tĶ8#���%.��C��k �W��2߀��8���a�FZ�� άx[e�����!�{J�K ڝjن���LTQE�L�gPP�EKMb<�w1�c��q��j��^�����靛�N��B�U,	�+���t�������J�_��s=��W#JrXh�>נ��� �}���W�\�B�2�-R����5�6q�|W��#@\:����h�)�l�lq�E�����h�͂+�����#���w�K�ʨ-h�I⽥2�O33ct��6b�MSg�c�@Xϸ��`�ފ�Z����p;�p��8����*2+�ъb�Oo`拥*ݺ��0�O� �2��+D���-�����4�:昿�gbQ}Wo21��c�	�cp�J"jl���}2���r���$����e`�r�sr� <��dp�?Xy�8-��%^�Yڴ1��%�4�d&��%�N�e�.n!�0=y2/�>��ئr?{:4&]!Y��oН��rL�Y|^� X�עQ��Na�ʭ;�͍Hv/�����{6�50&@k�l��9LBR�����):=� Z����Y3��Q.e�jg�����nź5}k�; �9�7I,����a�ˣG�X��82��� ��
�b��V�>-���>b���G	蔴b�Tq-}�oג�.���.� 6�4\�a?�A������"�a��)f��!�l�V�X|/�\�qH4r"J	NKNWu�o�	:QK(%��=v7�B��b�j&���{̚��C�TΠ����}��20����C��=��n\
�o��C��Q�=�pĄ8,�����&�u����8$_�:�ca���)�R5G����ܟ�L�8�Z@qk`xʰ���ߗ�3 ��c�1����@��֋R6Ȏx}?^$6���8|���V�*l�A���X��%[����u�7ʩ�L>�]B��@B���;�̊�����E�Ql�u�\���9z����{,�(���e�r��rD��ם4;�!��Rf�X�a+���+Y}'**p �m��Q�A�t��TJ���H/��23t��)�|��T�o�y% ¶n�a_� ����(=6�*�MgH�eԂ�Ie՟�?��К+���w�{�u�FĖ.k���aZ	f��>�ڰS�ڤ+L�M'1j�Mz�?G��x5��Dg�1��ˣt�kQ3�]g[ٳ���٤��ƧR�=L��6|Yx�1��}�؈,�l\=�
	O~?,8�F=]>r��G�Հ�}A*�"�i��G�]����S�FbU���O���2G	/Hk�0ޢ�x�\{b�U�Y�r�G��6��/#m���юG;zL�m�
gUR��쨗�Ò�O�^�I�����	����1RIa	�*�������]0ƾ�ލg�u�a$T�k/(���_�Y�����t�=+�z�8;������!9p���s}����-�́Ő�����;N�g��µ��k2�W�۪~&���:��`�c�η���lF�F���+$���ОNi��GtH۪��X�y5F���B�!_�?:��%��ÿ ��Sz��z	�"_�$�s� �b2P�h'w��KrȤ�L��%�H�Ν(�N���G�[�<�JQ��@?�]O%�����]֧�lİ��#k���ZV��{A���e�Oғz�;}�/�.��wY�BD4x@g��W�������֑��s��Xc>�v�vI���s�|�zޟ��>���}n{�%��i��M�J�~b�+��ow�.$��]?�źbmv���t��%�>�i�㣫H�}��?��N�d?8L����w��Y)wC~�*T��I-n`�^.n9��,�6��mw����m#�t���Ba��D�Pt�����I��J�mk��b��,�N�H����҃o�$6���,�e@Io���f�,[�&��v�	���uWm�>���&'"�L"ױv�Ew��� �xJsg�~�`{��R9�1�b����z�p�-l<N���b�SH[�x���'���u���v�\�fW=�O��&�~��$-Eր0Dq��D��#A��*?+!l���b��s"�櫬���q���.ռKԪ�U����	Z"�K1^fbZ����.w�L�$�'�|ۼ��,��J��N��
�8��'ŧ �`�n���̵���9B��p��GH��eI;H��EMQ�X����n�~g�E�m�v��[//�Y��5�vT���u��Bgۼ)�?��ȗ��l� ���Ap��f�H�l%e]�Y��;��<h��E颧���V��V�ȟ��U���Qa�iʤBX������x,���8Uer��Z=(�}Nb��2�A�`�M=2�,O}�����FiA�p�Ud���#�=N��9a91,�}_����pCI��A�A���`5\�,��j՟��5���9%*�_�y���,"��:c2N��3�ת����� ������(6<�c����G/,s�'N��� �C���Me��췵��ElS8զ��@��K�(������T�/���ī�V��<�&��=�,�8b�,UfTf>��i7Q�0j=�
�I����
���6Gr�x#�f��˝K��N�q��ί�� �\���G�[yV��i�<9Ny��j�f�c�ZT�K!Z�[H�T駛�7��7�<|�����z�3��7n���$��H_$ߋ_wᴥ�`jY`��|h�ꂴRU����1�V����!�d����,e.�5!�W�(Xk���3I���zX�U*`��������ue�o���`�Y�����4�J��;ic!�x,l���1�w�hH��a�k�ή�����X��_��w�l/f����;d� �j	q�>@�Y�����BKиt'��b`��]Rs��\-o̠�����+O�>+�"���/���MI�<�o�o7g��8o&<-"'��N�\k�ryy���� ;�d��^;6T�\ed=s}�V�zR�X������]���x�G�vL������x���g�Qg���~�,�jc�"�H�*�\�F���\�;����59����T��`3Y�g�q�8����oWn>L��W�)(W�@�h*���@�Ý�/d�F���/�W�1hՌ?y�%H���qz����M�/�8/ǝ�@�=rO,�i ��3�?�ϋ��Ы����0cׯ_]9:Լ _�}(S�~�b��F)���R��dm�w�(s5��[#�!^м���K�����<������%����2�%�*u.��%&k�cQKNߠ:~Oҏ���`��thg��\�D�i�r%�V��!��=�������Q�̿#�1�C�F��T��c@]�O�uTm\JJV���[&G��i�����j��$���?yS+�1����D�sZV�e5�n/�I���L��j'�E�^���ƯgN���}Д�旽*�<���b�iH}��zӌ)�9G ;����E�y~���Z" ���8*�Qxf*sX,Occ�֓�v�������E�V�%T���Ov{(�Z�Qd�j	�=���Sk���v�^v��0�����5,�הFM����i���5�͕>i�֖�P���oכ�d�~D��1?���*��_�S��ɓ?\Xx)��T0� ������	�2��h�חي��}��d�·�W׭k"��*������u�uR6��_����O���\GD)}M"}��J	0tt�{��gX��&ȳ��Bw����XkE�^H�Y$��R?�s7�I܂����q+A�� ��?�s�@1{dq�^J�L2����*�ӡ�����f�0�h�Y:���]�cZ�)��$z|���6�+����	�k��F��̹8�d1gHY.�}XC��N� 5s�J�<E�j�֑�|F�����x�G��7�Z/�y<�,z��m5�S�ڠ�Ϋund�qٝ��j ������7���ja�o�����d���v��k`n����x��O��jVs>�X ~~D�9#E���l^IƊ�SE��~a�Q�S�9)����ϗ_�6�����Hw���]g�&�]�����,Y�-
yN� 1���%5�l[�?j��S�]�������]|JC��o���G�q����I� tP�~�[��i�o0��ŴMxui��,��.g?� Sg�1h�DAv#�%qXB�*ʛ6�x��c?�B�E�zZ�2��S)<E �l��p���E�Qva
���x�W�����s�a���aE~�M��8�O����=�Ą�?`;�v�ws�ڵ]���(�hE��s4)��8�N�F�"�tLE�`���#��������)?O���j����cN
��JW��*'�dͤ���@T�M�Oϥ��+��@##��^�/�dGV4~/=��@���m�!��2��0�,�Y�$hev�V�wOPlޅHU�>�~Xօ�l��\�0��)�`��yo>`gQ���C�E��Z�8�7f�V#�ɔTg�R��V�awF�KY�M��Ut�<߇DFf���/h7�W���G���|��[��Bz�2�ۈ֘��N�A#��V���A�dn)S�.Z6fDwӄ$臾�ތ^gڨ�Y�o��r{ �W�&�@�f��j ��2��X��o�s��r>���#;��"ڡ��Bm�ǔ���֔���?�J�iD�f�����磠BQT�n5��d��'w���;=�	6̶�#��.)����)�\��aq�7�SG�<� L�#x���W4a1ڱ�7b�eYϽE�E���i� <��Ch���=�hS�a$
x��K�*�_ߢ]Ud"� ��d�t�O
Sb���x�
�l���n�s�z!
眀}�R�qO�A(f�����R���?�j[(s�y�ea�����E����l�%�Vb����i����n��`��`��ݱ;������b������M8BK;q�b&e�j&��@Ē��3�Mv���{W�>At|z�9��L0���^��<WFvf~��G�d�_e�T�zlh_����U��sؾ(�Q�;���{}�@{d�jr��U����$iiqd��.~�
!k��S��*�mS��[d��!� /��N1�yDɧ�� p�${;��곮�fܔ�_���`��Ic8Pb?	�ܫ{e��,�8�!�LK!��j�8_�[�B���3�{�h�K�
�����������嫰%1�g=�+zxK����<M� �
v��w}���έگ��9%RwU�2�h&���m�r��� >� ��>�]I��`�Z_[��r7�"��mT��W�TA,���#G�v^��%M�׹��bN���C�c$�#Lq%/#���j�*$����I�R���D�I�v����U��S���J[�X��3	��QRm���r�F-��'��	��� 귈�r|D�اNqC�ܔG�Ȉ8��M�e@�HC�XL���,G�����c���$�t!�*���Փm/���lGV���Z*�)AE}u�
/�I>��7VˢP���L�{���G���7�NA�������<�T�㌿2���?	(� r��۷�2s!��פ�ŏۡ��4&�4�\�DDF�(���۩p5�&�W���A��h��0�X/���V��(����6��s��ދW�z!��6�9$W���}
�ʑ�Ysu���LC�
�:�.��g�E�Z�����< �"x�i�����9v��S�ҩ�Ͳ�O�?]��-%(�y���d�6�ߥ����5��4)D� �ɌJ����8�!�����9?��çy�ǫ3�jg�|��N�S�vNQ�ۜ��/��%&8��#���p�f��p1�Oa��l�aٮjt��;?��q��F�Viq�A�&�z�k.�/�P�0<z����ָH����h�v��ݱ�Н/�ֽ�ЍjW�u1�?�Z�Qa�d��Z�4���qJ���8!�!%m���;�z�|t��tR��vE����W��T'��tzq�s���1�D�Ϩ�@PMٷ�WF'B��(rUd&�d�!��k���=���.!;K���z�J�u��cT���D���L3����t�*j
5�C�F��?$���۰�-C�S�}I��f4��{�e��F���,3�m������\�����y�q$�8�t�y��wlY�+��h3�su���O;�B�����b��� Ms
��u&�=QM�)�kkֽDO^�W����}�+������Y�&,�Dn�jb���*��:3��A'����I��A�(o�V �^{k�#�Gf�4��Ѫ�*�L_q!< "> ��>JӲ��9�=�J˥-���#��[ ��_-�զy�e@"Ƽ��yϩ�3�e����, ���XJ��C�2>�#(�w���W����j��di��y+�]�G�g�VQ�|�^����tޮ����`�S���$�a&��[ J{I.���{��(�ȇM}����G�D��9,+L�S<�/M�
6is��LE�{,fU���W�ZϪ��fw(�R�R��L��f�(�z� $��zl͎��[$�Qc�5�U��:��N�h��X�3����3�a�Y����c-�6'����3�?�B�p���qLx�wոUSCOL���IyY^U�U$�>ܿ�q�Iڂ����Q���@��5��8�L��޷M4� ����h�kN�!���7U|$|���mG��O1R��gS��B@����b��\Axڃ��<PL7��,��f�[0��yض�|��Z~ϣ�ä�L��)�#x{���
g��.��Z��K�H8[���k��ҪM�����䳮*�ȓgs�zD��.�޾a�;S�d�1#�Rſ��]��Ac^<�ބq�Ϸ.���*K}H��P���-�|i!�,�8�y�Wm�/>�w���l~Н�nP�΄k-ʥ��K\�[��8���>�ߊ�
Uf�hA�t.�Q��plL%�c�jY^��:֭'U���S����?��u?�F���k��OQ��CCQ92%�c�_2vf6Nl�'�	�1���Kߖ�}�-*��ّ�I��.�&�{,�9Y�<��D]�~M�ؿI��k��zҩ�'�*�A�7��.N�M�E)Y�{�܅h���M��L��'�1��[�+7�����CU�Ɯ
;wǭ�t'���!�k��艦�y-ч��LV1�����v��b��yIU�ǂ=7FZKo���������`PIz�-g����B�u��E@C�G�gj�/	�+��0�U>V��0?wD��9cf�;V1�*�;J�Tlq�v���e��i�Ig�R����Oޝ��0�y՘@�Ĺ��Q��Y�����#0{�����j�&x�����Wc7Y?=��4kq�bp�����Ϊ�Ð.L�2L~1[Fh3�����S����������1��#��6^+4�J�x�=�/5�cs-����Ұ�=+�H�֑���㹦U&å.	ڇF8�)�C��k6`7�Z�P.�����x�[u!,�E<@�ba��t.�s�<LQk�1`3�C�����z��1�5�ES~]f����������ah���ӹW���C7�d���G��<�ͱZ�v�M�ˑ�"W/�+�
g g����TڏO����jͳ�h=P��S8A�O�-ȷ����0���jK�<�٣Z���փF���\�R�vƱ�oX�c%pN*�p�p�-�F��@�Uf/�<�A7���]Hs.�i���4z����;*�Z�t���#��7��_�=}�$�5c {�>��.���+�v]�@�G#
J�(�v0���YX��y�Z�V�����1)v�������7��F@��h�v#[��d�*�JU��NJ�z �
ǵ9P輣H�����l���0%6f�!dy9U"���$[�!=Z&���qڵ^�֪�H\ N~�5�5ߠM0:.�sk���Τ��Z(��5�g��4$o����]��XcJ+�
f��\W��[SY>Ͼ�z���  ٞl�f����h�ώ���6��8�2��Jي��Y�|SS��6�.��3��vϸ5�jq�V���M�]T�RaHl�>p���������!h#^P�Z��*N��1v�z��D}���9(D�P�E��j��l�& ���wz�o�[v��*�؎~o/�UE.pI-�� �%��y-8��X!��؅:���߹��0��9;[wH�^*�_|�o�⒎�aqU/�e-�&�$%U%�ž�c���5���R~�ۧASh��"I~u���셶���� '��s�6gv�eA��^���CS�@��>c.�7�z��Y5Oa�!�Sw�6/|�f_�
���FQ2�}Q.���(��T~�{V�߶ŀ-h]n��������KGm��vQ�Ȭ}��F����_T��e
"��/�6���	��}�E�!D|�5�̉{ہ�J��
���1�	&�g~B^�O�蟈y`���yT U�6���H^��.�c3A�fJ���4=��ޗ�Z#O`��S�m� Ls�5��*Z1I�+��G�0R�L*7�l�U�,�����`z�1)i��T?�b�o"��P��_md� �Gj�����;��2���)f��Y��Ż[��Aɞ�lѥ/���f��<�+|v�TX�v]�e�]���B����զ�j�s��š�]3��CL-�	�@mkvӺ��m+��U��GUcF+:Y�z�g��|t�ʯrRI4��:uo���:�$�}(�B�u�5сt�~Mׁ��*��g>�k����8�e5]�	���.p
Q翘��I��嵋����j'6-# p-KBK5���J�3b��Z$�������5/�I��i�'GY��6�<&2��ݕ�%��^ԁНh�<6�2�H� EChɱ�ˀ<i��+�T��UC�(d,*��sTeƏ����qroC?q����9mB���ʄ��2SyB���I��
� X�SI���xK6E,`�5
�%�8���k�����_�c�^:[a+c0�ދ�`͓��U��������g�������P�	�_m�-.��M^5�`5p�l$;�Ԇz�9r���c�Osi�#$�I�1D/4�h�3��|�lR_�AtS�0s�L㒲O�_}���b�T�o��O�4����M�̕/"�d�d�>8�f�R�O+���y��=�Y�7�dm�խ��=rT)q��z�پ���y�$���ѿ������A�Ƶ:��;7S݃��s#���_v߄�x2ý#I	�����P�gz���gpl�n��^]@�f	�aFwn�2�vY�mPtT]�u�j��	�.�$�j=ǫ��r �-�M2��ʆE�ܺ�X�1������ c�h�W^R^�*��r�k�^߆���E2$Ufaw�*7��9�Z��}eI����z��ڛ��)vKxS��md��,��+�*�>~�G��om$�O��j��- ہ�ЏƜ��e�1�f�tH?�̀���k[���auo׳�m`�3d4��7�Wn饪?��ާ�'+�+�#[OT��^f���qĬ�M�	��ȷ)�T�Hh��Ůz:I�$����A'���3���4�:f�?S�u"\ё�Q'�'d+J��1Y����U��'RQ���ۢ����,lG��[�#�m�v�A��{�J5.E�=�L�J�ne�^��}���eA�ӑ+9���,9��AMѤ�ܟB�3q�ʄ�MҢl�����ؿ�rVCwMC �S4C6J�Q	��jؚr9f�*ޓ"L(E#�Ǩt`f
?5r�(�5��e�]6M히�I�2�vN����6���y��(:�<��5hJ��7Q�Y	���!��~��⚑5�`ʷ���'8�Mo(�E-L.��%M��"X� X�}%%�y�;�A�f	~�.�B��&j\�``��s'N�������$z�Gw��m����&o_u������M��D��1(vjU�V������ �lBmR�	��η�<�5���]×I���n�'�m�O-��T�V-+���Ӈ?���3���f�[g����e�����S�|L8�z�Ǔ�ʠp.�j�#���>>0�4y~��y��ɻJ:۬�1��JOoq�.WS.���ffn�xE�ُ���ֲݑ�{k��A~L_�٩<*�y�# F,�=49`gh]j��%:����P�@{��ڵ$^"!g�d񡩣���_���L$&�:��v_!V�}�ް!�S>}�''�����x4`	���AO��.CZ���H��:�-�"�9G�b`�A����l�f���M�+�A�P����u�v�L���I�iM�;�O�B޵����5��h�����x�.�(��%���DxKtl���}����Α ��g�/�Y�?:������s-�/$eq��X��ϩ
�L�̠�W)��j��]z��*g�m5>��Z�	��!*u��(�R����^�iwo���h�����1I�Ԉp���xI⋸^��t���7�4�L�Dn�_�a���+�B������C:h�+��7�U��_�T�>=��E�7zծ|�=�w��꼥{!j��s$�>�0z[X&mDƹ�X�kzD��n^<����)���TH��&����l�5�TN�{��
���ٞR�q�[��M�zt��s2o�a� ���m
{��Fg�+�LfNb�xr�a����&eY�Qe�p7,q��6 ��$�#�u�Vkڔ�z+$�����yj{��u�r�f4��"�&7��U���Q߭l~�=`��|���c�)
rA�1��0�ƻ_��^���F���l,>凄:]E�baL+3�R�oTi� vۻJEz�-&�Պ�QC�u�4X$��`E����9�����yW���{�<��յE�����*��<����il1eM?����,;C�^9�D�>��cfx�T�^h�شf�R���9�M�P���~-`���;�㧛�J�0o|�3X�I1I�p��`�~qD�m���2b�CW~~Y�I��1����2����:� CV�e��n4�`����㩑�g���Xw����GpvS�f�JԄ�'���a������%��r'ꀸ�+a��O1T�q8
�/Q�|�qTR�]���e��ZR��C���W	GV.>��}@yv �����6���'I6m���Y����b�$����<0�K@I�)]�Q�'F~l P�.J��$D�`��Tacv���dKM9� ����n��=�	�M?���z��Uƨd�\�܌���ќ�{CZ��'6��l+b=&;Vڑ(���\C 6�e�9�p��7cTw����\�	@��'Qk-`��2{�Bm5��+jV����%23�C:$c��,�������' �#"F\'���gτn�|���I�5%fq�4k�x�	d��F���ǥ_Ѳ	�0&�sg�E0�6fֈz�+Sφ������U�6�Z��O�X��圊��q	[u;�ZQC3���A(��jO�1;��Ou��v;U�:�p0"��=��D�>��g�+ktO\���إ�ә��-����w1�\~�f�E�����7ʥ.>�_�b��#a�����4L��Fx������P^ 	ʾ��$2I��Ϫ/��L��\��s����Eg��I�F�8�4��	A�R�������e�S��*�[x\=7ؼ[��O�Fi���Ц�$�e�*��A����p�pU�BD��V��2�QE
��X����Q��\�%1���g��?a�L(�u[<�(���o8�+Bi%��q�1*9�d���ӳ˂���9��v��s�����:��%��h�'$ij;B�@�h�F,|�|�;� �85�8ٝv-m���+�����	J���a:���D <�H,Aȯ���7�姩ؤ�[�&U�jY���Zk���fULw2}�dޅV+�'���fI#�����Z�Q�K�$��D��U{�+�6(��>����4e`l�{�c<h�i�=wa.�+�����ݵ��۞�����B�a���P)� ��.��
G�[-�H(��2����޵%�;�s�>�Neş�j�2L��,���s��i�x��>���-2�oA���ڏ���7L&��b�5�Q^��7szc��he`^Rp�|�b�A���#_��Q��23X��s�Ș�B�DẂ�є�4�8�$_fd�9a��x~�Gv� �9��@���?l��	�xȚE5���A���.0�"@5�7�EM�F�](ټQ��[M��eP�0��������Ա��\" �VO{q�ۿ��ɕc%.6�Mr������D��#�l�q-Ì�!��s~ү9��GK.ͧ�6ķ=����?�^+����؂�"Y��ȝ������{����@��A��=C�yO�^���#~��MhiS�;��:�po�.>k�Z������{�_��]�~����}�1��s�ï�Oͫ�2�̉�彗@��oEٱ8G�.5�@Q�H�,��
E �:L�f���w��?�-��`e+3{a��'@ծ���B �J8���p��R�DLAj��H�,����%���Q{����$ajŽ��C}���gn,�@���
#��&p�T��� �<�z��WΊ.�NU����"��Q޹�z��e�N+��Z����d���༩b�a�Lu��ѢNrg1�+􍀠X�n:W�Φ鹫���a���MÄ�	I���t$;�<���i�Y*�����+����/��=�E�8)�u�Oӫ7���8�z�� �߂h�}�){k$A��{d T�P��6�R�j�b$H�܂��l]�,�B��}2餀���@�w��L�8)��[R�uy[b�g�7���/>���
�7L�^�8�%h��@�,���[�$�SMm���@4� g�b\ҙB�;������[TL���\_��1m�}8��Bq�Fw��h-�?+Uo�˱�+G�:�%��9��p�/�C�~��*4!ի�nQ�_E�P����=�N tݳ	�Y�<ˉZ\�+�U/R]-&R��D$D�0I�!���JN^�'�Ui��ܸO����!�Si��4���iWf��l_3��j�@/�j�_��#?Q��mv4S
s�U,����a�M���(q�y@�!�G�p��`�O}�B�Q�ıX:�S����*eI�������xdWT�~9��{�O�A^��]/���2r{5��Ҁ4#x�*8��n{��)����*�B�
��t��0h�o�V��0n�94̀>,��D��(J���D��S]�}��;���&��	�����\<L4w�&����z�@�;r����h9s�ҿ�!GՑ�xy�X̾����	�=Pͷo�~�]�����E�'���LA�cr��}a޿k�&ɴ�B꤈o�g�u���j�>��Y��N"i�L�a�U�w'k)h�.(uC�O��;�'��u	Ę��ύM(�F��/v�q��*�!,�8��=�܋��v�o"��)J�V#%?�-���M�����)�F��b��L�V�On:�\j��f�c���DaUz� ��
�Dl\�� �2wpJ�ٹY0�\�A�r��Y:����[K1$WX�%1#uh�<����k�v4l�W�ʟҨ ���f���%5����Ϩ]�;*#��hЩ	��j[u���s�E�[���ۄ�e��8�S&_�y7��M�@_���Kq3+-�Ƭ)�&Z�'�o����a�68n�#����V��H��ѯ-��3�xr��_7������䳵�4=���<p��M��d���5�T�",1=WeP|M5�.�nNYS+�X"�^�`�XD�Gʒ�]l��
�k��������xW3��6Z�_�_	�qȢ
S�� ����}����C�Ph���ʿ|�R@WH�b����d�`��̙ ����v��kB����I���M�KN�\�P_�:rߌ�-���n����tbh`5�q?����ic����e�w�r4��a��e�O
}�ʴ�[|�d]�xR��n��!�Uh!I�q�31����.9A�Ig����&f�y"�
FI��-*Z_��yTj�no[=���d��V2Q��z�5Gf�@�`1j����a��L�7,(�-jո��e#�b �s��Y�Bf�$���P@�������fմ<�pr3�P��{���^�SIS���_*f6�b�jJ�aޠ4�g�f��
.�LG�D� ~��g���}b��F1,�ȜK�$�K�R�س����߭��O��@�@�P�h]#�/T��@F��C�fh`o��ԁ�^G-a֌���6���F�=+���$a���ko d�k	
�EA��x[�����g�ֿvV
	$�I:/ ]�^_�O�:��<:|PU��ţ�]	����U�`�)
Y���oE�MSO����k{��'}n"%h����(VI�x~���%%%x�/8?��lg�/���.Z�s\�K���i���0Fŀ��X��j���=�oq��1*��(]؀ϛO�e
?cen�_R#��2 ,R�wE ��>?����e�U���D�SFγR�X�6dx5x�rj�	��z��P�Ȇ�D7xaRZyiX�'�8A۱�)&�B��r��>\g(K��%x�u�f����D�GOrj$�"A��R����%��CP��
�#S��J��z-0ǂ?m�۫�&�V��yl��ÔzY�A���h�-�A,:zku�Dk��<��	c�V��q�8���5� q��f�*B�kGUI|F㪗�[�-T�
�U2����|��<ȆA��}Pd�#o��e`u�+.��,r_8[
�sk�C������4�~��Ga��ƨ���&�u����޵�=S�3΀C��ͣ�&�Oa�Ũ	��_Nst���g�z������:;/je7�(z~ 8�Lcm�\�8�>��#��A�m	�!�.��k{��a�)5��j��3i�,���V�%���pRM&�+�v���$U{a�Ŷ#U_�,�rN��eߤnT�o�	���a���'D����/K\b˯�MW(��"{�&����:Òx�E9W�3��]��UG��ڈ_z/A�9�}�)x=ƕ��%�#�8�x\'Pǫ>�hӏP/���m^�u+�0F��� /�m��ߔ��EVX�4+w���=��uߌ>=�q�3��"�T�=�*�H��V�?V���(� w��+��w������lM�?0L�O�#u�>��vjZ�e2�r��I��A��=q�d��1�<�!X�ջ�\Ƅ�֝���=�Z��i&9�<� ��!DA]��',�l�e5����z�"Q���uL���(�(k24.oV*����N�+��|sct����Lc%���̇������ocoV����� ��)/�叀�ᣲ0R��s(6��%E`L�g�vA�,��&�=x!%h����Ξ2�ڔ���x%��Z�h�h��4�#b%�:�M���>ZkC9��k�,>�E	\��f!��#�
�e�"
��������.�V��|�tu����,2S��μY@{�������T��M$�_�{������qJ9����&�G����k}�O���X��҅ә�&��]&� A@�@�J,��`s�����ċ����Ї�D3V+SV��l�$�5�����GA��%�Q7B�%媨�����>��&�E)>4�M�27���$0Ր���u��g���\�o8���K]#=ȱݪ^�C�z��D������x4ŝ�J��;���߰M�s�yu����6$�t)A�E,CVja���� q��5����k�mn4�j�i�sW�Ļ}�3K�����C�:����!R�5d�Z!"Ô��3���*��a�c� ��q���Q!��}�������@�9���e&ъDO^ض�d���6�2�3\Y��'yߵ��l h�O���5��ƹ�����YDQ�^!���c�I)�F�|ĿR<�'����S1"꿯e�E���oxvs�3y��\9r����/��=��ѭfn���%�=;�����p�7�,N���m��R�73�JO+s��"6_��ü]0�����.�-9M���x�9
&v+1!+u#F�˭U�_���n�<e�Х
kO�+?$�|ޞۊ*|R�0��/4̼ܺ4�B$���uvIa݊�ǜp��`��Q��cKƚ�Ay�����D�9I�y�Q�x�ܞ?}�Q��C3��x_]2�8�<eg�X�vq����AE��>�n��׳�부���T�m&�2��q�������}�E��u=ٵI�g���l}]/̴l��ݙ/�5)�%u��$>$���&�u'����F��%J����"�{}:��������������ҡs�,+�v,� ��0g�$�Pg��V'Tr����r��G��0WL�3D�$yF7�����<f�P���i�B+�YR��S�+��s9g�y@%�����������$��&��L����^!��`r�A{	�L=�8���C�Eil�҂�\�Qk���φŔ4�H�X{Nއ�?3�X�ׂ���������G�a+�4"�ik)9\ߺe��mAmq�+��٫��R�8�T[ήx4��!N;،����vk,{l�)��z"�����_ߘ�����삿7р͔�{9~H�Bwv����Ok��be�"�qh���T]o�_�!Z��V�!qr��4t����轀�C��P7�{�~]mR?���dA�o�"�7O�q��o�C�9gY6�G͑֫�Sv���k@m3�.+�	����� �|k7�gu�=��߈�s`��K%AI�U��{�L�(��X҇c(0��n��^Qgޖ=��U�su���HE�-�q�Ҏȓ׮�ϰ݈j,�~�M��%+�["�O�#8E�(�^�'p1xx����w�Ӟ�
}fup������tB���N�+&��]68+u�/�v
.��� �.�k�w�FH�V�����"������>9Z`�=6�M���P���d8˖͸�����#<S�~��À#,r��*M��إ<��l�ѶE>�
؛O0qGv� �v8���L�=/����$���3���-��"��@	��mŲ�3n�r�ώ�(?Q��Dv����������Dy�eT �n��{{�8è��i5R�D�����$٬a��J��Q0wb�F	*�8�l����I�q�����@4Ҋo�80�fju��?�,:�E�I�"�����h�tg�x�-	"l�9��O�������JZ�Y�Zh��+CC+t���C�l�:�FX��D����Ԡ%�_I����XQ*)Н.B!dJk%,l��ۑ�d���2H�/kpl�5qu�@˂�7�g~I�n�Dh�?�Wq�}[���2e����@��ā��L��T����G�W�D.>��|�)���5�AQ
����UL^�+��$P=fj6Ո�P�؎_�Dl��Qs�`�I) ��n(�<���_���R,�-v6�>�T�t�?�'�О@���+���� fK�uP��W�k����
�ӈ$��Ʃ�B�L2I���&�Ԁk�B�Ƌ���or��dǱy�0,A{�#����Y}bgd���^+�q���d�WVѷG��6
5�T�Y�Kj�:�3����2[z_��c�ߋdǍ�\[F��}=Z\	wS�	�I_4[��S���U\�s�>�;3�k�W4�=�5뮊�eڢk��|�9�Y_B�}��z�;}�o��]��Oc��NB�2�2�<5/���|��Ǝ��=�_�涏����^<�L�/�#�";���������k/��l��C!��q�c��xv��P���!aQ��&q[��_#QYАV�Y�\��苍5=������tϤp��<�}�����D��%׊�d���SE�?����c��l�)\X�ga؃H���Aa&���΃,��>�x��&<d�vڒ&�ӏ����&��*��8Z�� ���ַY@�=�o�_��ۙ[������r.g(�vw��N�6��_.x��r��>�,~�T�V���<�U!{X�/Mu��\՜�>�U��+���T�����v�	��|4���1����)�W�.�N�DjD=5ɣy+9uU���T�ǿ
}�1�]�ez�ή�b�F�܏���p(/6k� �}�U ��݄����K��}��P����Reߢ�����n�`t�����9�: 5����6SŁ���ͯ/7�f<r�yF�R�N�����A3�II�h�"|0�>�V{uQ�4��[PL��d���@�kʵ��V�+c����#�yR�V���+�Gz��.vu���^`�kζC�@�f��;��#��S�>�o_vs)��$��D�&��!}�1}�{�8���$)X�Q������AF�CZ�]��A���9�l�1p����_��)�W�4���>�a'���[�׉���'XL�m�+�X�?������r$�ˇ�x�Q��k����h�A�x�D�)��0�L<��tP�t�w��:�����9�b"LIA�%�n��CR�t�R�>L�/�������dj��`���?�d�O�ق���%�P�L"�� ��6�Q�5�����_��|l;a�#�����=L5=}������(�JE�W*���	�_�[���p�:5�oڅ���0z�~x����ɖ���+lT�*gYS��l�Ƈ�b��Lo�!��v���΂#���������~t&���bH;��R�#7�ڹE���j�[�Z%v������j�\�=!��Lf$[��2�پ���D����P$��`i���~�vk����>�9a�+,��I��ze?邑7�@
~���s�E`��؃��u��q��`Y�h9^�1��#�>���铽�@,��5>v'���_N*�|�e���L�Ö#wڿ�i�>;�*������@��6[O��O�i"o^��C��Hj�P�6����X�q�պ�CI^����0�^J�4ڴ��~�ڧک�*;�VQ��dy\;
?�&ޑlޝ��exu,��g˿§-}o�?���֝��hqS���ȱ�B��Q�|E!��s6SǏ����zZ��t����as�; x�t��]�<}O�v�c Bb��z��+~*^���4��zҗHכ�n���
�s盩���^y����,6���FtH0��Vz�a��5
�k��"�0ƍBD8�?����t��WW$��2*B���i���Ć�%x�9
�(s(�׮?C?�d�n9U�Ԛ)���`�l��36�#!El�H#�{��_,	bF�n�-b�/�e�JU!��H��+ �Ғ��=�%e�����DA����]��nO�����d�1���3��	��)�Y�?��t4U�	f��A�P��;Z������{����4�v�-0�=̉�iF�	n@d�zm�5��Ԙ�kQ�M�!Z�B�
V���
Q��p��n��l��fnl�ii�ȔثmD�bǊٽ�nȑ����js[�lT��8���/E7��~�՛P{����>i@M���qE�^I��Y��#�7&�y��AX �����CE��P�zc^u�y���5&m~"4�����7vw,*���ҰS[��U�V:�Q8ᖯ^\�jy���m��x���[�2�&��4�MǁI��s��1������e���M�?����ND�dX)9�#����HQB�'Ơ�A6zj��T}� 0�ly���^���^J��Cd��s	B�j��4/KQe`?�b���n�L��8�-)��^�Ǯ����\��O(ol7�A��rV��xt�2F��U)����i�솥J����v{���,��(�?���g�G���8+���Yp�]�~C��]�t���hM��Op�v���^b*.�A�����X���h�)�O~�E6i�[;Q#�oY�h�����n�8����(e �$�>/�����B�"��3�5�	���'}�yJ=�����b퍨ȶC�����ntɧ#p<|�w�6�jeņ�I\p�Y?Ǵ���2��f��&�Fݢ�-c�{��:����B����}�/t<ŀ�FAi�����*��X5D�@ ��A�	��G��q���߭%��1�5�r��[Ǖ�t�h�o���"TT���	g��ǐ0�[3(�h�0��t����)���5�����(�������eE�(��,R��,�0�uǵ�(�wM���mi����~��H���Յs�j�`�W�86�ݎ�?��U�`i���#�~x���wwY�ip�h!:@7��E�G2"���2��|�)�H���F�6���P/.����:�(|�ƣ��I�+ZN�2��ؚ�~��Wv�4���E�x$0�ՠ?��|T�'İc49m�w���t�B;C�u3o��]���@y�k�v%��I|�Cy^V��p�f�U��=�n��,��`՞#39���J�p{�f$f4�;1S?Tls�L�;�VfkU3^:tB���m�!��#�`I���<��p)cڷ���y��pp�xB�����9��^�H&*(��N]\K�X3���x��^���A3�4���Mk$���۰Y����3�pp県���oL�v9[h���"ꨓD6��Q/�顾k���3M�ص����Z�^Mb��
�i�	W��$��-Ɇ3��M�sF�|�|_%f~=�L����(c��b�	��A��>�Z���n���{3*L����9�e3B�cm�ܟ�Jjr��h��L�
KA���&-�n;"M�jĦ,���'���4Fg���G�#��}��x���R��
�8Ȇ�.lQ�V(�E'����c*Hua�f+SZ���|��=洚�|ڶ>qq�H^]�>�[�"�;�8��XX��QwN�M�ɢ�l
�B���<���UB�b�b�B��Sz���Wvk�����*�k����
`�ƪ�_c4�!"�2nH�lj�2�`%t�J3�"L&у���t�	 2Z}�ϕ�K�/,b�����qoI��F��

��		������j�Y�h>Ye��|�P\���w��Jw�3�x;#rPVE��o���~�`0��������%r7A�������=��5?�NGߙ�!"�|Uј#�x�~��	�3K�f��Ard>5Y��{'C��Y8���Z�*�/���WR�w<�]Ģ�Wĵ5����40Y?�VBA3{���f\��MSUm��/�I��@��gG�XK0Ix��/�t�a��1�y_M ;,�?�=
4��o����-��lQ�{I��I"��늈�U��G��jܰ5B�n�K��혰f壙=�x�o6q�ɰ'+G��S��ؒ����P����gL��h��I�E�T�I��9�QO>����y#�i��[%c-~?��������7.��=����=�}������K^���]��u~2dl�y�Tn	��0��uNK"��L8�����GY@��X���πc�J���:��W��N��t��oQ�u��Oq��<#Rb����򥀰��xH�-���Q�Yո�ʔ��R�6I�,)_��r�˟�
��8��9����o]aK�;VX�d��tnu5K�%�<���)��@
g7xH�
	�����k�ؽ�'��Þ-_!'B����E�q.�	���Ʊ��k����x�)d�*��`���KXT��U�bp�.f�ME=�De(���&���8�H*+88跁��2!���y�m��u�U�P"���@�m@n������M��A,�T��)�sZ���t)�g���ޛy:��!j��@ܦMX��$c��o>� 9������ܱk�=��<@�pf�3�c�I�T��㖽���Q��_o� v�����2�a0��K{�3{��Y��l�v*�ʾ�5����pO�`w�G�Wfx�{�M�=�<�?�y�;:'K͚��r��}�}|kM��A%־V'���,���<�B<�q��-�GK�aW��+����l������k� J�o`��UV����l$t�[��9��R ����%ޛ�(���y�W1��ﺜ\{Oq@�^��0���e�:p-}ۆF)�V]U����s�_�_�)ݹ���E-_����,lj�s�*�����,i�p`���*U��&^���i���(rm�Ɔ�0rS�|�h��D7�g�׼��WY5�K���
��ymձ��30�͡~e�԰�"��y5�6T��e^w�7j��'�R@��i�T�C���Ү�bP�Ǣʎ�"d���_��9%�:4߀���^ ؼḱ�T����$��D���_�ٍ�xm�֪�Ȫa}s�O@���� G,���p�vW�4xFa,�z����aQ�MX���������5z�O�3nHycgg�������S�2uԿ�d����9Z�*�U�jq;����p���'���0I[�%�p��������{�T
�g��\@��]���q��>�+����g�֪��E�]"N�2;���&Ѣ�5�J�yj�."B���dv��ً "m�w�a�c�y��囑)�� K�mӵ��%�#[/�����~� hl���3rE0
+�Ig�}�"������S���i�3%@Fn������,T`/3ۛf�!��<*/Fh4�赣}4?>7���<;M�,���`���=<FJ�:Q����g�T���n�-
�1�`alNw��%���d�n����|�mF䨳htU2\��	��aZ����.TA� �M��JI��\f�r˾	��9�@7a`��·=�}.�%�y#��C��U�5�Om+ʫ3�a7�B���'�0��?�����qӗ6�3V���5'�H��X:���_�����G5H�r~�0[Gsqk5ky@�h���~�v��_(syD�#b�XL�_9�;�p����b���,Ŋ�c���u.cI��M�M+�t�� ��*ӽ�n�ɴ>~�_�R��������~����B�`�B��� ��*�9pu��z�Z�6�M��^a�X���_h�U뷎�͍��B!U��Yܗ�x��$�X��ris�	�[��#"�^I��P��H���W�X�O��Pєq�;nLfE����
;Gr���͈�#Į�Î�J��R��y"$Zn(`'��"�l�<X�J��͈��ɶ9t"g�$f3����_�)�������=��Æ�0�������A"���
�?$s݆s5�Wf���,]�����s �E&���,W�to:����(���ذ.i�48���/�?��,��.8�m���/YgTW���Q�T�ӆ�xΗ��E�L�H��WXD$�f`��Y�)�=|n�h�*��\q�03���HwsH�y��2�2���Z��,A�/?T$��tq���>���g�0��f��놠���o���y7��t�OM�=O�����b��٥U�!%�� �Ӱz;�Ġu��A%�ϣ���+Z��z�����C�)X���0���M~��k��eꔤˇ�8T--���C�q﨨�W�6h���_��4���Y��c���H"�3���q��lxG��g5���*w��'��f�$a��Φ�6_�'Q_�E6�{FG&�&���>7��*�t��ݭs+$�᪻(���y=�ӭP��_##f���Iz	I%�Lڼ���؉�ɿ�ۈ!���{��`&�N��c0�X����\�{W,�x=^ܹw	d��츌V"��^_��� �Q�Jm��D��5}I���R�<�a��=�=�x�X�C[��y�/���7�j��\�l/.�٥�)��`�e�@~�v��m^�$ҊsTf�x[Q-�xK"k�/	)Å#���ahի$��y�~����~���tA�����oZ�11���vS�q�[�+R/x����Bږ���歰�aP5��kg؂�j�5�s�-r�!}w��]��M�g��_��=ʨ����JK���J��u�4TBd�$���1�p�v��wal��ro{>K,}mAN}�����#�/�2�}T�UA��γv_k'�2��#
���BN�S��-��KU������[�ן^&痧�2�Iw��T���	*'��>�TӀu��6;v}R�!|�^FVI�����n�>S��^� 1�!�oB�3��͢��2��-ɜ+v.SJ�6�D�Y5����h�|T�At��
ȁ1P��8�\ne�#,y(����0İ+�4@}K����%?O���?æ�܄�E�]�vd��NAS
;L5�v8���5g�?\����!�}Yf�u+	���1~��z���i#1�Q�-��o�gy�Һ"u�`��{/M.��[L�5̰�:�OMY�h@�q�o��9u�su����4µ�"��ui7��4l��vt�_ ��r��2�tx������(���hm�.s�b�I�J���@c��¯>�GE��d�ѻ?=%���-�ɗ8@d�~��sX�l�	Elt$E9�Ud�vL�_���̏<c�7j,�M��C���,Ҳ�̉#���̉u%Z̋��F�����.�?�>rT܏���IU�ɝ���?���1^����H�sJ�:I�.o`��Y�ި�{����b.0B��$b7o���?�i��Чaa����_9WW�P�iП"�(6�C�&�71҆نiy���n��EGc���A�D\�y`^
黛��,����ݎT	�+ad�5}�4<����K���ң�	"���������N�ky�vQ�lp��v�wz��S	���tߝ��,XS��]�|��,Z�1/����&���`������) 6����.g���%�8��R���w8Z|D�_þ��P�OQ�^��&
r<�� I�y���5$��������wOE����*�,�����cA~��Ƈ�@y������5_�>�3a�aw�4��Wl���ڃn��&�{���ܞ��"���Ea��\��OR�� ��b)'NC�;�7�`�y��"���1��f���)��a�@��1�n�Sߡ�_�R=hGwj�E�X�}����g$rQ��!�^Nd�������z@֯�fH��g�\���՝{�s��QW�H���B{�c���o�D�uZ���X����:��I���� �͡�w��0��q%3��$C=@B��t����=?!�i���cp
��7g�:QE3"Z؟�$F�٥Y>C_��5F�y�5oTE�sS �_�u�ol�(6��j����B;��z�R��Ǆw  ���V����l� }��Hf��ʅ�zy���/I��Qh�m 5����E��r��T�U�} ����EM��J�u�5�F�%K�O!��4��jխ��������0������!�9
������p�G��D,@=d.|��LWW��<�]��q����C�˦ �3���n.%AU��ET`!8Ŕv(��?�s�kO�0�����{��
6ZJFV���z^�ΑŚF��6$������F]ʎ*Ӕ��k�O #]!4�t[D�Ȁ㶐Ђ�4t�KR��FՏN�Q����[�ĺH-���W!�;�&�fV�-���y����95,5�\�"-A���\�/g��ݳjK�����<��e�{kO$��wIZI�=ֆ<�%x�烅@l�Zm@VTc��3����q])�8-��^�M�=P�<,�N+s8o�wz���uʌ5� �n�L}��{�i��qO��!C�\�_d�'��9���Z��{b�{��q��U*�$~����y4�%�!C:1F�>]�F��)��uι<����Z^�Ȁw�zē���sz2���<} �j��ؚ��#�vQ
x���h����-q6��nN�.�]��j0��^ՙ�X}����Z��Jޫ.c�@�0��Az��Ɯ[�:�P�Ꞩ���L�%Va��
��)� GN��ל-�`�I�M��&�+W�:���~�s��R�`)�u��3"�!\��V��Ax�>�)��y[	pٌ�e�5�غ��gR;\�F��ſ6���R�(^w�0�Y|�#Y5�ZIX-���b����ޒE**����i#`�͛Ia�%���-k5s��h~� #� n��59���u�( ������f�<��ϛL���P�r�D|�HT���j��f��!2bV rG�p`�9�}U�a�_�L���И 8Ҩ��)��%L��Z_#e���>k��S�B=R4�*t�esA; }�fđ�\�/hK#�]��K�[y��!=d
������|	��&�}� ��.2�����ouT6u�D:!1�RVr~N���z�3F9��e�8�
�g.�H- �a����fZ�`��cmCQ^�23�O�l���bE��I<�AqD�	lu���sRwc�����I����M�pAgu�4l�`/�U�����*M�J���p��������)�U��F/pŦEk��2آ��9򌇇�I��\0-�QD���Q����0�b�Ar����'�Ǿa)�ҳ�"�YTS�rt�Ӯ'��FimΡ����B48��Wa�-&4��;���&ѲI��%Q�5ӍX�@�5Oe=<��}_M�`PہmRt-�vH��J�5&N�7K��SmOnA��i>��'ԃ3{~i�S߇�LO�C5	�'VW��C��RY�L�iHSæ)oH����j�!ʌ�4�璀
�|�<����k	G�[
����KQ��Gn�	Z���;
�m
��rhh�[���R寪���hW�`f�]ҭsR8��(�X�O��r�8�JM*y�v��R	�m_qv7\��+�~�{}�L�$j�#��� ��P��"�|���;�|h�N�W�1���g��Q��]�N<���ҟyҌe��v�����dS���EZ�38ŕ��
�=��S��v[��6���n+ؒ�ɉ����|J
�o ��
��y$�\h�dk� _��6�xM�G6܍^�s)�B� �)�%ym�!�B2�v%쩏���p��GJ^Ao_*���b<���Y`FJt���@�w񊏂��C�e25����\8�j?���/��vD�_=�v�9�%�6�a��b��Q��CS��)
�`���/���P�.]ʟ>�[�T�u_�v�x����� $[�=�tJ ��� #�����%�ӻ��av����ta;i��N+\�(B�@����m��H�����%�0�N-�)��B�o�(���=R���|j��{u1�#���%T���F��ÿ�Z�� ���1x ��q��xd��c�GV��v;`-��Jh-�T�Y�-Ֆ��k%�㵍كR��nE�%�����N��}\}��J2�s^��P�Bi7�������-$c#�O�(@PnsER�0s��k~�ܤ�@!��M8�f���
���}�&Dr�͘�?�F��,��_��|Vz"��8D$E��ApX<f�zD����e~l掗�.�@�9j?�@oaWN��9d!��S�#�F�u���\�(\1��N��v�]��VgȶjsǜQ��dhB�/	բ�O�8W�(1��Wy��v�{-қ�JG�F��r��e �?�$���R�
FF���"Ѿ��QH�9V�?���".@�;��]zc�Ѡ �ȍ�W���.7��|�.y)X�~�����;&�S�v�h*���q�rh#D| P ��.��,דWy%�!�(�T��� tb��4)�>e��N�@�-���6 ��T��}+xdQ�-���&895�UP@�	�i4�)�I!�h�'j�]W��6D]2F�g�e/aS�<��5����,�=��3ǆ�y�im���4b �d��'~��i�ng�ˮ:I�)���'���@��Tk��t��x\	�r�O�j���F�\�X�����U0@�/��q�"R�9X�dR��́���)h�tӫ8I7T1/�]!ӻ��w`sS͜��A_,��tW�v��$q�v�}��K�C%�P耰g|���A��m�a�h����P:q�����DJ`��/X/<�Ȟ��s�yZ�������?rt��J,��~������)�ױ?��?���"��&���6k� �\5�J��L|�/��C��|{�դ"�'fQcK��y�W{�/�*�c�0`F_����������r����a���ek��֊sTE� 0JJ��14��"�px��
���qf�ϡ����ʮ̨�}�݌�|��ċj�4��tұ]���|lLBJu���K���Dǜ�,����PN¯r��-�r�^�3���n�qD(	�(���|��f�꒞�MA����ލb��*d�4���J\B�5�ҧ�,A�a���k*�Gi���]��� ���e�Ũ;t��K5`�� �gx�U&;�M�z/i�;!X�!�m۵_�8*pr�Icڈ�kFbx��K:B��e�9փ���6J,E�t=�]��T��p����A�W�P�U:�vm���sM����4�0@?�4�j�qk4�j��|"㈙~��D�t"�A�� �<g����D���}��Rs6d )0�r�m�S���c��\;�����C"�·����S�܁:.�l�r�,��7h���ւ��T���"%�����5���B�~�}������.��*�)��kR��[1+�V����R1zc��C�u��_�a_=��X�Z�g���˩p��.��q���	�l����ύ.�z�%����o�#��"�4gG��e(#'���:�=:a)���/����8^��ϒ�.@���qwd�\��1��cH�A����cm� ����{��DU�ȑ�|�]���8 3��I��xZ0��o�n���s&��L	 ��cv�L5�����ڢ5��lI��Va)^�"��Wb�S: �vO�GhnSm*��ᩋ�����%�'�yRU����	���1�^&�ꀭ:��q���Hz�#A�:s>�
��<���=:�n���o��@~u؞�$�N��������9���`�4ߒ�I4,��T'�]�N���a 0v�VBȪ�?�Xi�����rt�J�'X���n9"8��n�v<������a��S�*��pѵ>C�`aW_���mmEw�<�
�j#�1gO��;�k{UV,�k;�}�G�������;;���8Q;�2��65:�:��F)�9�m����V׺��촺�%M�@׋�6�D�U���՝c[菡�wX�!?�W�quhx����!�L =6���~��X�N�[�=!�T�����r�.uCs$�%mc/0J�H���'Q���	��
�~ ���LwlZa�ؗ�R�����pL�ď� �\�����s-י�R:;���>��rJ���G�`M�b�p�N&�s ���aJ�n�4C�z�1f�4�bK�*~�R��� ��p+g]nK+([�Ã`:�@�"\��$=+;/�߳n�+L/�g��L{lշ�����d="�����=������0���];d�֏�)��(I�:ׂ��$ͻ��u��-0d�z&.3Y���n��@�1�����ê���$MǴ�H7Ug<.L��2#U�4��ِ>���ೢ�zx��H��r���xШ��F�����7r�c�w���{���I�Hb�y�"�m�K�8���
v������>jm*��he��R��B��3�,Ie�c�!��R���A���-�*�^3&��Fm�Ԑ+A���_#-��بuEZa���$�d��~ִ;o��)c�~��`���x�U`0����P^�ncnV�D��T��ZQt�A�ѷN���?e\qh��z߱E-8ۙ
�F�Q��Z�@�qE���w	iR�o(��}��p9���6S��Mg!��r��*����?�|g`����~a�,G��սV�����!f��}���W��I�\
���t�(y�x������wab��o[qx�^����2��ٚ�A_E���F�<c������,�
��
1M@�NUMm��F!�~��!��Z�>MS8S�s�D����ڤ�uF^�˃���`-��x�A9�P��� T�
\/I��,��C��ב�&�Hd�7����Q���ChX�'eY�y��5�ͭ>�|�RM��GDLXE�>j��t�*��.�p��E	�ҝ����k
�
+2�N�����,@���oFfE%��'M"H1/�j�H�D��OQ����io��D��䏑2vFRDYd~Hb�� ����ۖX���.Ը�Q����2�33���!=P:v����0kK]`E�_�V�
PE�/�n�������e;FV��Cy�����\ u����hI�U�\�{՗�:��W{��k�NT��H�.�_2t.���[��T�a�	�ʄ@�({��Nl<��Z(�S+{]�1n�W�`"�h/y�V9������Y:�	V�S��A2n�%d(�YT�k�J�FM�?a���^ŷ}�[c~��v	��&�N�['��z<е1�#T�{�#�N���%<�HV��36�z�3;����m|���� A��e���4�ŏ4�R^��<��1�R�x���i�K5���%��Vr����1hՊ��#ۧ��R��گ��Vtb�B��	ϣM�M͵����FK�0�P��R�ۇ�t�S�
cm��~���uD�������=�$|��u�i���u�E�#pt [�i4���5��]�+�B���b!�/}��\`����,ei?��
Aȟ'`b�ij-@�|IMp=���U
��\����DQ�4�}-N��L�@y>W�洃t��ƜC8�OrdAco~����蒘�=w�D�է��	����;"Q Gg�,����;|�,vN��G�<z�I����B���[��-PЈ$v>L���^��8ƊLf�'M�mD_��Б��`\��)`f�lc>�i� �?`&],Ƞ ��<W�S��D�_�|�w��R$������w)���<Q:i-qϱ�y���
���*�^藤���D�n�=��|-�,tT�u�{��ԋ{K�2�ǚ"B�v�mzd�T"�os����X�cl��2���P&���*1n_��5�җ��˝���������cUR���i{c��E��9��Ž�������z�k��i^�ZgUt���V�L��W�N����YH�5�N��sfhU�0i�S��}&J��P��P{Q�4b�z���{7���M�.��M�-c%� ��Ey�I�"2G�G����J'i
�5HL|�vn�!���Y�o��Zf�h�(=b<���P�	��H��Z���a���bP�<���\2���C_Rl�x���mdަ�/�J���X�VWG�Q�>�?CX��IX���	�}F*��=�҉pL��I�r��@���.�@(�:)����; H�Jz:Ʈ%� �n��jR)�8�H�P��,O��i�	�	f`��:�����+��T���&��)Zݣ!C���� =��&��m:/���r�K��H�K�]���Š* ��z�z��!�0o1
�Tk�f���fX)��9��RfJ��K:2�'�0��%�������@`�J�xL鉳n����C4׺n������k���cPf@���گtDc���Ze"`�(��Is`�(��3�~��"���9Vm _�Ѽ�)�md���-2�:���B�1zk�\W�׷Sד��{P�aI�hV̞�v���DC�?(e!�c�}���p&Օ>�}PNݮ;�U{��7Cæ<|j�(����}B��D�:T��ViOi��Oy���Ȝw�̊��"y�c��T���E�j�P��H���L���=P�o�_QU}����v:�e�|�6;���,�AVrH�� r�*���7Aq૥x���]W�\Ԗr�vvxD��˕k�`��:�y��;��*̼�:��hװ�G2b����E��'g��>�<�%�.�_�{�{%jX����t ���s3s�w�;櫻���9`��u�>8�p��	j�Δ��p�-�e<ZM*#��b��8�w��͸Ʃ��PGO5�/^���j�ʮ��&��z�\�2Iy��f� }�*�jB��_���q��T��"_D!��le5�z�!!�4�wfm�1����R)X�'�j&2Ѓ��O9��]����8�j�$n �x�/�,Ue���j��%��ǘM�<�q��QN�m�:�{k̎<�x�ܶ�Tx �S<^�ʇ����~k�O�<!�;�mګ�aơa��S],�F�l�X:RR�ʦ5�]KQ
�<k��� g3y����V,R�I@1�$/ ΍/f[X#Q�M@3�Y�X-?��V����S���O�����GtW�� �.�g*%J�Wl�^LO��3+�����_�&{0�$v�����vIB��=cF�}AmZ<p0�t=N�?aJ�FHP�&t�`�u,���Wq��׌�VzQMc�����
�^�P�
�|�ȿ����@���:�i][Z�i�[�$�䋥N��k)����-9%~���p [� ��>'?�t�<��ٹ�O1h`�x`F}D�+�סO9�Ԃ�<w2S����Y���_'�@���0�����LR�i�.�z@#8�+�i��'�
�C(|R��>/{UP��]��Q�x`d�Ȗ͊�һʑ_��pf����jHI/��x/���.|k�!��c]	��k���RV��wD���b9	DD����%���w����U�c������YE�0u,�L19�ٲϲ�>��ػei@��{��$ϭ�Ģ1�T�HKk���-`(�x���!��P0� �u*+�*��bQ�l�,���B�@ނ�w�g�~�K�PR��x�i[]�0,f��=[= ��܁��8�GX>��u$2��Y&sC3�8R��ʶV.(�蜦b�z�<�0�W})o7	���͋�~Ƙ���gv�5�)�ѱ�=@��gx}��S�V�m�^��e c2�͆+��q�G�ɦ�D���|TJ.�#�o#��j�q�h	BL$$$UC" i�������B�!��Pb�*����Gx�c���jQ�K��;��M��'��^��4NJ�c���#�J���S~��4ۇlڬ�֩�Yt�,��*|@���]��A��}*�r�Kɢ��]D�CY��"����´	��T�V��Ni٫�l27� �������h�=$�e>�+���dF~Q+����B�A��F(+����������wICW�A���>2�?OԻ0�Y��7��Y)�$~)���ꘂ�"�&%vq_�*�;�_t�I�a{e��+K�tn��Z�]^�^9�!�Uu��}�k�a�E�-wH���F2v���{+ϖS*�<��h� T.�U�W��P@���u~�<�	�l�J���,I2|�8��c��������˕u�fuj�4����˹Lz��E�!����l:�Dn����A�(aT���
0�7�~N�܎p��`r���H�]�򂩊�jY�F�(r�vb��+?��k�%�7#�YVE-c#��#�����_�e
�p�k*B�!d�>+��c��U�b�Im�O���m����(�V��Ə���W0m��EK�=�\K�X�y09 la^V�̻�Dz�/ma&�C_0���=}�=R�67�hB��04�����ѫ�{��*��1}�\&��Z�9dtZ�4�t�x:.����������=�W�:eLl��|�DS�%�0*]Xd��\��_�F�|����'�(b]������l]=	��D2]Ř����,��v��s]�R�_3Cze]������P�>_���d�>�r��9� �q��WW��׵�g��r���J n���O�淋2������Ǐ�ԫ��	$��xi��6(�[5��쇳c7��w��1�ūz��p��wƯ1����J�[2:-
'C���(�A�%�R��4��b�ӏ?'�"c�F�U��q�_�%N���Z�Mޕ�'x	���_M���6�>����|�`k�it�,ݸ�)���녙�(ŧ���ZZ#F'%C�<�~�u�o-���/�4m�c���7�qm�L�9���k32OJ�n�,R�DR�ܿ)���iU�FŽi�51�)�%�����	����@b�j��x�_Gk2�� �;�ݬF0��*�y�j�OdI�x��T�MQ����a,i«��&�V�8�x�A��ki�c�^C�<��6�������g�-G�l����F�d<��3|�x�z��������&�v>@ �|^�6�mJ�򩄆�<�ܹm������4�S��5R?{�0!�R���=�� $�����?U����^OE�u�KQp� �\�~�V�RP 6}C��T��L���M&���,O^��orʈ��[��6Ș��V�\��n�tz��	��;w�L�Ғ�P�UFC��"�vd�!q3����lذ8#�]��+��m6!��)o
��vf��I�D|���!�$? ���3��:C��8�����A�rTQG�0T���q�q<�d�rV��E�Բ5�S$=�h��;_<�T��>M��v�9��N��_�n(Sp�Uf� ���\��i������=���_���H��E�`� +IC�dH�{���^��8��A�B{�x���O��VFg���:i��s���Y���ފ����E�����kc�^��H�M�
��[������	-��
��]�j�&DBE��C��PoQ���㹒�;�2{7U�=�s�oX���$ǻ���:�w��v)��إ�>���L�qe�n��x���j�>�-��Ꮐ��.w'��C4�v�@ ��t�D��
\� J�=ϵ�`���C���$�w'���|O����
��K�#ìy.m׵P���o-��T��\/��us���E�����<�r,�-{�Uu�_:!���	��(�88�>�i�N�� ��)����#���ڭ��dB��i�:s�%_�C�٤����`iT/�Y��=[��t��u��Y�_y��w_J����w���~{�l���o�R��c,���Y�ۉA���&,�O��)�� ;,u�D�_�L�!dyh�b�r���c#x܂�'m_RXq�P",��	m����J��~X�&f���o���d�S#�̓����S��L�
�^�a��-��ud僓v[��n�O
Ab��1�S�lU�F�o*�mq
\o��su�����j�:��Sŉ�à�=��G�2�Z[5"���:��C�h뺞�`c�a!��{��O��#�fg�@��`��g���]C�������ҟ��A)j��qJ������u֢I�"� �z>��<�*T�7�_"а�L������/ �G�U3_X���d)����Ҥ��2,/��r���>=���ፒQ$��Po�F]���]�%�rv���y�O��s���J0�1zn9���=��6E&�S]NR��eⷱ��������P���Q�zJ�� �Tɖf�F��ޜ8�RN8[�J�`@��}�� �������F��[aZw��EG0�V����-K�3�&��X*{�k�6hQ���tK��c���D9D��rQ��.0�����>v1�#2B	$� �dz:�+㴬�RԢ��S���:`�9J)��,�mhD��gG u˔ ��վ7%�S��v9��ݝ8�1?I�����;x}�l|����k<_L}�z&�ҋ[��֏�&-a���^�ދ9#O��"7��F�2'y�,P=(&�r����9\-Z�QO�ز�J�a�_aǢe}�{��]bD��-]V�0�c.��,\=��{�q_������D;�n1z)�c
Q�1�F����	{Gb�Z�m�P�WS��<��'#A� ~]����5hn���U�(�>?GseoU�'�L��%��Xc�)߀:��`��y�6}��d�l�D���LPT���4�v)f���Au��� X�P`�*,I����o��:s�,�w���˧UvЮ~%��;�U$k���-�����S t��՟]wo��GN �-=K��W'Ծ=7q����O�QDU�Yp�d��.�Q⨥�DH�FK4$�f����X�A`>teE{8����9`v�}ɧ!J7�L�
�K|�4?H5=3�g谻�q�?����`��o/[`��$���t$��d��sbD�����ӈP�xŚ��B�@&y"����hh�����bQW���jw�*���1��K��g2A���We<L߲��7bMªnS���֦Y@B�V��^L@�o�=�w&Ciʖ9���FH��Iz~���1='+U�|k�X��\��ԧ�bV����UA��� 4T�!���3(
@�q
~��$�`�8@øzTd�J�>�:wTq��R�d�s���aK,�)��>e�4t1�bҋ�X}�%�B6�T���
h��ʩ������y�&�*� ׯV�p �)&�����}N�{�Fxe"�<�3�\�Ӎj�`Y)�
@t7OT�ʠQ13��G�w����c��ҥ���=� � �7?�gFB����<HhY����;r�<���f�(��ys���U�����K�oe����IAbU�:blB�mY�W.����}b(`�\~�U�_�߿x�z�.���y��R@OC~�=N��$!�#(~���Q����?(c�u�=�r���#b Z2
������*v, z/�L}��)�
�>�;�O�L�*�Q��؎�.����]�,�>oP,�%����s�q5�ĊJ�Au�=�\$2��p�t�s8�D	��yW)�6O҆�Ĳ���g� ��*t�s��R��k�0�����9f����b����H��%��5]qH����鹽+�R�L.��86OUFp<��N�F��	Ο����t�<)���=���"����a	���t,7PCK�jdm_�nb�##���2eR��T�n��w9�c��@������v�Vڧ�C��.Kz�^촍��+f�E��J�	�Oӱ���A}����s�� t�Fx���]�&-䮛�8��t���t��F�1���s���P����\݂m�H��5�/�T�+��c��}��X�>�^Ȍa��a4	Te(X1�X0�{	�Ƶ�@��{L��Gm 	�TX]5��\'=�Ug:3��\ʺ<�7�ף+T�1�Z� �vQ��w�P=�:y>��Ħ�)�mVg���,�xc��cVp���uq�	�LV$�8.!"�0�E��&��,E��E�iz��BЎ���:���>c^U��e˷�h_�
a]G�t�����-�=����u�n�\a&}��"�tl1���LlQ/�T6o��o����ٴ�zŦ��%/�Շ;,8�����=��؅Mslz˶��-~E� |��1�1���m���B'�mNFO���6c�p"7:�G�bTJl\,j첼jج�@��K1yR�s�;��՚��?��P���U�l|��m)(\�	
z�yP���Ʊ�U���1�|�4UfQL��t�]�L-��s�Β�P�>�9=�OӄN=���l�}d���'c��1��]/�ko�ں�Z����	�M��<����q�
*P`�I�[�I�~���D#%"����'�4�@F����9��C��O2�_2���Q�=fK��0O!�� �O���nG��▟��r���'�Ϸ�G{���8�HM͒�����:Tй���)��/}�)�g��M��%3��}��vj�E0��h�������[��x/�զ!?���V���̏�n���N�FZȓ�X�s���m�S�`E5��	#���D��z:U��6K#"9£�n�;��h������8������p<A1��.�,%����r`�ʉ��J�����GȲ��
�z�w�L �K�W���t&<}�
?�b2:�#��j�\���~8��p^bR�N��9<h���˰��ͧ���aB ��g�nC���M��8"��R�]=+,�;����X��G7�/��R��Ѱ��xZ�x�ҏ�cS�Hq�|��jS���jZV	�6�>n)h�� M����rڐcצi��S_��	��q����'���P^k��Tư"}�[n��v�f(�+}���7���6���]d��N�G���W�r� f���3r�˗�����L���s��c�@�5~HJ�ĥj�-ŋ8�T���m�$�� '�gFA(��K~�ڟd�m{�I�m�Bk@���)�r��E"��BZ��`��5h�e�s��b"���}��T˞Tܸ���;ns��(���@2���Uhг�A�s�V	�2��(��A觞Ojn�����[*�䋾�'��z��x��C����L���q��D��+�������a�<�vQP�T�?$�E���VB��W���4�?�E̙p��
E�-�sk���v��T��(�CN��g��q�:7�"i��.z�Zi��o����c���{�}���܃.�A��f�:��V�顨�/�C�_���p���w귗y�=�_�a�^��6�q&DWa�:�6�.Hr݁^�˔�\�lJx�P���W��K��~�%V��,$���,@I���k�r�����"��
字x�z$973����JZ9r|�GK�����0�b���ȩ�l�i�k`ߛ���oX~��#���^�oU��r���^�&����:C�7{P�΃��~�oK�.�48��V��U�eo�r
w4>Zm�Q��љ��~�\����4a���#�����	u����i/��ǝ�;l<_��(�nfz�x1�~�(��D��/ll�'c[���b]�hYQnB��.^:;Ni���N��p���q�J��9DƤ��\���7K\Su��W9�n��l9��~M��[[�s�-��~���*�/�=���Cu>+�]���Ǔ�S�/�����p����]�bs͉�9�#�@^��}*3Kܒ��`� mwH�O(��L�>��j�kp��;8&Z=L���51�,;ļ�#�� 5�`I�矵�%V���e`��.��-�k �YF��:+��m��`��9&r� �}X��7.ƪ�)f�~�0y�sQo�:���3Ft0\|�=t,��@����r�u��H^��vo8|I���"���B�	�$M:<-����J|��C���/O�Thb)�0��DY`��y�T�TW����m�3�Y_�?��-��S %\���!I-��d{���N�{�ݩ��= H��i(��]t��Tu�$^���3bK��?�8
���N�']��J7ߛc��1]���sz�^j�P�hs�.0oŁP ���ѣ�2�t�X0�׿,A�����.�\�+��J���@����vL3^`�?d5��pjs0�	><��I��J{�1T`���7�����{>$�#���Ş�<�U�7�֎p���@V�����{A����d�~L\�tG��`tv����Ĵx��W2�XX��&�
��J1��R��a��g�J�;���T�s5(x0��<47�t��&��'��!3B֜���9�0��u&����Ф��o)bj��E���Ȉ���5wͫ���|����-�������A}�/s�6Q�4��Y���A��HF��G��Ԗ4>��,bȥd�kJ;�f���1Nv�^�B�T��r���9d�D�NW���.�y�8��@.m�n���nѶ���b�%�o�祀<v+�b�V��yf�9�c�Z���O7��#��F5�;��$, �
Xq9U����eӄ�w{gA�⍚�0�AS�ʹ1>�ڌ��M�j�`�_���n�& ��[����m�Ii6oʱN�K�ȸn���n��t����;R������{�s@x�4��`y�%� ����u�}V#>y���M��������TToڟ\n�tkЫ�b�@s��6�� Y;��ދ4l$��vm��(�Tܔti����ǒ�RO�~/!�kՎ4Ƹ��E}yj�h^n�%zE52?�8�+U�"C��w%� S|����߾�q� ��8 6���UF(�aY�#�-mp��;[�]��)�e�����3���O��ts_����|j�
����#��+1.PE�%���֤;�,�қ�
�ȧ��������M���R>29�[~�m�R0�����ε1��=�0��V�i�'��p꿶����RQVY�[%-9��d���H!O��x?+�e�!��)�֩/�p癸r���;�������D�;2X�K�����Q�Dh@㻊�g�.�8'�㋌���Z��0PU��.$�81��(��^�h�Fl��ȇ^b ���f�"J��IC��~�WW�^G�<���i�}�n��D���^��'�x��p��Yg���~淑n��%w@�E������$[�4��1�qZ	G��ׇtCM����<H�h���E4(ғ
D�%r{4$�;Z�.�� �Q�b'-F��Ζ�Lb`���q׼��m��?}o�a^�3�����}�2;��TA�%����T9�;a�Ƕ�ڿ'�K��h�dR崻���܀7/]=\&�>	�5�q�;B�·�?�⃟o�>i�EE$�c�X������G):]/��'Ahm�(͢��=� h_���(Q�������������J�����joiY�<�
�{�*�@�j�Ք�,YI
[o��@lR��A;��M��Oqk�V�q�2��+�u��fa8 �c�ܔ_�u1�bx������}����~�Y��r�4�ϻ�o&Ǟ~ؼ���#�	ɷ,�ha�oj]+g˪̉.*��"�a!��gn��y�xKiB9��e]z��L��[��3�7��o3D�T7�6�jgv��zύ�N>�n_�P�pQ��N�j���w��e&-!��-��d��K��dJ�a`a(��^)�M�`W=�*_k�,$�N�hD2�D��d� Mc��|�0�����'N*dٖ�����ʧ�i 㥇�mb}YX�����}� D �}��R�N��}m����8 ��I����l��N�jDKhU�h�Ѣ��h�<�F1���R!�|����շ\AD�eSa����p�ԥ/.!�K�͛>JQ��x��
@�5�d_?��4i�~�3\E���o�W�S�-/�G�N��h�+��/�ED�{�AV#ٍ,��|
�n��V���lw�Ѭ��~1�TԒI�����J���r�I�wf��Ish����>�%��*vq>��HG�
n�g�D�R1Rٳ�S|��_�����=N���_x��ZMIS{Cs	W�p�N�%���b��࣓����*����a�����9���Y� 4m�	��1jy651��ң���?}
P�lV���{��#��m��8i�D�Ud�u ̲����:<JI�z/����� �k�|�(��ǔC� ������=nx���& X��iOժ�ѯ]���]��M.��v�!V��B�ɓK4<�AN^Ko	F�{Z����au�z�����`�.���ӿz:�B�,>�@�UC,����fY�]����??,�	&��C�I���WG�N�te�R�6��t��fn7=��y�B��ҟ?h}�6�f���� �kV��
�=M�L�*�ԝ�i#Q���C<�r�z�	�Q �9;1�@M���
ut�y;�|�z'Ԏ/��M�<s@��ӂq��D��mm8p����1nCs�v<�MВ�檍�L��i�ͬ�C����+ )�x��s�����5>�ɲ�@��&��C����4@��. �o8�̔�FB3.+�ٕ���H�U���,�WIi� O]c^�M,���׀8�HY��3#/�P����W,fr��)U5���js��P��Ț߯�%���I!�㗜e�/��G�#<t�kL�������'��m�j�U>�>x�NS��aq�j9�m�R#��)5�r.w&�'�A���_YK
r6���'<��m��EZ���1�i_�ֆu���S+��RS]�D>6��ﶜ㿤�D��.t��\+��6u_�]��gm�D��7�G�7��o���_�j�1Vv��.,a��og5ʧ�������E�0���wű
�AZ��=��Hx����D�2��P>������PT�L�`��ti*��SK��1������.����Os#��s���Z�6�(z�$��t�o)��4�`��;[���N2�����RX��!��2�9��u�!HR�iP4�ydrɇ��C]��h/��3Q�!:h��.������
3� �D�	�sE�?����_f�Gp�>��B�;� ���%��/vv����LF?7H@18xJ���#w���S�e������V�x�n�f4��l�UswJ��oW+�E��Dz '���z�#1Iz B#͔��M�Sb����cf�x�6.��'FgLzw��F�ϝu��V����%�=l���BM��/�W��6�c����NS�=�*�x�6EB��_�^8����K�o<���~YY;H�Jǈ	WJ3h�~Uyذ8��"F[���Э�����vș���������z;@k���,4��ïK&��qI&��A&�T��
t��~G�T��\�����h��
��D�N�
����d<Y��E����C@s�%{f����T ӿ�R�?T����� ����j���+n����$!�⦓8�g'JS��� g���!�g����*Ûr�0Al{��v�Q��nͮp�f�s�t=�-3nY�r�Q��Q+�kY�V����s� -��\�7 h����SY;�:��z���Y6m���zæ��	Y	�������< � ��dL2}��	s%�e�V ���y��n�fc^�>M�D-��I}�1�o��t�U�3.�y�O�:䫥l�m�=h���8*�?�$�~���W0�Ws���!A�j-���{&=�j�$51"�ua}U���͇����Bnw��Q�O�6��Ɂ�����d��Y�_d�1��jp���=Y�x;����WQ2z����/�u�-�d��'�iF�s<SA��qu�$6lX�?2�?'zP�v ��11 ��R4�=����у�r����=~�3kd��3Q��x3��nY�0#��x݊L�+x����'��+郐���\T��*<�&_�3�j�I4�~s*y�&`���u?������c����W�c,t���;j�t]Ѭ/sS_�p[�#0K��hq�"t���P��� �٠k��~w�g��8�T��+/w��t�E&���� ]�P1~QΟrj�U�m98��
��<̫dgPC,�)���\*�X(d3��;>��_�B�QN��k��d5.�o���^�0�YW9ʉi	�X�|8�W�̃<]-^��n��2g��I�n��	���.Ym�9xq˨52���k.o�-�������=~vԟ��6��`�}舫:�td86�������qc��U{��ɩp ��}6���60 4�b�^����r��|s���i�y�xe�~50 �eU/�OF�{�0�Y8�Q�զyĭ�*{�.;���|��	u��/Y/�[��W���9��ɟ-��s��1n|��yϻ��l�F�P*|G!��� p'b��p�9���5��'�����A�$�|K��f�B-f@Җ���|y��� ���ȶ~��v��O'����T�X�5��U��v�[���=���=�qU�] W�ri&Xc�dB������X}�:�A�h?�M��IrY�!��E̽� ��WO������/3{_&�SI��VN!V�E	Ց!�y8t�5���?$�>��S1Y����]^DAA����KR�
����5U������˾���!n�;�c�S�����7{��P���vg�����Z��G�o���`�+�o�B��;dK�+�`��=��'}?,Nρ̿8�m���q��� ��"����Lrs�M�=)M���6oɵ�En�fD���NQ�Be�u�'��^����[zc1}B�9s/��o�X��L���m9r�D��k땻=���I} :��Vz�'g�_���@���o����>n��Ÿ�s��T���2̠��*,P����P�9�S��C�R͆Ä���O WBa��,t;�y`���Ln�ꢾf8�^�Q�(S��M���[�k�#_9C��Ӿ�ˌ��囓�fo�~�!�o�XT�"�B���v��ab�XfsG%��azy�՛赊`&Uv9}��_y�>L��6el��������3��$��ֻ���x�*zIc�*YsA�͏w�T��|2�Ј-M�׶�]��4����M;Du��g�p��R���홗��K�v��!�!�S���(Ugw� �%rK���lѼ��Wm�C/��|��T��ca�]��h%e��9-k�'(s.�+PVpdY���_�{d�*~�֗�k�I*鋻�@� V����cW�#A(ēxi);�(�qG�,�����$KK�1;�Q�X���g��ӌ��QQ�I)X��ˇ�b����*k�!��d���@p �L�r��F����U(G}�v{��/RI'������k,O�	r0{���� &��|��s��Y|D��^�'2s(� ɚW�.)���7����[\�)�%�a4���]��@�P��2:��)�I�*���t�"�UAr	���D������R ��6�r@�����&����]ۢx&���!��-L9aU��oz������yXp����u��7u ���� �oT�F�5�ƽE��Qg�S]��;�ȗ�'L�),�LQH`h9ip�մC��:u����'(U0w.<�~�3P�D�{�E7T�(O+�qg
�R�P�)�dIŗ)˧�X
�۶� Xǀ�Ne��%��|�8�Nl� k�Ր�W�Z�9��I$2�7l~<T Yⓦ=ob��S8�q������L6|0P�C4$N��T4�K��%B:e�����<)�/<�[q$���p)O��v\�qU��A
�9�<�Nml

xœ���
A��	���@v�1�c��骯��1����q"2)��������;���ӻ�D�r�u��-ey�"�=F��� j(����N�x56̤��E[1��AO��ܸA��昦�ٻgU��@��7Y(E-+*��&�fwIF ����(E~�-���M�UbT�᦯���3����o�QTa�"�`{�lQ������pf!<�\��nƒ/����xG���sc4�� ��Q ~�j?���uRfԨ�6��F4�w�<��o�/
�R>���]q�<tS���UY��zr��D�+������$����*^��R�(]sl_]�k|k��^.�N��Yş�2j�T;�����L���K}�n�|�6N�����'sZYp/y㊇H� �֘�Ǒk���9��/%l	��5�k��=&�l��Z�l:i*+$�v�ۀ�vK�ϻ��Vs����o�L� ���,Lk1��!V)ߓN���җ�;�=�X�J�����P�zm/�dX� k�+P�$ܮ%�i�՞5ƈf���o��)@@�L��y�S�[MO�˻l��vr��z��@A��� xhE��/�%=���R��w3��Uiu�����zf^���^���TA�`ܞ3E�Z���$[���SiV���J	�O�MX�������^�}-(���.I��EfWP�=Z܈���D��A�3Rh��-$` �BE�%�;�^��Z��bf����m��y��:vD����K2��d�򉜫�Ŗ�He$dʣ�_�;g!A�?}��)X8�]~�!h�$c{��z�Θt&��W�?648j�41,��9�g�RE���<��[����R�(������Pa�F�Z��;v�/�8%j3�n^h�`�X푰����������l��&�K�S�<�5n�]i�ܱ�A�7�̠>iZ�`)iz�z��B �{��7���I� �w3��g֡sS ��_TwVI@>4��A`��$��������?)�G��Tj�S_�:Ϻ�t�^�	E�iU ��^���  �]�9�$�Be�*�ƽ��V�ރ�y��61&��peٵc~�cE��)Ձ�q��.������1�����Qe�k�9����Ê��ˮ� �D�̙��:��<���W�	��:�h%�Z�l2��-����|em��uo�wM�O?�w���vQz?�I���r3����׊��r�ۼ���7�K�Ǥ��y�_H�����K�������O����#r�,� x'�Ք�|w(������,��3�Ct{��6�m�b�;o5�9��0�o�	��Ѧ��Oqc$��D�E��ܮ*,��s������}][m���,#���f�� ~�bhծ��ƌC_v"p	�8��f_��)�`�\I�E�_�@_N�rXp�}F��uuXE�D-����8�d��uF5
��ZZÜ5�_�K�'������ճ&;���)Rqx��a�_L�v�V�[K�/�ڟ����&x��}@��P]r5����~�� 6�|ߪP���� *���f3a*��B��`Ϲ�KG�$��lix��;W2�S�7j�0��q�̚����瞠e6W��5����	ǆs��6w5��U���\~_����]<xnc(&U��zpމ:��(��tv�NO���SU��>ݟ�=��e�C���"8-O����r��3� V�1�=��6�m���f���(.k/���\�; [g�,a��g7�u�3?M���S�w��=�r���C�r��A'3��TЈ�Re/�#���Pi��槝�<��r)��N��^u�����m'�$b!�M�����khZ��)HU�ۚ����]P��\ p�8�GKKk�m�_-,X��tyx�����uv1D�����:�7��f���#4I����9�هQGz�(�F�S��ˡ�S�222I�$��YV�2G��{�y����w�E�Ē�-L�d�EΏ�Q��H�u��Z.�����@F+��0���d��0=��Z�%y�D+l��A�H���h�+�=��4F�V��*S�q�JF�]
�Bʞ~b�Fv??��$�w�sI�%��q3�^��oiTŅ"��H�&~��1����c�A[��w'L�r^Υ4�*����|c>�:Q���%��x�������(ѰgH���v�_P�}�M)� 
'P�H	��R^b�3`;a�v/L���ʮ5�'B��Q����߮5��h�UQ�N���$s�A�S��,s���\�x���.CV��u-w��A� Ǔ�Xx�_f����&{OZ�@ʣ:�3c�<�"[����E�0©��k�9NRw��[��c��LA9���Ϙ t��v��XP�h؝ 5&��j~S��Da��	�p�A�����7T�5�(��d}ԋ���g	sF۴�R��	ٔ��: Ԋa ^�1�^�����1���1���`j���F����������`�}���ą+(����z;{��}`"�`���P^�1~�µ=*�:��H��F}N�a�ˡ'T�vl'l�&�Ѻ ���z����3�Dz�@Y�ܴ�t������<Q$H稨��l�2g�'��9��럭��E��2��S!g7I�j�M�U+CE�M�u��g�r��
�u���¨����r����.�j�~�.��~�Gb�8��b_��J�4P|Ϋ��(�ڕ(��*Ҟ�&b���??
�OLk1~�3z���G�(Hff+c� �袳���@5\��%�� O�/a0�K�^��y�G�Sb�������>V���m#�$3"���~��\&�����U�����6��hŔi?y��2!�.ere#��L�����n���^��;x)ѤMOC����);��z���oQ� �jF��R�a�.i�ך�Y����vB��
n�D��%7�?�/А�%dW�O�}��x�U�ڏ�mS�Oy,G�[���|��'p�Q%�6����.�{���_L2Z�Y�2	���e�
;'�S�Ly�sk�f��X�C͘[	���(���^���L�Ϲ��ʰ6��a�f�^��BA'a�C��/�@$�����?�Br��=��e^W���r�q~�L"-�**����f{��r ��;�,���n3ڭ��8���c��I����Ib fG�(��ŋC����5>	��[�r$Q]v�cg�h���+=8�5��Ĵ2���2";
��9�J]`�l+y
�1��[�d�D�`q��� ��!�̮���|����g�js>�Lc2�[�~���v�ޠ�8Ā��)��ji�뤊�Q�mi#�lD R=ɶw�
;~	�°���8W����z��������{ �T0*���N��[�
v�BԪ?�3��x����8�V��F#��R�d�އ���!�A!���ė�Q�[��<� T�E��$T�z��<��İ�I��\��7ɷ��]��4_�+HW�Vq�\�	��1�o�m��D�4�����|� �h�o��X���s�4�>��(,��I����i e��5V�P,�cI1�bT���q��P�i?X�U٬))=����l���UT�ծ��[�����!t�8F�L�3Z:��U�/F����~B���ԃ�i����^�[j��X?0b�)���m�����$���w�9��3��j��h��j�(:�M~�J���OEC�em���%?!�h ��mq�8�>���-Ӫ�O W�^���6�Z�x .���(���xm.��%�g���!ŝ�So2�=ge��&�!�Voˍ�+�UOXߓ[۫D��pt�CH�i��b�ψ?;�>���d�R�����P��Ë-�Y�	dE�"	$���.4W�I��S�Q@(����K&�"8�+���
�ܢb���t�����u�U�2������>u�#��2�"��f9(�y*�,��YU�~!7�lN�yLLw��l� ?�q3�[�/����Л$��#�+��#�����M#�8����+$��i���4�>'v jӾlf���P9�'ui�{-m�ͮ�g�X�$�՚��?���K������Ap:W�Fj��7��x�]Y��G��MBݲ�2�ʏ��O�	b���*y���b�N$C�WW�E"ʏmH�ߌ�w�8i���0�+�Eۉ���R�s���bέ1Q�,���$f�����=v��s��n�G��{@����d��<�D�7�x3_��US��rm��鞃ҭ�U��`�{1�3�6��0��r[n$�s��@�t��6ē���3)d(�tȉgy��<Hṕ�g��`z-H���um��g<���W�,��0mFH
Fz��M;��@��Êũ�K��>�����{�k(g�q\g��K��*��$&�c�K3��q��z�׸�t�#q�qG7H���-��,{ ��M���u!6��� ,QTeR��:l����$���}�|�??�,xE��>�j���r%hP��f�wI���àVR_)�r�?�l.����/��w��Pj��_�5��-kL�U�Lͻ�ޖ� ���3;{��&���G!t�4m�@6���:C&��d|�bu�������!Н-��&�W>�~������]X���� ��!��a�������o��.��S�9Cf�y���Ny�t�|_���0������:A�����P�����'�=
{x��arļ�ˣ�u��,�2�p�����%��x���n6J�����7�r��	��h�
�_��- ٔ@߰J�\-��*��P���b�f`K�6����R�"-Q�<2�3 ���a;34w"�9n�I���dg �7�*�E��$�qf.{�V�ҏ��-�O��5Vq�GA�'���b	ro��!� ~�E�+��A�zF)$��CL���G^{�օr�|sJ���3W7T�U��s�c�b�w�/���|�wzj�R�]�8�oThS�c��L�2Э�
Cd���қ��G��K�� qK��IF���yA�۱j�L�j�˟� �ӛ#D۳�*x#���뀀c%*���P�M�����:KT����jO��b�q>jC��:AyK�rY'�F�P>���[��3kwB�^�ߜ�ރ��O�*�{�`ۃ��k�v�`?�����[�x�U�;���}��;�� �^�k��̿��̷)٨�d7��DD�v�6�t�bWE��s��6�?���Jz�cRN�d�KK�㎹<�Fl�X��L�<��/�H�<�?ŅE�޶E2��r��Ujc[��.���@U3�C6��C�"�d��tf�~�:�i/9uRW����G�_N�=��1%��m���E�Re��p�ᵔ�[r���{�Xqa��N@��?�I3�t��s��6�r%�(�}T\L��0?mx�
�!��������E�!3�;x��(6�#�R�Z��-����}��O;�)$$�$F�[~]�¤����>�G���:0xcZ�HK�h��M���У�F���c���<�W|Ǽ'�O��䃳l�}�#2��nd<�S�J�(�$���V2�¢��U]�W5 ����<M���F����Š��F��M��f�%�3tf�E�@SO�/��~k�Gy�Gddp��,�] �D5%��L�c3�5�)s�>�����=.ic�).T�`%��y{��C��ԄeZf�X3 �WS���f�����:�����f�Vjŋ#�J`&z�0!N%�!oH;$��؇X�6kP��(��]�A�����U�9�����/�D=��}�	�5k���&��H���GΌ�0�x�z���)1j�
�W�]��G �&<���f ��x� ��5s9a�N
Mc����7*���6Dt˔F�L<����k���uQШ�=RCȘ�)���x��p1Rh��x��p�GƊba94S!��a�n@��8w9|Z�H�F�T�ؘ?%ء��B;PgD��P|c��h�⢹"�&&���iy��H��)OS�e=����ŋ�%7+"�)2���ÚH0�źl�w��p�-u�����V�!�����S���&����9���U��+3�UB�f�~ik^e3�X{�I��?ټʼ���0���D��v'ްU��PM���o��]�I���0r�]�Pm�p��GS~\�*Q���zQ��7,�N����M��r������fw���b�%D����5�g�LW%8$q��\�
����d�{�WՁv	�ެd�)�m*.�`w���Q����X���f�p^���A�R��c�p�3n�Ӟ7��&M��t��c��[���N�y
��CYy*�����@���ڹ��1� |���Ke ַS�l��"����Lb����]�ӓ��/yj�efvN/�Xf��Bo~b��y5��q~'6ϰ�!�4�N�fd�)LH�����q<��
G癞�����N�jŕ��Y���l�`E�M��MB�t������=�?�O������c#G�p�TRlӣb]Xu�L1�Fp�-���}��t]Cs������U��p�%��6��s��N]���P%&�n=��J��`0f�p��zB�s�E'�*h��Ib�&|�:1�Z��ٜbgN�� ���4|�]��jg���e�=&-���Y����[ QZ���|��~��.I�R�"qwO�]���8�ɲ�]E}O�h�=\��'���x9�X�@�Lt�:f$� ��G½���6K�/���L��1@a������)t�J	���r�/��T>��A@s�q��w�/]u���g�����/���܈7���y��=ɗ"o#IG%�h�8��jL��;Cy\�yfb9n��dy�wL��כ$�.
��2�-�UVfk���ܼS�$�%���)=����]��Ąt�.��p���O/�١��ͲwH|�"�S.�2�ē�=��YѨ؊S���U�M||}��~!