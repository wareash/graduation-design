��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|p�n�U��d�&�VQN4��'�_ayQM��r�oP�Q��G����o��`{��0^�1l��H�E�u��pɻ�)��w���tO:@�n�D:��8dQ`k�f`$��p���R��|�-x�?�/����T\��]�����QC�#�u�tѫ�*x�S�y�o������a�F��"s~�,O=V^��s��S���g�'�j����nr,_�;�-�T�!��>��2@( n���+jF^�d��t�J�w9���g���E�.������Q�P�k�2m4�2*����Ӻ��8���8���^���i�7*!�9�����8�2��~�6��uO�2�,y���}~��g��l�����ua���� ͚���8��
Y��r�mw�m�u�T�`�)ڊ{˚�{aD����-�y�Z������x%a����C/�0���!�mh�+7/d�o1�"�jLq]:�W��	J��`&��:,�bn�U�C����ފy�D��c�+�'�r�5C���Jd��8���d�סz�uW,�8�h��L<�&�𚯥��w�㒞�B��3�����������z��7��c�+=z���\Ʌ�9y����bF�����������ھ|հ��\�˴�N���ra��H2az]}�����4�Y�'�l��/�2��؏Y�r��j&7�r�ï��۾�L�=�/e�����mr�g��(j~7��	ۼ8h�;`�	r^�Nfk�O�����r]����������$�(���9��M_�����C�Wb�iһ���D�:?�����}�F���h�� G��OH�M~c��Sُ�z*d�0˗�9?5�����7�����?�&��N�t��!��Ho���I=1�at��8<��׀�!�z�l��,�ģH�����k��M�q=�j��An�5��C���F�{���[#Wַ�qEj̷�F�:G(���-pT��?��D��Ǥ�GR��Qa��z�����W�p�WzM�9O½_�+mh�6��"0�JuA�N�k���w�z�nfٔ�䈐��O��ͭ�{���dPA�Y�--����$�kԜ�Uށ���}�0dh3��('�{��Y#Ϫ�#/aW��z���[���2-9~ƛ�;|�1Ň��dq���V�bY_%�_�.H�t$��<_�&��Fc�>�	�zJXqhM�in���022^�^��P�K���?��O��~�W��T�Acڵ�v���{�o�-���%n5#����B�$��~���qF�����4J�Cr�f�6����a�8�}X`�_8���Du������:�6�u7~��9����+��	o#)��W��HK'�q��-�b�Ż��׷�+X@�_�Ű�l;�:0�����Xtt���{��$2|c�"�T��-�=MwWH�ފ��WS9��糶��>��&�%�����z&�j+�6��Aצ�P�|�BpY�w����{�s���8�b#�s��a�(�x擞�H{�_�¿�K��<����I�fF~@�Q���S$yݭE��Dc�s �!|��9�6���z�hn?�aφ5��]�3�9;M�]e #CƤ�J��o��^��)����)#�Ģ��)0)nMsC��@DI�5l�R�C6!�qF�'HH�9P�Бjϳ�|��Rf�7��pbR�jR�!	�����+ H���i�ծ��ΐ�"A�]�;��D�H��f�m3Eۜ>p%�l�]�Oz(Z���N��>�\����"M��U�n��1|UK� ��p�giT�^�=��:,�ϘM2��*��Ӂ�Af������T� m��_�;Ʋ�Y����f��,&-��@Tb�qqx�'������@?~��~I����ʌ��n��̤�vXcr�c������u/)�`���?����3��� �,�N9�a�l����5�V%�58��!�V�Ďe��~�N.�����k8<;�5�<�w@�rǌ
�9a�eӡ��IĄ\��!�u�ޠ�0������U�{ؔ/h�DڢH�LX��I�)����(�4��}���>��˲��$�[���`6�Gz_%[��7ӏL��YG�� ��$���uP���G��t�3D��kmr�t�>�m��1�{De1+�����B�c(���	�vkZ,t�D݌1��y�V�=�un�Q:�A>�G���.��?|	��t���.z�i#Nɠ��go��Y��ӑ0�{���w�M���k+�5Ag���Q>s|�؄4x� [\���b��1<{�BX�t�.������造Y�էdI@w�̵dˆ�xr2�����-�ëOp�~��Ai+���/1�;Uw��i�f*��ؿ��uhc��Y'C����aӦ��84�UQ^Z�*�ϼ��g��s9�O�n��U<����hB��ͥ�M��MhS���U�-�k�S��E(׀��z^$�;bƳ�m�T\H�tN�֮�]�ka���8�߀�ы���m�g�髨��c5���D��F���b"&�� *���y]b��A:�Q;W$�*�vTo`EF%�{F�R��Q��L>KUK���v�?��r58��ۻ �7"���(��:|�tN��Ąl��ͣ�4��Onw�lj��0��*q~nbN�v^_;bz�S�\�~���<�ȡ?�gN�������^��;�Wi�K7Gu���V*0�~� ��/����uy�m�\#-���u	sC&J����R	0��tY�"�@���X;��ny1�a൑�)Xę�)�]~�ZU[��ʊ8�n���X�_����:�ٓ`N�Xs����+�WRwI�]%gl��%���vL�8m�63��#9_u���{�"Hp�𷷌����{b2�� �P��%'x`�ۉ�^���R��i)w���V6	^ NS(�?���{��X��qTΞu1v�F�i4?�z�}��(#ff�.t�6��p�ͯ�0u���-���$�5��oi;CnU�S�v��"r�%,s-���/͑�dU���k�H�6��i_.!�}gH�O���j����GQ�HH��RZ��W����){ijv���&Bq��/
�~�n���;���bX ������V� h�QG�Shs�s���խh�	��D���?U��~CqF0�wRj�N^�~jU��ݨ����O`�p���q�dRm@Q| �_
�F㱗���(Rl�7�f��D�Vh'��9O�����X���R�x~�`bI�>p��<k�Rjj� 8�����.^��4���I+�H�s�ސX8ȡ���m.R��U�g�����Y�}�$�F!gnv��-�D2�e�V���ɤ`C�]Y,q��<j���b�X���#C(�},He�����j�^�(s=�i=�_�.�1-���q��-;Hۿ�'Ԛ�����W��S��4��=Ɇ��$�O3�3�$i�f�<�xG2a	;����s^�?�~Ι�X��m]RI��<�/�t�?x��(�)ښ+bt%0-�|!�i�K�3,ӎ7���BKk�%�,t�c��d�����T	�,�]�z�^B[��z�͋�i:s6����+��ؚ1n;�T�δČ~��B�luAg��^?���}/����!��?�6i�.�9i�;P5�0�$�E�N��E|7�W������$�{����|)��=��I#�[ի�;��l@gL��EUe3�iԛ}���g���>:���
&�1����ߎ����=;$�
h@�؄��Q#&>C!Υ�����h�jg�(W�~n��[����x����ǂ~v���?�������8����.�,���4`�^�Ma�͡�j�!�n�^�tt�?��y��4|�r�ipA��́b� L�&�e.���闱���_��2A2"��U�Ph�<�Eg0&�1�H�:���k�h��Y�,mg�������lx%t�Y.��i�_h����ǓFnF�".�qwE���n��D���b\�q�w7��:v�&��B��؎�<rE�{��>�'ր8t�)N�"4�DC�94�}��)	���'�����A>(_����/��C�-l'�[:��l��
<�����ޛ��e�W�>�����qc\hW��ۖ��+�T�JF�����D��{[���sh��c���W��
�o�?��+�I�Q�Sɨ�N�<�uC�wNR�ʆSf����T n��J6��d�I?{^~�i
���Cio&lz�IVh�4�ຆ�l��R���Нp~0D~�;\����e��w�.�%:zh�I�Y$�o4�۷C
�j�z��l؎v��$ �狗^dUWMA���Դj\��.��7o�ٿ���B������/���YІ]�����z�p%�Xt��m������>-�5��>wPU���-�Ѫd*�f�c�����*s�"L�c5C�vp��1vk���ZKk|Ԅ�Gɖ��<�!�y��/3���u�3�5�?t��P��t�����슢��H.c�	7H�VQ� "�Ýt��I� ��2�F��ZM��7����\;?�Q"��_b���M��%��&þ�8q,��F�eJC�GŰF�F0[�1�G��nh)O�v���a	M Px&m�yp�$q֕�A+ir��\z��<�j�p<��f�>d��z4���٣��r���*�����̫��';[��ڊ�p8|�<�i{$f%�;H�X�w��~��xnS#�ONTy��*���h�V��vc�3	c#��%g��NN�T����s�gd�Pӳ���s�������5턙����X�w�]0#�&e�>%Q��@�RxS�SV@�(@���i�(��S���da����Ȃ��ON��g�]|d>�V.�k�'j�_­�'�
���4>�ͪ�8�Kթ�"[u��&��I�'����s��E-���j�E8jn#��%|��y5�c�H�0�#>�fY�o����Z��剿��8��1��F��mGQX5`$�5.w��ݖ�@��&:QQ��O�Q|�WT�à���ܝ������y�]�wP�X�t��b(s�lX�>��Mt:=���^V�nN��E�>@lH�īoQ��R6cN�d��0����;�!�����+p@�@F�v�/Ҭ^��B>�P�]�WuSLN��ݔ��������I����ju�>L|�����jg��R�����ɔUT7=M�4_��n�W��-쓟�tT3ł�n���Q�"P��S橫���o.6L^,1����Gu�a$4(يY0Y�$�r�̨�e��1Y�E�N�A*���$�$�hښ� xp��9]���1���}���)��a��]ZCׁ�^��WmgKh(ù �4���W���{�/h�O�G�t�-ih�����F��{LԂ����Rc4�t��Fbb7G��K�z�)be�5h�'>�,�H3�Y~��b�É?���r~�j�G=������ ����M#z��A����KQ����(#�����#^���{�|l_0��E"e/��f�h,�9�'�����J�Nd��x��>^ba��?d�+�8��n4�~\oaNw� �x `[S1��Sˠ��U�c����Іz������\i��Q˗�`az\h���>�j��6�J�2�b�A�'�Q�W2Zg~����a׋X
~1	���6p�Y��s	s���u��\����!�!��]Dj�|'I5ȩi(M�Ӭ��<t;������K)��a���L��o�d7�1���U�搲��"������K�8̥��'�������Y�fS�.�?N'��Z}_�D!�=]�Yv������ki��`/]5�����¢ߞU}'t<b^@Y����0[���C1�&r5	g���R�v���Ac��3�빊�2\�vT�A��2۸8���/���X�x8�;�>��,C�tW���}��m�d�_b<�(A+���j��Ta�1Y��Q1�YZ�w�V���/����o,�$��'�R���갩�@;d4��$t�q��PF�D�2�<�� M%�����3$��gtP���3��taG9��XVBc=�*�xD&��,W�X�1����Tq4<�@�l|/gUw�0Z+$7�Ӈ�eui�q��sC��c�((x0�	2���}è��l�oF���3.-1DP\ �"k��+��ybR���{���%\$�*M�.�-��`��j<��fZphmIS���׳q�\�;;0Q(M�߲�#�?�?��.ʖ'+�{6&y�-O�:Ǌa(���*�/cӆ��a�(�1�z6 ���DiB�j���?H^>D�$ޭzP�.+��_��I �����?�e�,�[	L�� ci�R �. �/����;)_�7&aH���̒�]���[wئ�n�IϽl�B�!��^^ *��s�k]�A
�o(�sԮH��?F��>�!��$폸��e����Qͮ�\{$gK���CV��g���^������Ǒ�M$�}`��ҥ�2�����  S���r���&�?��c1B����D� �8�_=P`���%����00Z��kw�G�k��nXG�DO:��*��)����]���3����<M�\eݒ׊�߻�c[~U-'�6#Mo��V!�;-�t+�x�Z�y�Uh����{Bl�%�����<#�w4H�(��	��?g]��U.[UK��X���B1��yH������@_��_��pT�<��7��w��p��k�bܝ�~��A���r�&����*��k�)#P�'�o6n����$�H%">�Ƒ�����Vo�<�ʳ����>C�^Y ��Jh�.�җO����iɝ�od��"Q.ℵX/�.���p-p�+c�PT�q��!�ޮ긾ʇA�}Ih_�q�����ώx����)"����2Ri N����f�Y�%��m%����/C��Xm�1���)?ݒ/���	���/�K�h�WP���<d,�^e �kS�x@4��r�ƴ�u2�"��/qK�< ;=n���w���/�����R���&>�[�(�ܡ��_���Uk��r��������&���ms=� ��&T�^���v�@ʒ�&���b�Mm��%zz|1T�/ێ�RH�y9�M�9�z�㓐S��1R����YF����n��&�� 
��7�,�3�����Ďv���V�|�eBT�"B{=@��y��_S�"#Xlj����a��V�n�>"���&�?��D<H_�bC9VK�ѝC�d��=�s�V�Ϙ#U{(=r��O�?�\���i �;�W�2��m��Z��GJ��pD9�j۰�{;��?�R}L
�ꬵ����6��ͻc*�5aC�j��.�u:+0�fբȖ�1�K%�E�~2[�|Ǎ�o��I.�jK9kU>���_���;��q!�G��O'ҫ�A� ���&3�D��3�BHuX��챂�T��wT�ǢP�Rb���)ׇ܌).�KD�*'�+b�
��1ۋ@k^3��ӑk�ә��h��_<�x�ɟ&�4<|�	��Q�m��	W�9�beQ5:�B���{>I�}d�4n����5�G�	�eA���*�6rQ�mHK7�����&{P���{t>�^):���a�~���ą�5�{�wEg�fe�VD^�"*�YS�W�5`�iǖ�Uv�]��<��
�Ë�->�X�w����� �f�T�$�K���}����6���
�;ޘEEu���l4i����g����4�>�����	5��Ыv޲t�#��j��@;�`�Ƀ����j��7:m�LI�k��-�8�Sz��mXf�_KGY��2B�6����2'���&��i�Օ��򤞸�+��	�7ɠ+�|�yNb�Tj��:C�Sz
��ʣI"h��y�c�I�ŉu�{�~�DyC]9��M��;a��a�l;>�͟�=
L�9*Ŀ���1ݪ�?�DZ�NN���{F�S�t�ˌ�)�&�x���x�x��@���o���vP;�P��<��#G,5��7T���v*���	g8+�~ џ_��ƥ����[ ����Q�'n�V�i꒖��.z	���4�[k�����x]qL�����$�(�ÄKt����E�ݠ���hؗ�pǅS���t�J��cQ������J�����"t��c;(5�S�Ѧ���{չa�!ؿ���0v��L��Z
-�J\6���9<ƽ�<C_�z�>�EN-i�6ޗy՜n��zp�:�f���a�S;�J�11A���ξdU�������p�X#�{�w��<����B"����������&�Go�e���"����i?�f���TFS�cb z�A�����l��P��7ͧ�6��z�6M���W6�"|:�Pm�oj���qC��~x�/K�~X7(�����|l��?)B"(���ǫN��/�[ؐ&6��)-�VϚ����m���Xk�~ߓ�>�}#�"�L��_-+��^��\� ����3	;C?:�a�^vx�	-�8�笇-�&p���������#�&E����|n��06t�����p���^4�������H"���a�Z���Ao,�ҵ&��4�0�)1�Ͳpt}4��/e�_N�M��V4L����U�I×1�����Rcr���*lx���m�(��A�����[�5��w54E1{'��Q�',�!n�|@���N��%��z%C�\	��w�M�i�0qZ���j������]'\�bׅ���t��fJs����L��l^D��n�~Ǚ�Ta���;����M����z�і�L��(-G!�M�P�Jϛ���\�A�^�nFh#.Y������*���5ǲx�����8�h�o��Շ��3��)I�����[*�ځ�7�+*�a��$V�p���MUcހl�>J���66\�1D��e6<�R��f^���X�B*p�b�B��b`ӄ�i����������9����}�t����U���S��f�6.L7���
�Q<��b�<�,�L�@�S�7�J_��|-�m�ax��t��G�쐬���~�2`gB��}��C�~�	'���z�r��z�?N�@�x��fim��qRɈ��\�v ��l��:�Ѳ,\)��R�C�����\Q�ll��gZ`����x����kw8��㙌Q)���)���(�'l�k'ZQ�\�K|y��Ah��F��=Ǡ���O����A��=�	S�_	4*W $�0���^�˿��L�Z��<�su<�:}(�'� Ww�v�j���Fp��zH��L�q�#y�Uss����bð�6���4੼�扡��Tq�d?�v
�� �~C�i0�A.,�Nۤ.��,��9� �66�\�a�U�\������0�QS��'.��O�g��W�V21v#B��h��w��g$�q�ۨᨊ�ʞ�$��0�u��,�	�v�5�צ�*QfE�[p�!U��{q�ՁX�%��$W���>mN�u��+��CME��������+x�b���P��/��6E�3��L�i<tI���d���0Z4���cB"�6��m���/л��R�	�j��?7�v�DLW�;d�>Q�j�B���퓠��f0�N6mZF�/c�,@��Ǡ�9��\�S:4�`wK���XV�GO1�H�_u�E��g��@�W�yq����)ǥ��'���%�|F�z�ֱO�Bf�XU(��Ga�ZR:��<��l��]�s�gy��-[����VI��$*K�p��h��j�Ǫ<IǯS�p� nvI�:��������'����S�V �hl��3�@葮4H��|�;�~v�x�����j�$9z�˫�w�k�O-p|�%�c�#!��2f�5�]�g�DV��8v��;�
�;A9q��Lm��� ��P�;�f��K��b�7��#�P��mH�w�<�5�Zt�x-Lc{M����, ���o?w�M�Z�����.f���o��mf��&���vb��c��Uc��\_�@���i�7F�Ztt��(��A9���xt<��9jp1D�����h�!�~���K��95'��(���������΀�
�@-�,�y�n�I[ B #�� X�1nh@�̔Ζ��!3| �a�'��:��Ae��gp���\9��k#�g됣�
�p�&ۿ

�ִ/�ˬD��'M�A�41�f��y��Њʳ�u���5R��k�M�c��iY@1?>���ӃDJ@0�H ԃ��Ծ��g76���#�~��4����&!�(GQ 
�'�"G�D��jǠ���Й�����As<,��κ����K��@i�R���G>|��N@'H�Mͣ�N�=�R�CD{e��W�i�c�F H+���T�9���\1x���Am��	��� ��ץ+�����.i��RK2m�����R���0�t���&��	REsa|����͏M�\�H2��{S�.��-y�?9mX��M.�?���gH�T�Jv&-�>�kU��z'���+�`��`/�zX��YVZ�C(��~������& ߞd>�Q4�eU��л�t����S����.���'W�NL�9s5l�?�q���q�ԃ�nQ[O�3��l���f�s�?�g��`VR�p�9�4O2lF���6axО=�T=���yun,�I���ks [ZM*���c]$<N}���\���� ��:��1�=�U���{���
���Z�Ƴ��CЛ �^g##�BjX�!ݝ/�J����c��;U����%�&TRT�F}6����mN�T�抆��� �!���?
�{��P	�soWeS�#l��i�v�@��9�@Ҩ��`	��g�ޣ-}R����s��8���I�� 0�x�R�mJI>�S����f����ԺZ"(+�Cz"�>�t=��:�2��}�ݸ.v=���	۔^�<�JKU̸W�#FC&4	i2}�XcFjXq_���;Q��C�MJw6J�a�/"XbH��K�d�Ŗ����Ů��y2Z��%��S�����tU3��f���0��I���/u�,K��}�U�<��jw��F��{����	^�����s'?Ԝ�Kp�<���&`7�b-N�)�]�n \V6&(/��i	�
���[C��������z�df��r���<H
Yv�b���B�T��;+�Y<��9��+Q��hl� 8��M���!h����3��]�Zܸ���<ϖb��(�M�v�a�j`�@��lBc7tS�u1��}���~3�� ��ث���]I��� �#�zP;o���R��͢��)� �M�*�q�ڿ׾G����Ǒdp?q����M"
q~��<9�d�6ݣ�A�dYv	S�O?x�|i� X����?M���WX�?nP4fB'Ɯ�tu��k����(+���V�E��%�t-�B>J�6�2��USґj0�\�#Z��O�h
X��Ǯ�)�k�h���,gW�T�' ��&"��*9˺;����3��F�	�]�������/��1�}��&#�-��a�͌�5�ۖE!�-lc���zaa���(�ɚ� �A(�C Tu�]�Ǽ�h�,����)�x�.4�6��JP$$�7��3~n7E��񝄆�JD	DK(��M
`��jJ1������-U��V��g6�������h9e��Ф�Q����F���{��l���L�P�f^���]6�"vn��N�j�,����F�=Mf��Q:\�}��w�e�xg� gިV�wX���W���7QW{����ن�IA��2�tZ�vBS,�5m���%@�6蓇<L�c�(�?�� ���m8{a8�k=6c��oG���M�O.X&���V��JY�(=�݈�a��FRp[;��Q�����v�^xĨٔ�.��(]y��R��%�#�����������,	����v��#�7��Z�Q�(�����G���4�!�fÐ.+�^\7��̠P)߂j�����Ȫ��ڢ�)V����ڥ�ZȖ�ߐ�t)�1k	.%U0aq�X(��X!�h��O���=�fӽVX���eo���Zx?20���n_O�~�����8�꼬�)����s�g����[�y����DC?�G���x�P%�)8~M`K�k&V�꺦��`>ͿDT�����+�Ji���-=�g��X"5$I�~�ȋ�����Uk�kd�6Qp/��p6Z���'v��jAf�{�_�&|�ܨ�vܳ-Q#~�w������d�$ڮSO�=#�v^�%]V�݃�/�E�/̂҇�'~�跴�]��8�`���.C�:<��o�S�C��Ti�xr��4|N
�� ��9+���i���G
pn��x�%�#��wI]����Պ��������M�-�p*��?m��q�JS��Đd�Q���Cjޘ��ǻ�@�3��S������V}��"���g��Z��,�~G:��"P�ɴz)Jͦ�� ��Pk�'�]��p=������xq�d�"�!��o��C�Mʹ`�a��:��>��W���&G�7EE�2N%/�Ih0kFM��Y�WSZ���%�R��e`��LÓ)��]����}��-��A�sy#wY�c:�З�i7�˱��|j�Z�`NR.�e�������ys����s�";�0\pW�@ɔ����yD�߱Y��%|����г1}Jn�q��\�&}iL��̑�%�b�K�*�Z�@������ot�a
��A?�����AV���d�~o/��ˣ@����jx%�����N�B��K�t$}��2�(!O-�M�D�wM��`c��7C�{���� �lR~+0��Q��`�&�}oSG#�Iz˘A��1s���O��^�3�>A�qt�����u<1|=:ఛ�>�2�7b��Oɳ\��39ρ��7 �mޒD� �*tI�+b�N��ʬSIlB]�t�_gz��J'y�/�͢���p��.���?"`�۲!�%��t�*�HY��tB�֥ȩ���X|z؇���WˤДl��R>�k�_��n?�9���u.�\�٤�Lf-!_��௸�����P�!J��&��NUT@R{M'�Cx�����oz�	�^'�h��������N-єUZ��Ɂ���C���[�o�'���S��oK���j�.�=]	Ϛ����~Y�#�(*#�wFH:EQf"lf���%�R�##ZI~d��v(�U��U*!|i�@?<�'�~P~*У%`�%c5����q�=��:����2}������~�BY~CgЈ8�{�n f;�L��)2T��J��\��-�Rޅ��N�㝜;��k@,B��]+��I-=C��w�-��@�L�!�e��Ǆ7hw\��v}�gV~Q,To��6��f��~#*g�1i��ŒH�Mރa��)�M�T�9ω��A@A�_�-^ U�ǝ9P6���_�$�9�6`D0Ip��
IMI��Vl(@;�$����w��[-Od,S��� w"��|'<먄 \	�L\IUI�Ğ6ak�L�Z��S�u���.��Ÿ��[i��J;C��'�ek��u��^�^��j!��
�]pU2,._Dm�BV�BS"����+"�z��+i�?�ka̴l�� �ޜ�]���_;�ݑ! �-���ڞ���)��+"N0ӃJ�q|3����r눫Uz�x�["t�k��_�r��l�r�ed���{�J�T{��❠h�.w��C��0��������EX�:����˖��2��"!	�|8	���fnk{N`�mz^UZ6?y8U���$�6�~�ACZ�@m,�rr�?'{wUA���a���г�P	$�d�|�N�6])��a��3��E�R�8�^���rT�����-�Xed��0�њ�|�S:kֺ�:�:����	��ec�a���S�Z�ft�}��O�C�>���3hR���Ϊ���!�R�������}���:'s�Š���dSM��5���C]��0�K�6e(�Uݪ14^!ie|�u"K���)#:��9#%h���u��x��~���毌<&��	o�W���T`���a=��%�教�3��Y�hPE�.zބ-�[M/q ��>2[O�=�k�a#dU��}EXՠ�A%]�nMn2iR�u&s4�����t�9��� ��[�[��BV�����I�N���ϖ��8-	�����>���'=j��xsv`Ę��7Nx��E�]��f�eɧ�b[�{����6�nD�׿���"����&>�ߞ��9q��u�:�Jd��$��� �������31s��lJ���Y�� ��I�虷���mvnd����u�Ù{~����w���2���tB�9�d.=n���,SX�;��m�"�?Z�_q����W��ah�>u���0���pLФ|0�X�nLj��܆��#M�h'C}tW7���Ŀ�n��І�>"��b������p�X@�F�����t�����9)A�&CB2��_gi����[�R�S�="H�M�}�[�����40���mէ�B�=F��d�
�S�9p���D,�t�rƙ(�$�.>������K�h�7�+p�;=*���w|'s�	�m�J��Fu��@�b��7�$�q�.n)�o�'�n����^e׺+�
����F���:�pI�r��%�E5ߖ���3a_a
��̽��n�p�n0t_�uϯIAYQ�i���]zWQ k'A������]������WC=:��e ��¼�R�.�;��vy��B�yuJ���iS�R��.T��s
X۬Z�7V'�Ye�J�mArN5kΑ�)>'��3�c6F�}N�q�K��8'Eմ�����I{P���a��)�w�n��p�	���B����B�$�P�߈$Z�
֒�ZB�q�x��½BRm���CWp��v�g��l��#�}-P�2��MZ�D�)*�andV(r��<j�D���5��F^���s��42\�f�B�l��l�L^�z��xU�3Ԗ@P��z]g��>:-aW��3�-���aV
�?� ��偋?tmw4C
|i�~��
����s��P���M�ǟ�`���$-8\oi-�-R|Jw��	JTj��]@Q�l�I����4\u����$1W�m�q�^����_$鶵 ]Ƶ"!�M����ΰ�Ҙ�Ho�2-�;�	jAؐ��rf�UUTe��X��yU�D��	Ϻ�_�y*�����.�57��o	-)��?�V���������j`6�8�f��1�Q�F��l��� $`L���W���7�
���CWs��m����؛�cK��{�[�k�)���ga�lPt�	'=��i�f��� ��1m�����C_��g淁?�U�䴕=���9���_#�E��̱@���v�e=�ec�_2��##}�q�
�'(�mI����a,;�T�Ӿ�'9f����h�������h.	�hݱP��� �p@C�G�Ѹ Ǟ�e&"	?s:�bh����_:�Ff���G\�4�,�S��)��59[��D4�U��]��h*�Kr�n��TǄ���X��֤A� ��ಀ�g�@�3$�C�S=cє��43vO�j'����N�1�?oE�̉�l�4�)$	�a@Oq��i�/�
B]��U{LP&=�z.�11����=�������i�z:�|Dg��
1����V����b�����C-�K�{��zM�����E�~����v��h'���amm�e ��$S����"�;z�7F��SB�J����+���4��l�lyK�C����r��	��n�o^�M�t�C&(���� ���W1�MA��E&����h�L����;�� ���̎��=��u��Iusy Еx�%߽��� �?k��Ah�/�N��{q%F��Л)�����ÈY��*NL��c9ū�꒎��?T�6��Q�y�?N�0�7B���47������Y�̺��U.<D�?-�@�L%���5���-��X�S��ŕV�Voh43]������TO�D�Q8q
D��k�gh��K�!��0����ճ9��͹���qc ��v�f�~��fԝ�|���*�4,���+��'@PW�E٪��]_k���8lT� �����-�����`����Ԓ%���Z�%�{eTE��	�}�x�'��I�Q���?Aن�ST�2t5����v�+}��w���^d޶ҷp�q�s̎l��L]FR_�Xf�[IZ�t��#� <���:jv�~�J�� �%Qd�gU	�{���)���$�)0*��e��%,l�>P �
���G&���~�\j�u���	8�aj�������B�*�XBG:��nsZQ�ۏ�K����{=(2��wσ&:g�еKv5���`ݯ}���R
Xid�-fqJ{��I��vD�8=�m�q���{6��Oe ���5w�qC�Bȗ`Oe#o��xle��Mk������|.��������ϩQxG�伓��[�2go�������R��*z�{�� ���]Pn����=�d���u�Fp	[?Cj3K>߯<����#�n���`��τQUX�P�R�ch�����%Ě}K�
�EC�v;�Ǒϒ��~F�q�D��_��� �wcY��b���f����H��<�%V x ��A|��V@�U/�������܏�zJ�P*�|D^���W�(�Ơ|�`�Niߍ;�ʓ����LUha������X��#3�����A�e@����+�zT��n��Ϳ�5�(�M:R����ݾ�Zt5�P�5��/��}~=�-���xƂW�5ۖ�N�������f8:'�<
7�߉�'o�ߚur:=�֋�J�,b�,@/����N�_���Gr�qV��S20KmZG?�؀�['��a@N��5�h��؈U�N+K��AG?I�fɓ�B�Dv���4�x����Yh����wZ�ap�X��LbD�q��E)��JhYNw���DxLl�f�ylX�����n�{f���w��j@]3����_���X���4��ӵO��)0g<�m՚��S���m�V�M
���!�4���a_p8��yA�ԏ�[~La���*7r��r.Ĵ�؟9k�S��k��=���&vn+ۆ�Y�2�h������S������+	c��*��ͪ/6dl�r�'$� ����~Ε��#�S�எy[ċ�H�ק��S��Qn3[�b�ΩPg�w����NC^�t!�q'�"��ѝ�HOod�b�%�v���aM{�DfӀ�l|�~M ����M��\��r?�wKr8Z\ds�b1ۍ���a� :�Vh\�e�[�c�Ro�y�J�M=+�����1]P��'�v�Ԡɀh4�5F��(�5�p�KÓ�P<Z� ����!��I�0���gOx���^�;��+bQ-F$���U��.�m�4wӻ����% X+);�9����^�O�dԁP��~o�Sd,K<-y.�:�=�o�<U λ�&�-�#ʗ6���V���y-��_�As�iҗT��]��Y�JC���0
X�2[�����G�d�b�j���3�S�����fE{c�=	�$u��I�o�-L�v�tSV�����[>}�g�'˛;�J�J�0$�@����N��7������j*���+�-�3��0]�U;���7�sK���3@�����-x)rg�F�����^~��M�\� ��Μ�.
�����.�PjR$R�9��FZ���6��)��}k�lP�����Q�����S���{9���	p�L(l���7艴+��zPw���=�LN壥�����ra����^r�< Ji�s�+n��d�ų���,q*t��I�r����,o�ZX�HVǧ��'<�;��W]�)�E,P�e�����nz��{����� �#F�_�=�q�*"_?��#hn�F*�+t����%�m8�	�_Y�	i�;�ҭ"�F��q�ג��Y�7� l��L� ��·��)������1�L{$�[R�͎?��Zm��TD(yʙ	6�ts�wkE�u�߉�s�m�/����3qJ�D��Bҵɳ�����Cwʬ+�1�@
9.3�?�����\����@���Z����JL���ػz^oc�uk+��}t��.{�D��a��^U]��8;�������Gw[�I��GHUD���s�S�Vĕ�z�.\@�YK�hЮ��o�ni��6� P�S�R��L�:��+ ��_*�x�c%�:�F�T��"u���y׭�����U�Kʛ��I�?���LE(�8�2���z�Z�ە��NXEQ˧��"U�h���0ۦ2����_�O�7|�03��<����%����������(�_̮}d����0�O�-���ϞdT�O�aOr<��x�b�OB�#^	��b��Mi)D�q+�2�,�" �i�o[���NM��\���g�)s�Lw>i)�Sr3� �J����$c��qi�r��g0��.�P�G�����D�G�3��<ը���()����1��
N]�	2�h����{öS�`�&�ED?�	��1�a������ZC3/�/ǹ���'�����OQ���Mx���(�����ւ]U�@ ��H��ip��L�BNۋ����e�6�ݦ��*�qfo����jd.蜙�SyepG�/c*&�����b�R 6��x��_�5Υ�q�����@@���y,!�&9��:4���Dg=�W�Y�w�^5�H$�CZz!��,;�p�%�1�t�gR��D�Vyc�(1���G�@(���	\���w
���>`|����?��ީY��~i)��R�AF���/����KqB�L:
VVA��J9��Y�`{Eӌ�[8�Ũ���L
�b�m�[����^��O��$���}CB���8GW��XA�;/o�y��NT���3e��q��|�8	��w�p ����i9�'�~#�o����J���up�{���nɯ���b�wW8ק�?�ED$��-�J@����D0u1�@�3��;$7�w�)\=��R�8�}޿��]i��Bw�b��h���:�5�N\p}�7_DV^��˄c��܍��YP��oΝ7�j1��81;�:��l�3Eg�<��¸���L'����V�C�r�`��{tΘɨ��D���i��3��'�c!���	�1��������%U&��
��6|6�zc�.������ܲ�{]�(i%a.���74*��NR.���H�^p�32���½�H��c�����SK_;J��2P�.�-��A�%C���xX��x}l3�����k�e��S�7�NH�0[���k۽Z��O|�"^�}{��')lC��A��K&�]EA/�B-���E���/����ʌ��g��K*��7�;'��E1��vm'��!�jԵa���[��feJ2R�69��L���j�My�׿�)Q+�;�E��Y��D������G"��#���͸�o	1Ĕ���7W�����!/����<� �d��  =5�=Ѩ���7��]�$�E9�|�J�$����Q�t�� �J�V�k8�܋��K���V���UHr�a[
����Ơ��z�gjs�T6K���O���y�*Y�G�}�Y!+����G�lVT��7b�Ȟ^\�B
n��WCkG*L�M��kY��
��	b����;R�ɵ�kV�V��w���Q�c�2p�-��|.�ܳ:�~:IF:�@!Un%Mmd$u�(�uڸd�2�@<���$�Kx܃��H�A`u�Ӽ)�z�t�j���-�7�I���M�NȘB*4i��}Ij�����:p	N�;��C#���-X�N���c7bL�&���-��|�\�Gk��LP�яd�c��]Zέ,K��d���"��x�a?���@�0�J<�v���Pj�J���o���v1K8���/:���:s]s~��*7�Sr^�{����W�n#-2y�d��M�!�������}W�τۮ4���8�Z�0Ɂ�����n?��O��@�uEԟ�X��xc��^�*��| ���W��E���h���t��|�9V����y>�l����C\6V�8@��hs�����b�v��6��2ϫ��8�
����(F����f�d1�=0:qF�_PF��ջ��O�}[s�P���-�f�PA�xe��_��dHex��-F�*e!����3t��3-)RvC2����N:F�����u7d�n� V�Ӧ�u�S�Q� �^�w�9#�� $>��X|�Z��^��.+�%v	јF�w�H4/tP�jo�?�R�9"���򴡴	fS��V�����7U�!��,)�����	#J��xj��K��HY������Qe� 2��n�b�R2��D�v;e�jA�P.gE��N�ew��-�`5c0�Y�a�V۟��W�Eč ��d�R_�P���I���7���~���mu}�H$5_�-u~${������$��Ui=����|oPw�_�.;�i7TB՟~�@b�%�bk~�ӹ�y6YhnBP �2���8�9�0�D΅C��F<����O�Mj�ד@���T����g�������z7�pQMn�$�"����=���f eѢ�����T/8\f
�m������\�d���0m�d�LN/^���}�L'��_�_��>�fLHRa�kk��}�g_6��E�(C� �R�=)�a�/��L.��g�3�����hn�r�/d�_�-��h�~���	o�Y�V���P�n����Z���	��|�����,�C������X-�Q�[	�r<"t�⼅��{B�n������.]�Ԧh�r(-���+���N��o�D�P�.'��D���
�y���Τ��P�P��\N�)���|]�n)����~N���MfO=�*�[G�����5w
�Imɋ���|�����j����MQ�E/�ғ<d�o��R��0[����-����HÕI>'@��s�}��'鵪��i�@ʬ�-��6�����t��!;c�e�����t��d���.&xl�L޻4�<\H�c���Q�3>��F@q�_u,T��䞛��U�d'T~����A��'��tH<�x~2��pO�@�H���xL��H���$JШ�['�>s�#m&!�͠���kh�x���I��!��e�Y������sv�ϒw
��UWؕ�.ϳW<�����v��e�7�'$��*�`Zy�u1�a���8^XU�� ���q���(���&��˜`�&`�O�)��)���L��P1K�+��S5��%�%"�y����|�D�����LYBMͿ�-�p#�}E�jdz��`=��fz-��T╦���2{D��+��վ�s��>����]��iQf_�M�ܚ��ZRgsKe�Spj�H�
��C�E{�ɳ�ף�B���(*`늀]Ȃ_����pX���C-�@n���)tI0=� ��T;�����y<')�A����on��OǮ�+N ����E��n�.�9���1��.��Z��Ӆ���J�]��fp�-B0�<�M��9�[�'�2�fR�$�LPhT�G	 EBU�.���T}) ]���ȡF�{c9}7EXį�&m�ȍo��Ƶ6����7�':oHy�i�}M��ö]eFƯa�o��8#�["�%rx��R�1�6�O�8`:����-�܋\N$��X����W���e�;�|s�C����\}o�^�0mz��� �
�v2i�pm�A�ʈ��{���'��}�G�+�N�O�L�I�����9��6I�!���*�3�OmQ�p�'����ߩ��� ���{�fj���5����В�qJ���	(��;y1+G�ӆ�+�^�.�B�4��%Ȝ�.��0ڳ9�����k�q����8�#گ(!g&S"d�R@���Ƨ�i�L�ǷPAř&\?�d��⣴��Gg	��a���m�o�hV��M����U�_�X�x�_��	e�5��H�r(k7ެ�5�q'��wh��t�vc,^#���o*R@<�1�_/��,�բ?T�]���~q�X� t�P����	P/�-+��O#������2e�3�\�R�Jp,��N�ɕ�T��S�k��{�B�#z�'Е��QLD��yy�F�T�	���r���:3����A���j�vu��o���,����.C`C�C˝����ˮ3|v�^��������=q��6`��J��t�+Ք3�՚�����M��\�T9��ۍV{d�_6���A$���o�Ϸ
I҂eg(��.��d����.`w����+x������B{N��[H03�������.Ot��������<Zf�d�ˤ���{�����8�~Ɉ#��,^=��G���ۇ�)^P=z��P ���Υ[G-�ub�7ǚԶ!� 7�&:��5U'�di�J�R������n�^s�$�G��)�0V��؏'EպA��?�����Iα���f��Av]��,��*Ó��I����cB�}��R��3Z��\;�U/@pRg%b�~q%o@G���eQ ��(����րd�+9��s��!��������i�=7c�dm��Ή0X#U�p�`�?{R�[�*!����?�g��*�n1W� q�uU�l�8�,�V�<8a�����_\5ͻ&�"Y����L6�aT�}����V�N51���)V����o�y�z�_���h�j����Q8?䔎@�kT�&�~��6�6��9���1�5
GxC6��]��l>�%-4e+Rn�R�X��Xq�X{)M�-��ċ\�A�Ō#U�G�2�%��l��׋������;�;�|#E�5�� PC�R�޵(P6��B�;�k'�/�0� 
$[�G�����[;N�Q�����x��&s��E�(ْ�Y�m�o5ߓ�U�V����u�f�m1}��lT�UU��W�v�V�~*�K�|H"�Lי"��Mbf� �ҹ$�m��؈בduX`�n��-VP�������,s�:�#Ok�<zqh��b�������D�`�?n6_OQ�)��G�<�bۀ�6�Q�#�|�;�����������LM�����`���l�B14��>zƼ�¿�0������w-��"Q	��'l@���=��&=ǧ������K�V-pG^��Ԛ�ײd]�J�(���'�
�r�M�XfDJ�x����H@b��of>�aa��N�|�C�I��׾kf��j�b؍R{�$~��z�yo�4��Y;O�	���P�� ��-p~$�b�w�ǫjNQE������9�E�ԡ��G~���4h�2�7ײ7����:�^�A�۹��X�~r�Q��U�Q�P�� �dȘ�V�N�m���F&n�7����ϗ<��{�˥3��A�]�FiM�<��Ŵ:$��{t�_��ԉ%/������TNg�Ҥu��Q�\��"�������\�:��Z;tE�%dP�J�.�j�X��'(�}W���遙?��m+G�q;.��<�]�/���8��+X��=�˭�p�!c>�"���,��o��X 7S$[�]�sܹ�uh'�()e!�~����MC�).�f5M�~�'d�Q^i5�{�D��D>�