��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jåا{�\�u�?߷�dn@6�zf��r������;S�����*���	:���E6��(��1��V}������5�B�����+]��Hu���'s�(�����}�ؒ�*н���Z��x�z�9C��\Ԙ��&%�b4�^%��1J����F�P�a�ȕ�S6�5m�;����3�#��:�S��r��[�j�@���JUȵ|k�H�&�ǂ�,t�L��[��*�:�¿Fa���* ���fP1{*���C� ��+u��\$�ZV�.mp�jNj! �6N���p���woN+h\|��W͏�gyv������q��`^i$�\\���J!�G�K�^����}O=hr��vD�+b�7��t���%w��Z�}��t/�8M�T�j��X��n�l��܎�����2[v%�a�P�_X*��	�2�5
����|b�{<��}Ur��w9y7M�^}w[=�r�I:�f��4&�;!S%`��͟N&��m͹>n��yEai����Z>��={�] �q��6q]�(g�-]mjB9��T~��f�p�/�!Y�pU�;|���lIo�U�t�pI�����:2�jI�p,��j�������Z0ޠD�.����[A�v�U��ۏz%b+��{k:P��=)�Ja����Y��.V�c�>�[� ҈Es{k��r9���I�q�Z���pģ����P�4]���σ-!��#�{_O~��ה�sY�
��#N��G�]�Š�:�[+����Q1�=K���'iu`
M� 5[�ܠ)p����=f0�"�a_��h@
5gC�2D���Ƥ��zo�!�B��xzZ�*�]�����2=�]u�VS5�R�����SWj&b>�������$J����4������qS�S��׿ũn�m��A7/P�b�	��J�ϲL��5V�cg�[�L����	�QMA�0�f���O����;��k�	�>-��ɦ>�����ˑ�\A�a�����9ߢtg�����8����L70�֎6:�g��9�(�t�\w���xh���	��V��"V��g��c�K5S�)�;y���Z�uJ����C�>.��MH��H�+�p`�ti[�S�A��������y��
N�(���p�}�{�J�vBe��5�<�]�1@�tT� ����w���˗9���.폆P%e���: �d��K��G���?��ʨ^^p�XN:�:XJ��o�'G_?�x���o�p)����C� �?��?@h�L�]�?	T��(&gr�&��t�,������z���7t������vKt��`��~�tuƭ��m���WڐCP%�)$���+�5��i��Iн���t��W؞����G�_"�&������bŐJ= �̒��I���B`���-T2���Q�\Ӵp����B��@�ʷ����@x(�G���8�������@W/WBRa���?�H�� �|/J�n�����o�-*8��¶ǝΈa�m	?A��r�F�&, ���|�!(�X����_�*��dpM�[N�27Xkx�`�O%���]���Hy��Q�V5��T�«�M\2����t�����2�Œ��Ȝ�s.Q�QL	2Ʋ��Ş���_�%d�;��֪}��C5U>uՕ�Ԕ�]��9kH�N��`�@'����|�������Y#����?}cg��oC�U3�����P��$M���Gݚ���X5je1���c����]�7��l2��~���~�Z��|�,;�$:�+9���<ZO���\�^�kn�:�i�c�	�Ǥ�]��Bk{Җi`܆�%�&���c��:S=!hڪPQ"�{%�/Ƈ��eW}�LL�.��0/_�"Yr 0�Xu���<1�그P��*GN|��1Kw�ӆiN����C�Hu ���J��Ҟ���$�+?��SLp1l
�R��=���2��aݳ1�l�#,-ν7�(����Jn6��L�6*	DB҈��\\��|�<V��d�0ԢR�_6SX�d��	�������l�닑��ZOY��Z�H!Iiˊ��}� Iȼa�Zc\�Q[��k_�C�g�6�9_z�x��	1�b���"����q'���Dy���Y�/$&�;�/eLV�Ӹ��k;Od��MXYz}�g+۲��Y����#`���n��V���ܯ*�-6x��C��K�$�sO�.`�Y��X}
����W@W*�|���a��R�
i�� v�O���I��J��"�k�c^������CSW݀C�-0y�J�F����1=ݚ@�:���"�y�`>p����V��ÑŦ$hG��n�|#;B���"!Z���y��ҡ�a�d�:�I�ǿ(o}YFiX��E�)やz5]2���^�5%v�h5�¢T �'sP^t6�S�:��*l=|zm��(�!�ٯ9f,:��1l��h�pSDa�@_Em��.��ɰt_��c沣�|֚P���>Qf�׋�����*�e�ҤcSG@���̌����~��)Z����Δ�ش'�O���3�[�p3h�{�ߛ�/i]JCmD"����ţW 2��l�m��/��ݘ��3<�*Q�.�<��]��(A�wκY���
@�n���~!�� �]��*�>O������ P�����\Q�ּ۫~C�.d�wm��I�K����m2�P���������؏/��UO�����{	A� �`��G|g�k�̹����"���XP}��f�81��g��f�tIi+B�u��M�f�]:�
�f`D<���!��^���P��qYߜuV���*�`e�Ѕ2�FH�r,,��6pG����:������E��a�U��x`�3f��#�����p�Q���{��{��v"Ȇz�ԙ�Uş*���1���e+�a�#��u�ֻ$�Dƺ���0�ݷ���L�t_P>���x�>��:!��*22�
����~J�b8e;�aU�`����!N�k�/BJK[�	�����ӽ�]dl,�hYP����7F(C~@�>"��h��<���'�1�fV��l�X�	���o�X�Z��_�I�����s��>���g����W�h�򇔵U9Naz��~\r�t�(��u�[H��̰0㥇j�j�#����X
~q6ƌ��6^�u*�wr;A�t��P������	�kdLq�Nl��m������ᤥkU�r�O�x�2(���Ч�&Q�Y���������Mz�B2�P&�<,�YJ�����(C�<�����N�� g��k�ք)B���2<R��)��� ䷠�
��F7m?�+�������8M1�����D���s�k��=�A��=���;Z�!���E�[ߕc
�vNrc/5D�?}�6��M���E�<I���:&#H�{�ռ�3��bɶA��rvK�{S�Q������z�FY5�c¢�YZ�K:�|���kq��kR%f��7��]� yq���� ��F�冩m��kx����tΪVz�x�A�t�O���lOd�v(�6�\L����q�
S3
��g]���g%u����͵AYf��	N�ԓ����)s�-gY�D^�3����o�Xr�����C�������(韵���Z]?e��&��`	$����s,1�u�]�T�v�r�1KE��j2�������r�G���e������5{Q�fi�������c�_3T_p�[
4vؘ��0Ć�����G��}n}��F6���%�,�.�����3�ʸ� W>�p���t�$	�����GG)O;����٩[�I����q�3��z^Ό8�b�{U��OpF��xu�D� ���E;Y�ŪPb (ߕ�>���W\�@&�i������A-�/xV{["ϖ������ {��fZ�nc�53��f�,1A ���"[~��?]%Ѥ�.�\O+&��'7���d�{#h(�]_k�ީ�'��sc4����uj{����7 S���M��]���zX��w���x���I|1��V�u�1y�09�Wn8激B^B�Ұ:��\�?$K%���-�r�b��k�"����eөC`�$��#�A���N��2eb5�W�����Ddh�3�q��O0K���)�B��R����}�Ì�0�<z�8�L��Ę���ԭ����Ǖ�+I�(_��3Orݯ�q^��)�7�

֣�8C���*]�aZ��r�)����Dԋ�Ȁ5U�;�G��H�2}.р�$w� �9u�Ŭm�)tD�R8ɾ������B7빪[���q���g�&Jw�]�p?