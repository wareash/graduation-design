��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jåا{�\�u�?߷�dn@6�zf��r������;��1��B�	m�)�OE_dx%�~�,�Xa����x��
S��Z��S��7ԧ��� l��i[�:���b������ ��U6ݘ��lM16�u����;o�35�8��Z
e;`�߁�E��s�|��0�����_��Uh+�XF]�YmP�ҕ��������h���a�������W�N3�sIu�� ��tz"/+�;J�t�5C�{	�S�H9dXL
T]M���FI���F�E\)]U�Ǔl�)����u����)OP�9�*�z�m[�J;�d�<!_�
)��5Z����h�0���~�����CQpc��Q����W��ئ��V�9hϵ�U5�ת��	��i�q��d�"��0|�Z����ȏ����<�%l��Z��,YJ�p/�T�׆ �y�ȹ���nb}*l�qy���ߓ�1��E�L������*����bg>�s���E��pWVL�@��� }8�n(����� ��o�-��\X{`�:�U�H�d�[l�3O^�Q�m02������׋h�=�OC'���	i�6�JT��Tv�Qn�T�#+jL�%�p�⤍=�[����r��� �4"j��h������
;s,l������_^{+^�h���NBF�Qf�+#\ܣx��!B tt�q�4� =g�*<m��38�ق��d��p�LrUw���l0�֚���ɹ�P�V,����G� �1�r�92�%,�(c�S��V��1䔹�%�Y��{D��^�å�v�O�4�}�r>�2'7Y�P�� W��A��F�"q��%oۭ����ӯ�9l�	�0/��J2�o���b��cE NS��'��y�8R!�n�X,Bfڮ�`�^�|��r[�;�)���*��=��k�:�*�g~</�ϯ�L�Pi��,]!ɳ	!%�W=�Ν��Z?�ſ_lvac�`��G� ·�=�LY ���H�s�3�Hτ�(1�Ư�u�Ǔh6_!YB\ѣ��1NI�whRG~��1���nu�J^-ai�|��\��{5�F�֙����(�W��h&�i�K}�<�	9:����K��A^Wx-w�jVeu�ԇßF�[5��S�qt��P����z%Ǫ��C�ǁgS�]�K!��ri�A6�{��MR����(����
ݔ���Wv���=��
�(r̲��6�v$	b���0������P
�Nv��e,P3$2[ɳ�X�x��֕9�	c@��t="��>yD�������R�{�1ܭ��B���`��i�!�{�N� �?}7`�+���W�l~<�Q�!
��>����B2+O�������f/urz.M�և�����X�� ���p|" �Z��s����U����g��pLdZz�BZZIZ�ӂt���[��G��h�Ă%k��n�dڎc6V4���w����?Z�D�߻���@�D.�(�j]��9�<k�=��,�w�HXL����gAm�yK��F�#�ȼ�W�=�?�1!��@���8�;���{���}s���~ZЛ&:���(0t�^��c3�����[���ǰX&1��r&h�@@t�	l]_tM꼺utϠ��"�S?�����^��[�WJ1x�
�fU�AD8�`6KԶC�/�^�$����m��Z�{�����8Z��8����o���;J=3��o�,�3ӮI��"��	���PZ�p��}}��G�W��*��SV����C��b[EL�cR��i��E�y�;�8)�"C�HEG� ����� >��9_��6Ty���������!�]Σ��`�!I�{�g�6>�JN�����D�!�K��[EZ��n�N
 R�����i��؉p�"�����D���'�%��kC�!�2�P�2n#�N}�R�.kc�Md%���{�A��c/�T]2لX����2��=��:dt $bg5��UZb��+�ϴ�C�с��@�����Z6�Ћ^�"���m���)�s-�7�N��ʄ�&0�#�!_)�`~�"��}�ӌsb�ʔ�W���:H�	�ʦ(���j]
:P{�*4��]��y8���r�M�w�`�fϯ����Vm-%�t��\
�0
g&��C�����rג��ѧe��j�����r3h_��%��P�(����W:m�qh���B ǠIu�[g�(V��r���
��!��
C'�I�Fۙ���h>���%�ٌ��n~�3�oi�%����*�Q��nѢߧq�F�ԟx� �������<7*�ȇ����&Y��k�1��^.g��E�f.��%��_��v�W���y�h��C#���v�rc��nv�V-Y.
�m������`g�_�,������*��G���W/V�	~�x���.��mh��> ��"L�B�������t��ι����A�>9��Bُܾ6x,*�����	ݦ
�/wE֮��$T���@t0���Z�F�wEu�+��/n��[��_l���n���Q���OqC����I�D��vq���]�5�Y�R��g0+�k}3�����?�3���ю�ē�ػ�>�o��T���q�1����D����r�׭/��:�K}�G�=a�/��G8�j��F���3T�mWv���G�'�6D�ǽ΀�'����&���3�b���j�t��pQ�
L��a�dz7I�A�/;0��kp!����[S9�|�p����Ȃ���
]����'��Jm�e(�RaeA��,�ADF]��i ��)̹��bh�fS¾�\X�y��bݠ��u�Lm��~�L���\�%�8a��*;y>����X2����-��+G�G3݊�p�}g��`꼹y��.��h��~/f���}	Wviy�lG=��=� �]!~�'�!̴�JcLZ�R5]'�`7��@��/��Ĵ��(�w��s�|�x�v�V��UY,�|$�w�.���fd�O{��;��ևL?�4���"�Ѓ��6�FO�CM֘���d�2����ꎽ�.�ҵ>¤����)(���+���Y	G#�G�~�������� ��o�g�}V��-�o���fŖ����I])I�vͮ�d-t3������g��ߩ��vC��3|NM�l�$I1/���8����{jkX�J��|�6��e�5݊��rc�3�NE��^U^1k#(��b�}��ħ�d�-��`rWtX'�߳3������0 �Oʙ��SM��1n���
!V�t��g�Պ�ERG��`&L�u7��(#�L�������A%N��a��߫�0
o���W�"Ov��OY-\EY4�	+�4;G/;y�Wj_�X"ϛ���ߊ�W�Nv��8�l1Wy,6(�G�3��~��"��#o��`�P"xT5n�$]uI���04h�c��e|w�0v9q6o��0D����q����k�:��S=hH���&6~��oI�Vh#	�%ر�In��c��Uۛ�G�����A7b�x	g��Vr��"{k��E����ăI����-������6�����нH����?�o�#m�2�=�C��7���4
�ncH�{u�M�<CE�&;�����:��ئ�\��7��j�M�ק��Ϫ�k�|�f����#
� ����+��6g#s���;0}�#1D㓉g�/Ya/J�UQC�.�l��i��g6�qAޘ?!r]@HT�_9R:�=�&�![V����	�}������n���Q���E���S�����9U�l�:)%I���J.���F��q`��i�>�C�K��3w)t
�Z��|u�*��������ͯ�I��(�q��n����m�-��vYT�Y�%�{}�y�=2޸PxER�M�����C̐L�:[�ʸ��>�%R!��G�(�$ `� қM�o�ĝ��-*fYa�d�9 ���5( ��q�-�6�tl���n����l�M8un�r����F���}]o-/�4����l*P��wS�xJW���oW�ge��̟'#��㐸�b�#�j廡rEߛ�.�b���@���9�WÆ��E[m30�h�\zG���N���j��⅘�q�w��Y��Q��f=c��
��R5����U?��^��� Y]@a��Tԕ��v����%�	�����}0���fu�&�68���Ţ>o��=�i[>��N)Ui�	�������@�Z����ih��axJ������R
��".����³��W}����7��b8�K��rmG��C��с�%���Ղ�2��X|U�"����>J|�I����nv�}��Ƴ��'IE�(�8�N��V"��f�]N(0k���8��T�;�)����?�d���P3�r���mY�=�������
�ٽ�-?�.Ҕ�W6q���BC�i#�^'���A��ʣjEތ"�j�Ƚ Ȫ�ʹH@�tPeY�)�(��հ1�������%\a}f�|�!�2�wx.�^Y7V"0/��
��.*M�`>�a��s �0���2Mba�=�� h�v!�oQ�"��E%S��:���s;��{3�n D�I�)D����P��:М�0j���[@Nf�W���uL�UUJ�L.{�!� j���X^.āN+p�P%-�X�N��3�{����a�,�k��O(W�VM��e�)I,�2����,�<ꠂ4=�U�T_K�=�?����'�]<$�!�=�,h�G�X�o�0�u;��~ & ���\����q���CX����Z��|��
���ʜ��)�:$�i�x�����V#w��d���Q��-�����{�5}������2��{�g����W�}�&~��?��B��R�	�fz(�C�q��e\R�D����a�Ս���9�s��/j��	T&L�3)w['O5/�$\L650J���*���D��\�WȺ�Lac�N^��[@���?��/�Z|��(�l�[��{C���)YM����1?6��97���`�K�\ hR�:�����''������j^���������e"�Z�L�"�����~��Bh��r.���T�zU�o�BMB�4����gI��}�v����і�pˬBy�>J�U��[���R��J}��3˞��!�H�6s3gor��`"d�+6��p��)��*���C3�;�ŧ$M Ml��c���%>���yG�(�h�-+��YJZ�C�g��8J�tF(d�	onxma��ڄ�����o���T+�m�����%?V�4���x<�Ȣ:�S�x�9�PT���
E��p'(��72��0-�n���"�ǒ�r۰������K�9��W�#�Q4Iɲ�k�Ӗb���[�>?Vx:�v�Jׅ#0G���?�3���$�{`��
�ME���d!�y��:��`��uT�h��F�ý��w�'\���h�������l4K��	1�\|f�����w?lsJͲ���
��D���X:��7s�.����
��?O�I�b[�{���ҹ.Y�/CNV�+�ǞA�,����9�)�%_i*�!`�KX�:p��׶r������e�M��6 ��Z�������f�hbBĴ�W����*����`|�M\�фn3��VsU���=,����6J��!+gR� U��d��9���A���I��g�:A�?��B�㴍�Pv7��4�>�ŀ��Q�?Dq�]0Ng ��D
�e�hH&(��\L�Fg'd?n ���Ru=M>��>.p~�"�%�~���m�GZ��c0�⨿�X��,^{|V1�V�4��y��CŰ���4)��=#�����#h����u%w�j�h�//l��8�00�u�S�+Jg�P܈)��F`������Uܸ���L�Y����k����7%�����afe��@4��rL>��qF������I��r5�E*W� �7�kXS�������7Ք��{m@����n�}�5D��6���?����M`��u���hvM)b2�g�?X��A��nYc��#62�e�D�z��d���7��;�B|���fT�V�O�MN�.�%18"d���v��u8Z�Qj�"���K���ڄ}�s��Z�%�CkK��#Tܷ�#m���an�T�?{����WA2��YPb�x��{sGB�Ҽ-HQr���oS��k+�y_w���,�aֻ�T0��n1T<�L �p��7��ۃ�(��U/�9m�cH�>�
G�EM�^���+[�z��U =邟ˋ�#�p�U���^0��㋉��Ћ�F����=~ji�ၨ�1��i��U3'=�H�ɲ��.9]E�����*}��K�4�Q����l#�^��!��\��x���k��w߮�Y��{`��C�v��pd���;�B7tf��+��Ѧ����Myf��_s�!6��#�� ~�}�:��\\r�˗z���p��R�`�RO�X�2F�s���W�
P�P�l���ߨ��A ��D�e��⤀���N�k�ӫP�C��sV��D5����ܾ����KW�H�Ɏ�a���Z�KS����:���OWիo ��:�9�0���_��쒨�?	޹M��@�^�㆗���y��4�{�`0D�}�*�6 u ;����1���J���2>�P��#O�S!�����km�S���O_�Ƚ�`��r�tk��Y�ѻ�êfQG��R>�r;_�n�[V�㖶Y�_��{�y)n��둊��_M�(�հʩ�١�R�
D��rႰ���Z�@���U���LRB���£-��wk" �r�۳���ȊG�3��[4(%%�v���"��y"$d���2�I�ס�"�,=��R3�a{��2�{��qF#�^���<
C�R����|
���8�%b�o��>�4�Q�I3�+�G�A:���7&�A�|.��+(pz�b�N��(����l�*Ut�)� z�%Y�Ga;�*��H0�M��o����-�����騮,d
��m�e6K�)mB� L��X4X���0�4l@q�*�~�C����Uj�`�,P2�K^%vY��a<�a7�l���1�Ϸ+��gN���M�6���|�;!(�޷���G(mŇ�S?�t����+�+E�{�Q�9���0�@u`�j2����W�պ��kܾ�i�{nb�:������,���4�g��w��Hz@��t���e���[�� 4CJ������tu�� 6�m~��(J���Գ]5L�n�q��:���
6���FpÝȠ�Dz��
�Kc/�L�Ε��Ą~�T�=�U�I�rEAfR��۠z��7�g��6ߙ)�����_ �����6��c�~��� ��I�S|���t�4�B���1�E��d�'09�������p�j+{�.�Z�(���c��H^���T����.h��j-M�>��~���b��v�,�{e�#�32�I�$�u;gK5'�,ߥ954)^Tş�G�#?B�R�������D}�N�����28����� ��;`�_Z
�؊�h���;����oq(��%\�<P׼��5g���{.��9yk9�/������L{��"/J�)ǁ(*c��=��M���p?M�#z��띫H�.�Q�4�6%�)O��=1����Zl�G�WA)�rj��q�\�lKux2�ƲV73���H�<�l�:3|��?+�8�s2BB3��T3�~�L�D���J_����4��k
}|�dt`���m�p�ik�����y�n~9aqʺ�p�ԋ�����E�l�.Nf�b���f9	���|�Y׮Ϡ?�l�ǔ;�sЛ�b����1K/�����E���P�Bt�t;��}���Wԛ��?Xd�/���c}�&�A��&� 61z�������
s��װ2e�u/�j������33Kz"�$kJ�T�n�ƈ��"���|5����y��6Hr�m��8'_�Y��v�\E���	H����G��љ����q
D0c��-�]|:ӑRe���c�Ǚn�7�*a����N0�%l�A1������li�eFp��� u�im��^Q ���eJ������h�R7�Kqg�9��˳���6���b?��W�ʿ��R)C��1i�� 6zҀ�Iñ�h�0k�N@W~�z�K���%(!c&���Y����B�¹��<Q�2�nB�w�^��99>���r��B��	G��O���Ǹ`D�ކԞ���������=��+ ��"lqN�UP�f�K��TX��`����	�E	eO�N�?W'�^-��=����}��{#W�,��k�gN�[ڒ|�#�d�у�Dn��rJ�cq�=KN�kq�lM`4Ŕ֌=	�ǡ��8�.C5�ʫ�v��Ynޣ����XRT�R��ו0K�7x t���������]�r�g�~-�]�Ӽ[�yj�!=X<��I�x2�hsmn$(�/!�ݵ ��=���ّUB�| �+��"��[/��q�3�g�Pe�WI�ℇ��c?Gn�L����P��jd�xT�ː2�*F&U�_P���U�'\��sX-l��N[��׶}$�	�P]��#�5���t�`�6B��hV\1>�u04�U�Rb|�5�劂>�N>c�l��Fo����=��(!q���ŉ�Z�� H��#�ʸ�4�����	�汲z3O�~[�-�Q����3�=m=�ړ%��"�7��W$
�j���wc|5��G�,�ɮ��`;����N�[ݵߖ
��X
Lˀ�.L�-��e���I$�u����q�5M9c�Re&��������^S�K~F�᪥3�T����ڕF"Vy/������C�����ۭ�����i�j�'��U���t�tb������T����0P"{��CY
 ����Y�[t�D��u�y���t(��r+�^)��I