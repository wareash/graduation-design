��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jåا{�\�u�?߷�dn@6�zf��r������;^��
pt�h�s�JH�iK���R*�e��MN4�w5X��2k���E����&bA�u��\D˕yV�nP����ѿ�'��+dj*��H�v�g�-gD��/�P�fz��'�|�VP���~E-��@��&ou,�����`K��#:F�\o`��]q�2~K*Cj�j��78�f��LW�<'P! ���=+�F5�Ǉ�N�Z�`���bщ�5�q���W�A;,��v�����Y���#Aq-{5^�o��G��i؏����_��Q��{����רN��b����7��d:�	C��91t�I�68q͠�����Z6~���-���oA�_;W*T���hV��9��9����$(�I�M�ڈ�\�T��0f#�3K ��E?A�R��n�|��J�z��S�@�eO����HZ3lN��)�l
�����R��'O��@�P0�L�N+���k���H	|�{fr7��(�L�+Iܡ)�_:������oe��;7%V�Ha�ה�:�T��3� рf�`Ҷd0�,Z�I*��'u�	�@ͫ���mM���>��
�RONM@v2�x_g0�e�OL�ÿ�<<R*�w��!<6?�]q5�� U[�A��fW<\hN�J�+������h�>�\���g���m���J�"��2�'�T�4j$�GKzYpd3���'p���MA&��P�=��JX��`]�����NF�{��?C{4���w�d�Y�(K�C�
�);��g����(�Tq)��`I+�]�^� �a�ٖ�,�_��1�x��ph��#�d���l���,F�$	lu�	��	�h�RQ��O�b��6ȉ�;�?+�}(���<�!�>ܳuVo����L�j��dT�Q{0��~��V4���	 	������6'����سO��GN��h���6{�D�m�u�F����1�����|v=	��8�*�d z�����������-	yM�yE5������\|����ÔVՄٽ�Z'���H��C�مr���D��������,sԂKIQ�FuKָ��������J����J��F��p�jW��C^�����)�=ƛ����@e��n�
fMH����?[$z L��21���.���Mރ�*�O�;"������E�X��`�!@)�Wg��߻ˀׅq�e�����5��ϋ�_��/i����ohߨ�	ZM�g�^E���>�n�t�
��� �]P���DK�l�u�o,#!+�0����e�~�P���P~����y}���D$y�Un�Tu@]�^�[y����@��r&�LCf-�o0�D\�q�"3'=�U,G��E��<v��2�]_a�E��&��5��=��$Z��bO�7�-i�;�Cx%x�X��ң������u0Z�k��*�E���V�S�@����>9���_�B~��y�5�Z��]<�$�o/TB4R�+8�� :��.�5�;��y��l��0�\	c�D�tܛ�a��Fp�ݗ&+⫰#/��.d�$g�\o����o��S�BԈ�D��t���'>TJGJ����n�|�wM�(n%Yn��iF5]�(�l��G����2C��ϣ�@��_�e���=�����8V�T���/�.b��A,=�|��F"���K�L����_�_U�0O{�A�i	��Iӏ�х���O@+�T� H)ۨ���!����GA�'l� �9�Y��w�����.���� �d`:�6�TQ`��l���>`����V"A,���0!��g^��a�r!��]���ks��}V5���$�齮[���_!����lmd��������A���(q/�}ۿ�bW�7'H�˨�B��@H�,Q2�����>���ئ���0�2�V-�T�Ew��\?U܁ҥ�6��~�i������g�J�
����O�@�'_�"�ho�45W����0w�B�6G�m�ֈ;�4}�q?�t�gt���&h��O�f��Ҙ��8����*��@��� ��2%V:؇�'y�Y�x�#�����Ud��i ��i7���ۀ��
� -�c؀R��Y�
���%�7f��>�9jX���c��ԕ�mG�X/, ��Z�m5�Eiu���ό݌p� �[-:�3�G�^L��d�»IM7k���RJa�3����2ޢ�?5
|6�������d�Z�d�S��p7d�X �w2�)�/Mrg����:sbPێ<�q}[	��d�H�ijV��w���<:'�x��i����w��F2OՆ��w�'���P.=A���ɐ����Zw|�ݞ�]j|������O�#�%����*���X��Y�.`0�,�?�4��@9C$I�exh;4���7�>�,��0ANwGmo{(�V=W�ݙ�ȭ��wtW��ߓ6�U���u,�gϊ�5�_x��A�D>=��JO�]�p��T��&��Eㄼ7�j��5��y����m�f���0Mg��mQP%�`�T�d�뼚��Z�\d%�j9}�W�L����2�H����]�>�'��,%���̂�ߛ�7?�����)L
�}�a#F�{?���K�S6߼;!��b�G��)4/�|f%s?���Pb�r@J�Fl%��D�h03��d��p�v�!$G]�/������O�F�<�����N�[n�y�%	a�"��b������5		*@Bo7��*�B*nQ��'W���}��8#�;�K8���l����.���b��}*l޾
r��d��Y<�q��8:�)�*S)ЭTP��S8������o@�*�6�i���)b/3����eH!	Q��E�_��0'0O	*��2����l����9n}>
�n�DV���*�M�º�bb?�߾�?s|���S�Հ���+�=F'�4K��>���A�H��N%�<��+��8������e����a�,��K&r�z/Et��=W� }C%�q��	��ӋpAf�ɰ9��/��d���8n-�xB��)z�*���k�$���r��`qJ� Mȍ��z��B������ �a�i�J���J��8G���$��H�Q�ZR"�h�w�c���䔶���UpX����k7E$�ex�u�J0�B��^z�\"X�{<:ֳ���a���w+��X�Ӑ#ϋp�R�#~��T�R�T��/�}����e�Tg