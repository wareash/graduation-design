��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�k�۸�m�i(b[�{�㇌�]�i�5'�`;Etg
<������H�W޵α���N-�`��6����ݾ�FF��eF4��_}<�ےA�[,�|{�?r+-��ע9�!�"��F�Wnb� �i��a��c��v�Ϗo@��Z2�[�Sh�+����,��ơ� �����Δg�Ф�vmۗ��!��Nt���Oa�Z]{a��x��8��O�uE7��P꯫��
���6֚7+�b�&Tٰ����B�D��=��O�z��o�Ӱ��Ŧ;[K��jl�o�%H�4��zh���=��-D�Bɼ���u�%hCK�#K��|+��$��f����[S��	Q�#��d���<d��P� D֖gM�)��<
���.�4��I�q̗�o}	`E�y� �=��Ȋr�gz�3�/�T�B[A�1�E������5�sn��+s�n~�������Y��)�p-e���Y�#V̞�!HO�	'��E2��^�|�e��5��&�f��j�ݶ.Æ��BC�᫞00.����͆���Э��5�I���N�#w����h�������u�z��z��R��>s4(@��v��n-����������	�����+�r,�bۮ��b�y8"��I�sS�mMZS|�W/���i	v��5�N]?%�.��|��Z;DOHS|(L4rQ��9�J��S��S'X(�0�!����F�MYR�}������-r��䷠M����Z�Ϭ��m�^b|�ߘ�^}Q��X�Jj=��k��l��5�	�YQ���y��kj)��EDz�)х�5`~~��y��)h!~�m��آ��ӔU`���*�,�ؔ`�*r�]kBH�	������@y/�nW{Nרn�|��Zh��ߙ8 w`������@8���]&s�@ݯ�S�qa����r�X{e4�kK��dZ$������.���q�Vb�npRЋ�B;,BȐ��2@<��_��5R�7=��d�l�-�xp!���=��������b�1}�ĭ(8i��y;K��(�hf�Ϥb�QYA�#��!�:+���U�"��|���R�:XM�Z�y�O��y���H��I�ິ+շ�+�2�#g���J�H��D�����,R�U�n�Z�&+'���l��NX�5r�v�����8����/�DN��oV�'2I��g}�]�H;HS���_��iO��#WF�
T+bd�����v�{�8s���Mz�����W�ȈN�M�FY��t s��*Hĩ��Lg3�fj%:e~�A{�֎xK�4���Z�){�ẽ�f�"��~yz"w��o# {�InVL�FS8,o����ξ�����l�܎<���֕���Quf9
6	��C�����7@6��vn�4N�����U+yP7�'hN13�y�ftB�4����Gƣ���W�z�=��2B�,2�P���z�z6!]_�U�y�]e�lN�+5B���B��*���>=�#����L�{>l.�>A�G�/p�kj�7��P\�W����s{�y��tbkY|1���g��r/�sL�������!��Q�u�����#]��zCbwu��Q8'��,��A���$U�O�ֲwh���
)��C��.so75�8���w����I����G�Yh�h�6�FSZ���d󛒷�@.g��i���~�@Ƶ����������s����՜r	r^>��M�T�0��]qc!����ӌ�X��?�V���|��mf�o�Q��*&����M��P���=]�1�*�ż����<,]���<ψX5��y�ԩ�R҈ݑ#/%牐��{��`�^&�ۍ���aP���g VwS��/TI��X��D�_8�=�m�j�wR}�/R����,�&��������
+���9�M�M����b�Ze2��5%:'��#$���U�-R��<Ŏ,a���~nkj��[變NV�I�p|���Z_Թ�~�Lv?:�o�eAF��欁��0�4��[�(ae4����_l��u��=����rHoZ����1U����y!I//�Bg)�j���$F�O�]m��E���Z�߄O#��q�t��i�����{(,�,�m��4K��fw�L_Y�u� �d�e�	��@V�ay!��I����K�ۺY(j3ZL����2��Ǭ)��.��x����xi��uy�I��|۳��M(����Q�G�
+�8UP8��,I�X[@{F.�ł��r�;�ـ(�\�3��gS��>M	'C$m >O
�#a�Ë@h9^����s�cTt����m���n-X��7ˀ�| ��	e�-l��FTl�B3������ ����n�T�)r���M:�r���N����9��t��A;M��{��>z����QS�-#Ğ�tc	�s7r�k"�n$�'�}�!Tpv`���#�g�"
.Qs�6(�M�sk�.J���=�t���� "3�f�xg�A��Jrj�ڙ9_�h����|�kVn#��?�_�ǱW<�:9�+s��M�Y�X��u=��zr�)���Qp����6�e�n�L��۶g�F�;-�
�;��Ke�m�k���А6r-X��b�:��N;e��I��X�^ݻt���)ܢ�����L\��D-$=�m��˵u��l���*z�Oa��.��L�����Q�Zb�>�|to�M;0��B[����wM��s�ņ@��on{&���1Ej-.L��4�����V�j?h���7C�ut�rT������oi��3'"��.�z7�HI�.�)��V���g�#/ꯊEĺڨ7x"��&N^����m�� �{K*���l�nv�Qp�8zUz\�+�_JL�����n��D�����}�6TPE�������/�=E�ά�(���!�s�נ��D8@���r���n����K^���
���	�7�T��=�[1�04ˆZ� ��߈�)��Y����Y���mQV�Ɵkɺj��ұ�b.\`@��g^EG#��G�m����V�����$�7�Ր^a����RS�7�8�F��5���VD�����j{��Q���+��v����HۚR�W#�ཬ�TX���N��6��ػ�����"�G�r��>Y�-W��oF�f`UA��}N�;"$l��QI\�j��>����\#й)�4_VA\i=ֈ��I����*���K��˜]��E���z�^����M��"(����gDxI�%,���� �A���Ms*���P6.�C�����`>�{�&]|�Ci"cz$#�kqgɅaw�L�ߊ�$��;�Sx�fQ�h��zy����o��Z���#����3���`�>���:m��f�2����Kc�h#�y �~i�q��A�U/(���.��,�tV�(O�.EOm5�?���E%f�+H��A�݇�&�����'o�HjElԠ�H�P��c��s���p���;v� �Q���<�cO-��_��h.+GX��%�@�)���NQ�d��������4*�O�X_k���ђƬ?��7u��a�t�ai>��#͘jgF�ˋM4��=�S"���?!35Yv.�H5E�ry��\�ب9ʔ���!FU��C�UY�r����ӕ��_�>��9d䫁42���Py=3��I�%�L����'�%�TpG�:����|��B�����Uv	����a�m�,���Jx�SK��(���v(M�/��4��'��E�܁.��{#Z���)8�%�2 e��(�6%���#���IP	�5��#�V�eV�-�ڎ�������&)��H�fH,���R��<�`��5�P��кq���_ݎ4;����u|ߟG�+��L��F�KE��W	�����"��f���)s,�*#�� :����jv�F0�[6s����\ ���܋��ג��~_�0q�d1QA[>���j�lJpw/��_�oߕ�7��4���!O�UM{~~^�ƞf5	W�r�����dM���ޠ�w`�mN���y5 �݊��ҽw'p��k~-��{�?��P��sr5���nӆ^�Nx��w|���9�A�U��leM��TQe^؛-��.X�!�����,5�������B=��'M;/��m 0�r��h�<�