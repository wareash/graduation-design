��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|̪��q[�d��h�xM�+z�D�._�9�e��M��g��WE�ώ���Ck��E?~��z�����^'΂��dH����S�6�%�.�Rb� H�'*@J&P����v�w��u]l��{�t�8����mԘZ'��B��N��ݶ �Y�H`#ǙAl������}B7����J�pn#oJ5P�0�g��IϮ�e���'��#�?�xO��|�B}Z��\��z
���܋��Zo�!SZ�Xg.�΋���R¿>�B[mH�M��Ü؎��03�K����Y)�}Y���Pd-6���M����.@�ͲQ;Ȇ�M��� ��^��8���dj���q�]�QK�[�;r�k����
z�����`��2��iW���.C?�}}��H��dy�T@~˔���bhw�����[�U\$W#%q���c̟s.�xp�$�Vy�� 8�M�΃�`1�4'߂�k���n�=�ԍT#��4��Ɩ՗ #�ߣ��Lg�"� $YAۓ��Gx�&��������K�rr��C�af��<�>s�>�y�#�(SQ,��eT�>\�>�\�Dv�/HxR;��P�+�
}�I�/۷ �2���GtR�6E ���p��L?j	3`A&X:s��>z
)��$��ym�ģP�R��J��Ӷa1(�,��5��\G8i�x8�!��@��$��������a_\�z+T䒧)�R��9� �Q�pxgS $��4'�j.a�6t��)ױƨ�W͢.�v0�ō�>�Ii@��
5�����+�ÿ]�"4� ��� ��:a�h��v�����������?D���Z�i��k���1�:��`�g�9���ң��w�ɸ�i�[�s��k��ka��LtE��1Z3W�
f�Ƙ�5�j��z� ^���h���=[{M$R�P��a�1^�>�b�V�F����^o"���nH�m0��c/�� ��c������e�k�X��?�HErJ��(T��h��Вյwʠ��L�
��#�p�'�P85�:�}&�:sQ2��\��+Y^T"����ɇK�	��gH7dԊ�A�D�2���`�=Ŭ�#nX/C@�"s�ZU
��	c��-��bNN�- S�XZ��\��� ���8"Gt����ķ�M@>�%I�A��2���+�8)ȎR�}-��ыVg��=	�<h'w�gp��m~7��s�ړ�+��D���цV��Ϝ⁮{�O垎'nu6�2�p����2+���,ݙ�1;L�L����U�����|(Ǟ�,w� +���4�X����.T����G��:�q%#��P��V}�){�Јw�=;�^U�F<�Z6�)�LO�	i�v��w� ��%�D_�Zo]�´5d�����4�vg	�>�!'sM%�P��ݵ(���Q ���B���
��#q�<�ڡ����K�%����叅�֢�]�AE!���7����;S���3�ބ�d�@!�aGb�,�x���ćdb�f�s�D}2�L�����T�է��&���v����r��S*�q��V���5QD���*l/,"s\�7>��s�skc�{�zXVO)�#g�[H	!P �I��Sܕ���*��d�Y�KJ��.G8QO5���y�VGy�u���h!y���G��ϼ��N�H�4��R7�m�,�O����$R�0�*�/�:�=S�R/u�D����~5��\#��QV*`���qY�2w�E^�>��zy\�ng ���9�KJM��ף3p$>��̭����`Y3]���.n���#�(����(ۄ��z�݃ff�ha�8�	��N�˛�&Z"!bCD���cF):l�]�G�8���a��������Z6��P�`ij\[�/�k��z��ZД�S���j��:�}^'�H)�/���a���k��)$��4�0������Y�&��ʄ룬�>���hG��Xa�
ys-�Pxٷ���윸C�[��+���������Yڷ{��!�a���
&)ڲc}�%)����`W �@!��1m_��	��Ҽ�=�����X�xR�ܷ���Tёp��1M1V����h6�VcI6�T���yT�+��H��Q.�?b_$�dǦmv����$Oz+���D�%S�Ƶ���w�Ғr����{�T�ϩ���#x�//ذ���
�R�1#�˩9���h��M�S�p��i���"���|od�H ��Y���"�V���������k��1�����X4��	p���Mk�I{�ä����k��qTEN���Q|��"A2��n~��JV�q�vT��E�� ��D&�o6��O��!�F?^|(Tu#�*��H�y.f`>}��G� V�m;��4��|���3��KeV`M�F����*�ܡ��hDV�t�MW�}	����g��d+<�|^�6:��W9��xD���Z���oL$���#���L�8��ΚX)z�3�
��Xs����Ju˥�9j����.*�e-��V����E\�dxMjcP{b����D2(��0s3�o�~�SJb�1{A��)M��\ua�5�	9�Ua�ہ�����yk�U��d�_��Q���Xu�֭���z�lM�s,'{t��Wfv�I<L�c��T�K����*����J?�b�Ā��8��z�+2�����8�1��A\$�JH��TÖ�8��q�|��D���E�j:��׮��e������������f�m)K�`�lP�8�p��������nʯ=L�ڦ* O�$0�G��{��`l\ �)6̍���e�{��CO�qֳ���׾��;cφ���S'�'� ��i�?*|9*p�O>���qV�NǊy�D����� &���^�)z��$�Õ��X���%�I���"4]fE|6�:���(nv%�y,kt�6!�0�m��_�K����ȅ(%umÁ�(hW��)�:^,�-����P������美��S*���6*Q�(�܉��n������Ԛ�!��!�*��r�h������y�����7I��z���d��om7l�����L�tG��;Q��suJ�������ۅ�<�W
�t_,���sʥ\�^l ���J���,����W�s��c��=�EN�H�l���V��a p��d%!�����4��2|��'������нl��S�'��P��X~? L{���B�?��ya��Y��7��*:\Ų��2D��r��Ξ��"����i��L�r�o�K�sѨ��PL�=Z�׉���a
oF ����������dƓk�N�KS�Y�Ƚ���?*�5�gkt8c�����1`���Y__����z��@��^��]�d��_RB����5��(�K�}���oΩ�����xZ�
ݑ����-?(Wtޕ��w��2����I<�x�ɂ�4��R���>7DSS�M���dRvD�$�;BM��Fl�z/q�*ߐ�/`7E��0w�o!������B��a�̴urF�=�CVYVp$�eդ��8&�r��t�`/�<�y6�=1���U��nǻ�&���{���?b�Q;	]�����X�B���+����q�BV-�	��Z�=�[��z/��_�����q����j������<c�^l���A<S�[�T�
��+t���!����:�%�U�H�*�q����	��I�����U6�`��p�B8���z�"�#�IU"��i~
��Rc7~��kw�`$��6Y�u-a(�N���6fU�uc�2SxLrX[�4�E����}uz]��mB| ����8����)X���<5ar�O�O�d��ug!l��^5���2yL�ZB O?5{ʉ/��~�6�s�ǐ�)!�l�C�V�G�պ��C���u��MN�G�a���j�r�v�'tk�V4^_����x����c��{BK�w����O��Wmw���e�O��m���Z�|�lni���Cu{r�����I^3(�Jy��T(V��O �p� N"W㊇�0!@z(�����- Q�h�{���Q� n�r[b`5t8c�W�� k���%�,�/�d��
��	�BO���;��!�Ƿ�S�}�qTϞ�[[K(;{j�:�e��o�y��,x��BB�yq��`kx(�}�Pd�*�[`��~��-�\Y	+��ž��8>צ�t�K�*�]x�g�����}�f@�hh/��o� �U�%E~?��s�Z��|��^oN��0\��n�
���e{}�K�I@D�=�R9Y0�h���nm�oIM3����������Qy;W�z� ��/0а8�*�w>O��r�`h�1���5�;��㉔�E�d��a����S^~tVz/.�n��7W<�@����#���C���j�c<�;�Ax�|ʲs�ۨ�L��R���q-c��O�Y�� ]6]I�.�WRL�[TH����cG��",!���^k���`ʊֺ�V�B�q&�¿hcӠ9��;�.�B>��x(X�C4Kɻ7����=�ǃ�������f��r��xU[�!}ާ�@m`'������b�:(�`���&.�:�`�"u��A�?�>Z>$HӶ��Wn�#���:����A0�7���Y��*��ܪ��>=w8~��!�4�j���HGW���؎����sѤ���ڒ�����	S��7ܔ@Yd�|>�����Y,I��i]Q��x�S;a�3��}�9,~5��Չ#s/�@1��#�\�
ȫp�J����V��mWP�t���4�]�7,��#�,������^\����ڸ��@|� .���JBu�T!�dE�����fKoPkbo�Ő`c^9�����/$߼ÎV�����:i������&�Нcqh�Ot����V�ㇾ���1��$��
iHH+1ݬ��E/D5(s6��t�Qu���A�شrx3�-�6)5��I�:}�=�<!Rd�9K��5��N���'��B��iK���v��ᘘ���m�r�m5Q��{�i?�X�'� �i���]SBk\���j�h��v#1�y�΄�#_'����g��Zz�V��^S�%�y'���l���ʼ�pk���,�^q������d�F���RB�-�σ�h�� �\��|n�}�6�V��\��wYz1�!L-V/��a���&=?g��w���=2:*Jp����36P��ѓ��)��c� �^���A���]+���V�}��H�p�/�i'
�9Ʈ]d��11���h�>�벤�S1�~�p��ә@== �[6[O�:�"���c��T�y�I�!o�4�JXH�7�qJn����Ǌo�`�V�����s���r���l���ūtb�{�CAo|��������ox�