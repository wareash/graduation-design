��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2���"WYj����i� �N�7A!�@<e�]ң�;��5D�監p�.� ^+��Rk0;Õ\z�7PF���p�e��	��j�kdD/���1M���(���T�e+qr)zD���FWkV��������\���mk�*
`�R���	j�' �� m�cD���9:�DhT]�����۶�����i����ޙ%��d7ܷ��	�:���U��(�����#���wv�pFc�o�m?���<�δ�7P����( ��(�����1���o.O����BE�l�pSX�m����
'j�ߑ?�a\����3!���Dꁖ�0�S����>��"��M���e����2P�����H��£f�xV��w�������є�����k�,@q,[�Z�&Kp�2BП�5�O��>�2�@X	&n�탛
��S��P^�����'��c���9��3���^��Cԥ���TzYB#5߰L՚��ѩ�ӧQ���T9�:5�N��y�|�#M?�U{l����A����x�H�E�n?�1v1Exi�w��h"���ѡ_��v4��)����_%�r� ��[��I#�S�V���I�sPwW���/���f��-�����p�_���ςTJ�6v�9�+�S���a�?�j��=A�3���g	eS�?�����Ix`J��,�wD4��}�clX�爵4Q��wU��5ҙ4ֿ�8q$����^f'���oe����j4�9l�ZD>�:{*8�yp���^D3���$A`*2��x�괽� 8�9�j}�����4��*;��Y}Z�nw��d(���%b ��\�7��Vϛtz����pN�<����&���hM�#�+��=���6q���f*���S�a�A���h '��)�4��b!
�d��9�\�����'� f�_��{�)l�g�l�I���e�����ea��_%Ԙ�h���/�_-�oH�� �2�����W�0����������������'��v'���Dm:0dvQ?5|���!Ͻ.�E��,Z�����j! �M	���� ��ވ�K�Z��_j�ԗݱB�!��h���|�'���vwj��[��:�R~���3u{�Z�P(�œ���bF�	��;d)%�܎���	`��iG=+�"9rYD���B�հxi� F	��M]�s�y96�g�#��%$�.sq4�$���M������N�6�\��9�
V�&���۠��q��U:R�D�(����p�&�6ǣ�����ʄ��cu�M���T4;�X�y���ɢjϙO� $�n�S��k���;+��-��9�*w�<�V��)����*U��ܚp�p����fڹ�)[T��XF���w�$ߎ�X���w�E�,?ٶ3�v($: �@�g���I���0��
*3B���{*J�5�gļ0/�m=�2��#�Z��}�<��d%�����4���%�R��,;��߆q)�"��� �n8k���&�ђ_9\���b��rJ:y��m��%#o�y�Uq�W�Ke�8U�r�u�����c��S&�H�2��I�ү�؞M�U<S+��S7��'-�f:�5�_M�Uf抙�\��5�H���(5��ؾ-g���x&X}��P렍
�n�U��.{T4꽃'�#g��xD��(��bS���&�y7���������L��\L&�ɾ�_�%��#��Wʘ�mxZC)�;Κm䂫���������@��0b�\�Р�* _'�@�Y J�g��I�㸯 =���.�sr�?BT("�eD���^�>0���p�ZH[�X��
���у����� �b�"��m���s]��M�D����b��j�������|�[7%(��;�[0��E#���L��_�|`�Ȑ5m�{
Am_�/F_�Q�c4 �@����U��T�L��mB:�c�?�ٯ��<U�<�B�+֮��H,t=�Y�!��y��5��"h�9M%�4H���Fk[�Ϭy�d��ԡX�</R�i`�M�sC�C��E⡳�>�\�s��������N�� :�EY�?	�Ӌ�� �Y�|�����#�W+�l����5c��D*9�8������EE��:��c�P��D9�VMϒ
�A�����	��c9c��;9󄼡D�AH��g�`����`��p�g�5/i�ת�W]���Z8�N�O���yx�ug|I�Z�k0��-Ȃ����J�ԩ�A�a������U9N���1�}c��KgQI����Z�m�k��'��d����)F:0*�v3"L�)$P5z!TW��9��.f�O|S�3�m.���]b]��I��Y[��u:g0d+��S$X��l��^V����P�E-xZ�W��}8�S�ÝF�
�j�)3J�%� �m�4N~Qˌ&<����������s}��1$E8�^ �?����!���h9�
�mM��U'�C�B��1�1�^Q�>��D�1��S�'��+m,'d �ͱ5O��蕎���ަ�\���4��?��i��};������Eo�i��g>���"􁣙�ߧӦ���?vٗ��:����]o�i:�������væ�)KӃ\�� 6iҹE,�Q��(l�c��*���^z�^��0V��,�퍩���^Xc0z��G=짟ua����M)��f��
	e����h��-��v���ku?ڦW��s�]�3�+l~��)�omZs��=��Q���6Τ���K�:�t���ߧ�.�I�I}�����:2��e,��f���T҉ӭ���O�t�F��[0�U���(2+�Pm�ګք�U	x�-Z�i}e�~�䕥b��Op��dJy�;X_�����9�$V*���(�{�%v32�&g�vsEF=F.+���A�a���1G~j\��k(�t�l6���C"t���7ζT|��XO^C�/��K?c��1�LH��~@9���#�.9�a.E�\��]�h��{r�e�CS��>�xΩ���"["C��| í\C�l���k���F���+��V�5<�'2��@�M��̮,��o��8�EI�מ2��� �P��#�Je����qޚ��T�y��g%��-����t;���1cGؒ=Pڞ�6��	:�9�- W))\?Da�D����֭.eU���ž@�\>��5Th.|�q�>�B~Z��6\ʊQ�	��xȴ��x�ڈ\����K��?f�Y¬x3��-`���C��t��������CN(@Ǧ�c^�)َ�K<���)AZ*�d�BT����#O�:���7c��Rqf��s�������]��Ӣ�qq�Lu���n#�;8�Yvk�������cN�l��<<? 7��T=����ґ_�e�^m�I՛K��@�X�#�4Q�^t��5��̥i�U[!h�圁R
GԬ��t�?���l"N�N��t�u� �&?�r)d�7�Hx<������4�*��J�e�3�M��l6A�t���hi���dJlQַ�D��ߺ�\(J�&�����Z���Xq��ry�Xx�(j�nt Rƀ�&d�<]f��E�eM� .�u��̹GS��9лlo��OH[�4�ME&#�17p�W6���,�����e��˚��ͧ�T�'o����J��#��^�>����-kp4!�6��:��������额�k�܇#��8qU��t�r�L׶��;��+?�����OxXHJQ���'��I�������L��è��s�U��a�
��	�!�~eu��CJTK���`uɪ�Ɇ����5c!|܂��H�L}��'|���D˵��Be� @��2w���f��N�6hN�m�'*�����H��A��5�`��]�dA�����R�Hs0f�!�7��|��7�s��+
:�P�G��c�ı�R��B�V��o屲��S�"�륊f�o��g�/�ǁ��c��d���9�ݛOI�=dl{q(3���/���8�W#>�>g?��C�7K-�����'K5l_4{X�'��_�O�?��Ǻ�����&K�m�Ot}���,;���Ʀ�7���&�H/��E.�Lp�����T}���}+m�F�&����-�c�5��}�sUc�����ڷӴ�$�Q��d i�S�7��F� ��6c�)L���i����X�������ŅX���� �ꍢ��n�z_��|%r�
��3�7ܼ,���&ĩIHY�~���p2p�dm��K�\y�3��"���ЖF(s�<KÐ��4�T ���r���RFb)i�e�bg̋y�������/%��v�:-�	�����sP��Ƽ ̋����)�۠!%�*�@����#�b���O���1U(d����x��v9`��)��]��<'�-�#4��5�����.�\�<�
୽1���{M
��Ey�	T��N8�6�mn
6�c�q���J�m�����&U�C,p�Á�n~�tx�R��ٚ�y&�ʫ�H@{�L�d>u�Awz�l��4d��A�Œ(����Q̺9%L9�!9�FW��Sw�^N�w�qi�M���<x��Mw�!,�
%M��N�i��4��݅��L�|��>�u��� @x�N!�!�z~�������
F?2{Sy�b��P��痢U"����?�5��Cԅ���&t4 �@�C��m�(XKI~f�x��,�\Q��!�+K����:Ao���v�`�z�^��	|B3��������/.��aܢ��`%����P����K�<��'��&��;���W&t=���^�>���Ov��pz��L�v��R�Vo=�59&*�m{���m�RbZ>��;,��𦘏����w�A�6oe��ףa��&7�v��i._b�K��u���=h�n����{ᳰ�JTT���:�K��9#�_$��c���� WNv\���6�Ö	@��?�*�)/��Ĺ�/lGml�����ѮnR�WF�L��5��MO2����(0�fX@�jY\�:�}́��C:���~N���Hi�I�w��誽S�ze	~4�F����;Rj]�e�kk}K�����Ջ�4
H!Xm��VTr���1r��p}0A�� �ben�id��>+�S�l{7;
!�`}*�!��מ�s�K���{�x��\�O+��M�ǌŰG3�H�+�>G^{:�:jDC��֔+b�ˉ�ޙ�dpL�:��~��.7u�& d 9͆L>XBn!Ҏr)�A��2��%W��V
j�U{�d(�8@����_" І���ϧ��������?��e	���#�|m6R;K��"�<��}J9T�F���0 ��4�,$a�f:� ����H��G�s�V.k'����x����&ѱx0ٝ������%gR����H�y@a�k��"朜�N��(R�=���g��A��'��6���8�R���5�Tt�{��*�$�f�*H.�I�#�Ϡc/1�,9�;{f��(C	ΰ�%HҺ�B���y��l��}��ӝ�'���=,2a.U������H�q�!�>@���2}z�u:E��R�DOGsy��r�g+�;�n�LtJR�
��f�M����ugB3�+����fϦƻ�F%3�4\t�*�h�Ϭ�{!-���m�<E��<�|ú+w$��'B2�$໿�Z;�'���cO}
��>t� I�� 9@i��\X�?�b��tjU���Z���hm�-Rc�v�nE�A��{��+B,R`@�r�� ҞM�H�1�X�a�l��������?�V>E�����i!�_��H��ݜm�b��[�H������	B�Oٴ?���k�Lxg3r��ݘ� ��/"��>��~A>��?T�`�$� �B�PY��b�=C�}��T{�Ź���! �DC~̖�_��_'AUu��D�Xܧ���ԋ�|U;8
��up�!��Ӹa%v��8l'����^����6�Y�	��� ��*�6�)��_p+O�L^)��>���A#�c�⠟�i�L��a�l;�rFsb|@H�A�Ux�HJ�Efj�w��d;�\��r��v��(w�l�v �tt�EK�L�sP�c<����jv��;d�܍r�}:�7�K�4����%W���P`���C�as�|��|]iS�U�W�Ɖ�\���a'�� �5M<M�0db���"�(�!����g��i&:���i�J�0V�����ؾћ����r}�Ք���HI�|�T�!�Pԭf���	Q�N��]�C}G{�Lm��o��GQ���k7�M.!9j�uOL���p�gy�-��y�y6���1��&�)�"JF�#�_��ی�5��ovMr�H����U�, 1@ �+�%:G{BI��C�&�+ ٴA1*pѣԯ�q��!.-lj.m��!!߀o�Z�S{G�S�	�����R4श�ͽ�	Ή>��7�e>��p|猹ͳ�pC㿰��w5����w���ڣ��T?�������7`]mCk���k�bzCσ�N��˻@}T5�S����.��N#��-|L{��oN��, �'�lR��-�l���ۤv�Ld5=������G�}��&5�/yO�_�Y�Z�1�L�D,O~���I�)�f�6�_���{� ��BYC�ۡ6�c��
O��nd����r�%*����"�D<�`N��k�Ķ�&���:�<:P�^�^x�h;�Y(i`�J
>&�J|q�{@��U�'<��(-���c��FPՄm ��_��z�ϻ�U��6�px
p��n	�z����%^D�V��[$vEhe�s)�us�;*u>�e�A�͔���8t��	�|8��-�v,� �j��v�|��(�-�.�`?q�`�t".��3����l��P�����3Jb,H*��B��}��ЎI�V���l� I�>%Ŵ*�O��շ��l��Z��`*ϒ�d���炮�Q��g�ӞZ>P���S�pU���A����Y���m#9�����s(���*���?�zp��F�[,,�0 �;�8��d�����A�j���������b�D���
�ܧ%ih�gW'��1����e�KD�C��͞��%?��F<;�'�W�c���DW��چ�N�������D��_n㎙�>'���A�S��w�8��z�y��J���m[~�~(v����M���n�EKi
�0�'V�K��?�]I8�P��p�-Qy���hY�i�Wv������\���`��0���8����-�}��jTb��t��(��vѲ[ǽ�+�!ǯ����� �� ݜ�z����;���J�o��>���u��汉��{��d)R�Q��	B�=�a�4v��H29>�����l �Pþ}-,+�*h�b��_���o��`ɧ�3�Q�܎Ɣ�6��i�ft���aǲ�.���B1WM��2̈ �2 ¬�k|R �=-̳�+�.�g��j$D���cͶ��'�O*�_q/5�t��?�*ל�=�0̮���}7 ��LD�=X�g�"դ;��@�� �ns�W�R�o,��:w�=�S 8�r�i9С���.�� ��뎸ɉ�|�f��~�"�����i�ݒd�ne&�ȩ�I��h���\��̻˕F�s��=S�=|��
k��,�Gz>$�D��qY�|���d��������l7t�ɔq�d��W�V�:��eB'�RV|n�3%�H�f��w�������?_K#�h��W��YE�{b����j�/he �L��U�~ޘ�x���� ;JD��KC#�jܑ�5����#*�$/J���n��]����4S��03jł�+�rG������-F����۸�,����=���9';��w�3�[
�N�3���_�E��=2��"YDz�CI�KDLg*�5���ם���=ՠ^c>xD�ǧJ��V������f��O*�Z$20Z�w�GƋQ�L���,\a����`5�X>Mf?>�'KL�M�@�z:+EB<%��+x���'X;ק�h��w4��d�+�=fg�&x�&.2&V$��?� m��{�G���9�Zd�v��I5>a��_tG�	ʠ�1`Z�)��V�S=h�s7�J�67q� ��\`P6�l���K67���Ex	���ձ꒒P�����Q*�+�gU/Ϫ�>�Ie��������e�=�[n	��-%B�P�=����!ܯ5x��Jk�d�_{���_�v������&(�gq�B��2�}�mU�G� [e��y�k�#��·����7������n��J��<���`+V2���	�	� �D5�N��`�sz1hI�g#�Z9*�U�9��8��չ�g��I�H|\����Wr��CY���t�NGg�Ɉ���|�sD�{��}�FP�~��hUvz>��0.Pm��'�	�H-}�a+J{�A�S���n+P��B2�$/E�6f}�u�A��8q��F������U��6�<�Ҩ/ɹ�Q�Q�5��61\;�wu���[9���l��Ь�h�M��,l��E�����LI\̔&hoqå@u۹��r�=�u`��3���v���	�|ٷS<F�v�F�~J�}���pFy8���1�p�ʯ���[�sQ����S��h��^<os�O���N�T��`�dsNSD�r�o;��!M�q4��m�`���RPV���=�in�aNY�{{��א�]$�*����D���;����iG�H+S��fČ'�������Н�l�dӒ[������/J�4#�Nع�uE7�B���iw�B؛�#0�L��P[��l�FK�-TB�5��YYպ�%� -��ៈ��� d��������gL�f"�hYv׼��{�����YR����|���K�x�:4����K�@��bw�P��v��Y��D���P!��IAѾ���4�e�T�U��u�ڛ(9���4+����<�-�*Ʌ<_���#��N��BɳA�B�6%׌ْ'��.�����73�n�OԶ�ѵN�3���3
PMa�T2l��?=M��S,)�t�jCc7�zvY%�E�1QA����D��?*k!�]�6Fk���sp��&]��U0�:��'c�U�m4�}k,�x^�R�Py�c.��h��:|(�ı4c]	m/;����^���]��f� ы:xMx�s:l�''��� ǜ�E�Ł��/�b�e�����ֳkZ=��洤���x�:�_�dZ%(���ܹ��r�e\&�"�2�̊�Ev$z�qH&�%l\Ӽ�>j�9t�4nڜ�.Ǡ�4^�gd��m�|�D�8�)���vmM��{�����0��(�0�H :�� �hv*Es}ٛ4�<)1w�̝8{ë̢�}Cqd2-��������>-��ne�bc�i4�j$ߐ.%�I9��E��9�HƯ�*�ي��Sť��OǬ�����
���-�I�@J�5�릈Q�Qm�|9�M^����A�u�^�൫�Tr�8�΀�S�p����tx�nl_ǵU�V.5
>�)uQ�g#�YCsI����_%^j�H�+T7�����p���H�݀F����~���8]S.`����&��
�����4�K�Y������͋���r��}��gx#���Y��DY1cߌ�7�)_R9�]`2lcګ ��7��ώz�!X�wt]_ˇp�N��}�WGa)d_�Ĉ��眴�U@o��)��V-����%=���}>�P��! V�>Z�'
$�Ўz3��[0�K��D�%��'r.{>���a]KE����t���?�y��q���$(�MI���eө��0$��)X[�:���z��@���.
mG�)��EM\s��^��r6�1TcP��q#W�z�09?��yʎ:�4=py��2��ܴ���Bz�D[�{$�K%I C�"�fU� a0������c]q��!tm(�}3��Ě\DQ
�k-���^���Ř���{(V��y�$�_��� P0z�Y�5���B�r��ؐݍ)Z�����p1�g|����w�'v��ޮu���ͻ��{��[�:�j3i�Y۸��9�'��YC嶮1��,���)4��(q�vR��ϒ����x+��u�(%��u�$l�j�*�$�#��&|,���X���vπΊ�7S�A�k�����������h�c>�	�+�XH���~�ĝ�.�h���n��< 7�OS���QV6	-��Z���3�I�#���"LC��*���O��(��{0A�ϒE�M�x�hQ��Mz_�����U�;z�s��S��}���lkF��A_���R� ����}�U�i��&�=��ߥ����yrT� Vl*�]��@{���m�g'-I�*Ė�E#2�X��s��;��E�	U��}3Z�*x�&�JGj����緌�>2�%�Rtwö�A��`U�\\�\���Q|L&Is�\i'���F�ӈ�6��x:�E0�W&��u {�\#e*j�Y�5���]���n��~�EK+�I�t�!�Qt�G��OŦ�O|m��Y��������g#y�����J&���?mﺴ±'>��� ��?�V?��D@�I^a�D�ӕ 2�´䩪���ȨU�38������������@\�G�?�
v�����LV�ִ��(�����^\}�Ψ^>)�iܗmhI�z� �[�E���i��C�1B:�A��:�-��]�q�V�3A�����	m1�M�U���t�&dN�_��qOb1��")M�/wP%q�W
��N��'ih�V72�U?�^�z�Kܛ�3I�����&}@1Cv��D75��̘J��M]��H�P��^�_Lu.��t5@o�^b2%�d�.)촮�W/&oA�Ú�۵B�E~Ee�$^q�G,��֫��u0��
uL�T�I��c���{���΄l�K)�m6�TLH��.�F�ҕڏfNn�Q=Ƽ#��Ƀ`��
�o3V��oZ�hE'�ɪ��}C~X�p}����[�'��"�@�)m�wlkř�u��w(���H�x/�C�օ:�+Z-f�赏Z2e�]I?���e��w�C!�_J����SI�_���QL+�e�4f�2��zS�H.M4Ҟq^5���^6�D6��-S�@�����|8HwH�N��l"=��5����@���֛Kr�����KK�!(�,wCߵ�>�8�9ߧ����@]�U�]u)��6_vA4�eЊӑO���>����
+s"�.�ɼ������2�F�]8�7��_�?I�ec%�G�)ċ���.!��X����&�����,��Ό3�R��#ؖw޳e#�^��a�� Li��pů�� SjCU(�F<�յ��R#k�5���K��^�Tu��������n;o�����2�7�br�-�������Ry���w����SvLv%IW���f9f�=���8� w�n���q�/����a���3��#�y�|�?��c�b�X���	�GI:����}i��$�)tz�!�WF��
�nP���A_��Z|��+��!"4�lU��W��d��vPDb����/]돾.�9��m���������%:ZxJ`Q1� �|[���L�t����f�IX�a��'�#^˄ũ'��K�D��)�ŀM�|�:��fkԆ�?r"�Ŏ��x��x�^�@�DEc�fFE��z뻀Mj�Ie?�ɽH߽t�3��2eh;��=��%��U�_pY������3nL��Fn�K8���C��s].N�a�m
�G�4&���y �뗥�|�=� q�O��V\DmU+��X��O)=䫾}e 3��@�8i�y�\_�H�с`%���
���8�B ���;�(-Of	SCC�=}vEM3+ ��#�i=_Z��dep|��KJ+�Ӱ;��$��z�� s��D+w:�aU����P����w�b��n:���$r��=)���4��2K�V]r��m�����	F֎��$���7����䜬+G�3���_�,�Xf�a�y"�3�,h!�0���eNXf��/<=�P�ۉA��H/�2�����G�7��#.1�^��Տ�xD���_��
��-B�#��H�c,�;��)՛fl��ښ42��@�W�ݴ�߿������*���A�m��ƒg�j���g��9Q�75���]C^\��%��󕊺!K�2Mi�t�JF����N���=�S��F�K��ȵX��k�
�/UEڋ��AK��@�K�57�4�?c�o���Ǖpв�;���	L�����­qMD��I>kg+X��xJˆ4[�@��)u��$D1���657O��;U,Ĥ��_�؏����|~�t��$k�B6]8���ߝ5�PfKѠI��Z_�H�D45v�L�7t�O�?�EN�Nrw?ǟ�$���տ�$XM��"^ʆy(���W�E�3��]�Ǻ��{��Ή���uO~*�Nb5��, 6����T��t����0TG.��f��5���8���1擶���&g������V��7oPL�d�*�U�ѵW���m&4>I�֟X���G���Z�]6@=��+Ym���ͻ߂rF�ı�� �d�1���B�ԁ�G:?�
M$(�r���j@E��G�Q��H��[�ȓ�h`<6(�k�f�Oa��E0������-�q��۲��~��i5̨���g@������A�ht���xoW�����w��Z�����1�X�-�@��\���f�GT��
���Z؟y�>�t�xD��XiZ-m��ק��V[� �j��k��n���B�;���Yy��������4�%���@�Ԝ�u�"1��ү|v�&��8��59�ý�*�°���������o�M�Q�e�e4��T/{4
L%ML�{9K~����J��D���6�P x���dء���Ǵ:��$��h��?���M$�=�d�XmJjK���������������C�+s�'8	�
Ͳ�3��L�a���I#�� ���9�¬��O�)[)̯�4}�����[��t���m�D_k��v2��I�o`	��m����j���^ �OǱh<���j� �;�HDC)⒇�:���S���!F�����~%��;�Au  ��ڐZ���������0|��o�=��r[�i� DVk�f��Τj�s��i!�:��/���ЩQ
�I�^�� �TM'H���Q<,�P`� ��#}��$�v;��O�]�h��,Q��{Ew�x�����kn!�E�ϥ�c������$�*��f��h�&3c>MI��v�v�_�sů½dq�����f
��gI��֝1ˤ��9��*�y� ����};d�/�VB}(]v)+��H^���a�����ї�LeE�f��nW*��)!��I �����DV�b�o��F
�j��`� iT�����52�o��}� ��~Q$�͏�/����%�L�׫i��-����7r�.��c�Rw�����������9�h�4��&�E�L,�|f�G�3�ɩZ�h��8�N-��.� �nU�Hɩʪ�o�
���)�}�ǭX�;�Svn;m!�%�:zPy-�#h�,��r�G��,�ݔ'�d��#W @��z�?�2�5b�l6��Q��>�ܼ�ƹ�)��1J��v��!�uD��%v���� �s����C�T(�H���{&�|U~2����|�u�� h��K� [#��IW$վ�U\&ZK��T��^[@��x���Gnv��nؿEuV�Y��#��{�o&}Dbe K+��;¯����I�z����C��I+�}	{��V�J��3�
BmO�(��H��{<VA�l�ow�}�*��u�S�Sڮ}��[��V?o;p�α/0�4����ؙ�{g��*��� �h��/��T^F(���@�����?������̭;lM<�x�^*�}<��X&c�58��
��P����j2�� ��Q����P�TCqQ��,���/	d�P_e��tL/��Hbt(���lYx;	'C��������e8���^����D�������7�u�������\�3 ^L���d�|L�9hC|��)G j3X��UY<�i����uؾƯ= �b7�ۋ��N4��5:�
�����]�c]�OIl�M���a�TߺC@��2�)���9�6���ꅾ$��8ߏ_�H:�#��0�hIt����>�D�Y��D%D̖�B?��/f�"[���ZO$�.��S�՚�
�hOk�����Z=��G��= �����nʐ�:J}p�_�Z��_j� Q�*t�4����'ff��~F�;����xw6C��I�w��R�M(�&s�uB�C�w���P$��u����C��	Hٰ���^S&W�I�]���(�̔V;�P������h�������nR��;��?u��w�j>��rc:�]��������;Ѱ�i�M�W�Xn���Ε��S���\a4���~R���p䈨�X+�뭆������|&0����s�f�Rn�a7ւ���k����d��� �s����������́�>�z� G�e�ն�%�PCfF��$����N�����VN��s��z}>�#�!;'�J��"�,%�&,Xf
��F���Ab=��%0�]�1G^$!�)���*[FC�^C��xi�TS�R����H��}��P�{|�,}a`��V�����?��|}b���'�쏏!����N/��PL�o+���d�\y�K,�1�;g��VǓl�� l���L��5���e���p���g�� �S ߮������&�=:�q�.�z�XI=(�~Mlm�[�+�:�������U�T�}�?'��%���*��Aٲ�?��p8���X摂zM��@p0����UW��%�4����r`�;{7ڮP���[����#N��͔�D�s�g@�3���:�t:d|�ͧ��Z@~�"r���}�X�^�O�SrN��i����Ũ؛ގ���b�qpf#�Q���HS���R�%��o����k��"q�� ͚�����ɕ��:t�Pd�"~�B֓�gn5A����.�dq.6j-�RP����5�A�U��i�Ǖ�����1����y����$}�
wB����c#����5o>H��d6;�<�I�1��c[E'Zb�;�G~}��r���ƨ���

��������u:�(�$�Vt��<��XlJקZ��.�����@:����e�z�X�n93�)���Rn���su�����]��j���ǈ�Ek��e���N�rbb0�
zܳO֊I�LN�����G��ד ��Т�$�R��o_����#��X�/p��Nb!���M���;��lc�f�a�ZU�X!k�S���`�?��0o��Iuf��?
��vx����	ӤyO�j}���ZЎ�����_y��>�niu��?u��#�E�(���m~�2�!�%s��~11Tv&����N�&B0;G�S������zhbSWJ�Y�'�rlE�
�,g�KQtՇz�Knl�H��sP����o|mJ�G�n�gU��Q����KaqOP`kLp�Ă�p��1�*(��5�x��Շ�V�tإ��U���r��'�[T�9!/Ъ�K�*��	�R�1@�r���G�F����}{�ᗭ"�����
���/ ߔ�L��<���|,2�-�P���3����vg���������{�\�G ��ʙmF�*nҩ����)�ٮל��V��Sn�j?�A��	qc	K�������W����#r=e߄4/��,�O���|?�����c�� �q�d�Y�����ǆ���3V�_�b=<1�I$ޅZ� �^\&��Y�E+l��I�6뫾���x��i÷_xN��-|�7��	���G!_��F:S�ZQ�*\�3J��
St9=�m>{�ؔ ��d�߿�d<?B��\���W�a\���2��Fwy�q��$!V��
�������|����e3{�υ7��c��	4>���\.�G���� [C<0��`5�ⱷ�Z3�f��oFLc�P�뜛+���o^�L�ׯ7�}p��_H�F�9�4{���,�a N���3�ܨh�.�k΀i(B�%`��u0E1D�X��4��#ۡ4e��j��{9^���$��� ������3�D���gEq�~�\t&r����Hȝ ��T�3lZ3EP��Wk����^�<�ʾ��|}c�y��7���v��J�WB�v�Q�3���6|�{9>(ma��ߴv�=&KU��g�)�8d��<a8����V��,0QXLb
|�ySzi��(�%
��T(I�w��l�X�G�c��`��kl(�߽�R:�aw���#h�l�N\Z��`���/	 ��8e���\�zCۓ��Mwt�վ��IDCjɼq�����p<i�'p�y��6-������8����_�����@����vzr�k��)���'�+�k��i��%��3�}��$����o�-����
���C=��&�?7�Ɋγ�Pu\+��80�|>���D����Z˶�lK�Txϱx���_W6�x��|J5�Whh�1�.���'r��tL]�7��]5����u�POz�Q���TZ���m�+��:#Yх����oV�)4��|W�1wF�u�V���(��-i��NN�{��XN{�A}}�:nv9ߝꓬ&������$�]�."��}����]��j�xJGH�]������^��kZ ��C�舫R�l蠫��ɣs����6%�a�#]U�
�p�m������R�ΫS=�^f=^z�@{�bQ���I.�rE�Euް"&�r�;�@Ơ�B����i��&��D��,���~t��\���c�!�+���`ڟDn\`s#����Z5|T�C�K��z4C��JE���2��T��8�_!�������N���d����f����cJ����u�Esv$�܎$�.|k���|j��j��V�j�KsH@q�(L�@���� N�u9j�2�<�Yt7�{�����e[g�s;z�������)=Tz���]��{������B��K��i��Ħ/[T�N��p)�Ʒv�=�v��ᤜ�����p%f�>)<{���>1�)�]dLk�sቭg�����E#��e�e�ㅙ}�g�c����_>�DT��>��F��Thn�1���~���ą��G��Z[<����KoZA�L���@�2��q Ƽ�Ph�rM]�I\a��C����h�>�t���Y�Η�5�Zn'Oԯ;ǟ=��Mp|�n�D�g#"�>G�o�3�4q�he�!<��{q����ƴ�˹��a��_t������Ƭ�=�4�HEl�%��8�J��8z��v}�q���X�t�J���[�	,��1��1�i��#�&Hf�	3c,p�E�0��4�~W���u^�I��ٖ�V:=�`	��Rץ6=�h�@��.2a����_���>�C��Е��n$�z03�7��qE�F�s�j�R1�Q��J���#�=�t61�'���u����2uʬȮz6��Mn��0d
�w䞋$��1&�4e=uC������IT�"����/���}���h��BN�4\y�^��&u&��&�۶KI�2쥚鞫��cf����,�p+�L����ސ��|�W�������Uˑۨ�6������냔��H��g�L�d���������j��Hj�R��F���ɽ�������+�1>Y�'ҡV<Ȼ^E^��r���!���,���7�`�MM/Br�"�K�+��c�2!俜z~�2���j
�����#~�`�Z�����E5��P�W!�[�o�I��9���
��V�If�ܑS�D��N�ȫޝ�16��^o���ڿ��=}@��rI�z"��`�����d�\\�zE0IH����$=ӞT���Z�`�ٵ?��$���8V!1���Ej�������u�����H6��YZ7�t���k8�OZ��<�3��&���j��c?�R�^:���N��OQf�J�4|�l`{/�W`�u�4-*@E�g��uzȄ���P��.|2R[�GA2H�	�ݏ)��y������������2L��ǀ��<���!b��t��ikdO�(	ܚ��:d��[�]D&om�=�Лx���r��M��$d��x���5 佳�\�$MA��
~�>�3�e�p)�����������,�5?I}g(�ϣ�S:<��^���;�nh�h��6��hV^�7�h�1�?#�pO6�����	��ܣ��|Dx_P�����|��t!9���_z��*J�����{�����������P��+{��L�bD�?I|? ~��^��3'$�����x��ڼ�\CZXгq�۲��iO;|,6����͝�ErtV94�Y�
�o��ϐ���x��h��
I��T�Q��N��axx�%�EIv(v�t)�Iq�*�6y g�jlmf��{���c��/X�q��
�\�ony��$��ᒟ	���.B�C�mh���1�%����0�-)M�����WY����D�k�Sc����S֨����ť[�b�/>����0��V���t	6�jM<��i�\黽�Ԏ�n�(�5������E>�o��m'3�B�{ �/�C�����B� ��(Sc��v��<��}�,�%M�֠�*u	�>������`��B3�j�����# �\ZL�-8�yZ�v�4��>��5�Mrb�]�H�����-�e[��>Ә�~�X8����{��M�;>Ѡ/�����W�( >��J���
��q.���@�-�#���?M�N�l$�q�#�����To"dv���*�,���0<bPv̲��ؖ�"C^����f��2N�N�+����l�#��Va;(���m���&ހd�Y=o>f�"F��Nߣ�['�1:"�};w�a�m
��lė]�	��$�ɃVc�|M�!�<���Yh�n�l]5��m�|9�jӒ���`8�������#0�g�9���'.��|�iP;�n�g��&����H�M���k͢�!�*�������4��Tَ��4�%�"
ׄ�{��ClX���/�:��wE�xHe�tbe��&8�;k�҄r)|_�Ȼ���S��P5r͂h��v݂��樂#�ewF���y�=�v�˼<!`{�^J��@�B�v����&	c�8�V�NXQ �ڇ���L�u��+�ذ|��0�W�W2�PZ�<��n{�\6,W�]�U��z.����2;X�»:���z��|�S?��/���(��*0�J2
u�ݷ`�L6�L� \��Z5,1*|�o��`z4jX��:��X4�\@�[}l�]z9�NǨ$������+�W�[\_ICK�[��F\/�*X����ρɺ��˃R:'�M� �d�cme��Q_)M��W%(��U�xig���{���]VT���O>ٯ~́�:���%�8��Z���c�U8j�Y�U��$��.�$<9�a,��<��� �R89�e�
:��n�x��NȧԒ�RV�=��;�<wq��s���#ّ�J�+e�������l��Z�&�'����h��-/�%jsb*?tZ�&.vȐm�NUW��G�%
�a������P����=]>g���`|�`�hQ���(�Ǚ��ƌզϲO��Øc+�*�1o��<u�T��"�S���~�oc���Ls�6�|�#��]�yՎB���l_��x��e�z�cO/h���dq�Q<��W���}>~���<�=@|=�>��|.�]^�HT2���}�<zN�M� 0�}�!�=$����V~}�;�������r�@0/����T���@�8�Y�c��@Oά�F��	�'S'�e��ci���m�3�=�a�'L�ǜ��PQwJs���v�֡x&t�.0��	�5�ݜ���m���z�\�f������ �\���QQt���φ��`WFX���,�� ���B�>��+�m�/	;�_��<K�`�����O7�*�BZo������>U�0Yѡ=z'��h��%����y�뱧&>m���I�6�i�'8(jg��?�C)|���?� �_gD�!Gȩ$�&�?i�>d�H����� ���I��i1����5���t≯��l��^,7jX�!.i�~I�/mU�B`�� �_��w�����k�aYu�=ׅ�α8�lt����5�>��z[$݁����k��Q;�P��-�TB��R9��D�X����.��,��i���V6�dR�j�`'	+��h.:�K�L���TOy/�C�&Ɓ�F�nk$��/�]Ƚց�;8����}�S��V$meOHWp��>m=�#��Q)Zw��S����F����������r��-�m�ʍ�Kȳ�������������y,$���C�6FY� o�<��7�Ģ�He�i���U|�A�\Z`+��8Xq����_��� ��YX3��l�L�߇�o�Q�{�"$�)�"�H���F���rN��M;���s�MF�q~	�Ձ��$�)���� u��M��-�X�'�qȉ��m�7��$�߸��jY�V�~k�>��]|~��{���H�([�?%,��4@d�'ixM}����̤{_���;��#aY�\>I��*ujI ��n}ɬ�.{�.,�������{u[w �g��&~ӊ�?�"ь�Cs�?{USnK阘��E��X�,\�` ��&����<AL�،;��o��e��I?��r%?��T��{g%�ɠto@� ��~�l�/.=zد����VLuB�Z5��~4��ƣ+t<{�nV��N�����H��c7� ��d14�>I۾�˟�t�!��щ)�Ę�������Ї����x�{X���xYQ�%WBx��N�ݽ����𨠿�O�`j�{W �/�v_������@�@���d�s�{�N}�� FN��s
�!�c���p��NJ^|�p�f	B�����|Sf>������>7��