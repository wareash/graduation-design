��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jåا{�\�u�?߷�dn@6�zf��r������;$VF�w�������Nd޴�\����@`���ã2�1��:�VU[��[	O�~M:���Ta�Ty��vV�^�xF~�E�rj�a����8N �B��%�>T!�i&NH�$'=�CJ��<�u�牣P�q\H�#J���B�m�qCM4�AF�$�P5�D����BG�*��WIx� $����X5:�t�ΐ��k��MWq�L���?�m��k����\.ٌ�����ytpv�ZXZ�wZI�������S���CSVp�֞{$��Df�&D�i^�`�_�rZ���	ر]���Xı^��N�;X��39\C���GƛJ���j�D�t�3=��㆏-�l�̉�� �p�)"4����v�/�Kf�L�΁�JCTfK�l��@ንr�C�8N� ^) @g���փJ���IO>s�'�0L�-K�^A6c�������_E98Qr�3�2=�lgl)�րO��p&�,t�Sc�ո�D)��zM�4�Ń���*�ig��R�[|/�A��	�yx	�J_��/SS����r*�c�8^S4��P�� �;��4+�Pъ��y���*4ө�iWbY���q����N�`����G�K·���_o�~睵�Ⱍ�~���dQbG��FTtW׍�5��GY/����h.�i!��q��e�l6n۠��%4�t����_�(���0�O���ku���r�e���
�s� �K���ݖ�F�V �5.]�+���"��\�
HQ䩛X!�9�(��ݮ%%�<�N7�l���>�I���'��#sK�c&q���]�su�7@P-A�PL�YZ�����QnY����$F�fP*�w\Qf3``�ehU�J��U��eS�M(*���}[#����V�>�^��G'��Vs
&`+$G�>�̩Ih�1�~��q�":9����' ��R�*ez���{&�,'��F��j���!a�#'��C�z3)@>�����3��&rV�qv@<
����~9�R��9���7��'kď)�XX_"�>[L�i����,�d��A�B�s
�*"[�ҫyk�˪}#Э\g����4�l~c�8m��"�S���؀O$����~7�E��H��4�v�x1���E)a���9��������l�@�X�:��sI���ZY���Ǎ*�x���T�ȕ�1���j�x�
���DN(hj��9�6��+��er	�׀t+er��k&��� t�oN�%�;�u�_.���9��H��nr=�'�sP��Qp,tjRP�7�?�ը���)sW���
�Fՠ�\%��Y����