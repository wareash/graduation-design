��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|/K�^!�� �Ϊ�I.F3�h�]D���� �1x�ϓ�k�K]b�ec���9�̑�2�۰�}EW��E�aǧ�b��S��+�/Aė �d��׫�~^^��y�4�4pjTK��~<OS[�EI|�ݾ�wi���tW3|��.�O�l�U0>�����զ�@��������L�3X��ɸn���'A��U0��f��݄ �.M������ZI�>Hz�����Q�C��ׂ����!l
��W6*��۶��r��6�3�\�^ף/z�س�����鵉�˞CV�MC��	��FKX()��fb��m�cVF7��=�#T�'�[QwB�/A죢,�D1�I�f�;a��H:W?FCP�C˫�@��"��o�t��8���,��4�`���c��1S�р���n�*T}�ΛnY�ptX�ͮ�� ��r���(��|W�=��H|��ǐ�=��Ƙ%�|�&��&
�$+��~7�1 >'F2��`+P F��o���`x	H���s��@�=븈L����٭J!�+F�0��Lko�<�ѯ_������-7���蕹/�sD�,$��s3�q\ဩ��*�6��ۄ�벱�m~}u>�U"�%,��l�)_G(/vZ�E݃�J,i)�k����>E _�o�+M�(�{���K��������_ĥ�Q�nYk�N�un4/W�G��$�s���5�s;�s��<�VL> $�9^Qw����Wh����}R}7A�����^D���9$g�ONoY��0��ۯ��64L���LҔ\92"����|�6~:e�/=ȇ��E)�u8�!�\�?��@�OYL�;r��=�͸�E��N�C^�H��d�MiY��q�#�2S�{5@m �&,����N�0����*�Z���̙�FC8]��2ƭ���o�*���5a���_`�8��̣%g;��mre��0��H�<��w�Hl�D+�*ku �C�F�%C+��ewD�ӫ�b��z�a���28�b1
F�z��f�T3�%�uP�(��_�C
�O�p�XWoΨ�4���^���v�L�@(��H ��$n��:*���wGe4f{���f� ����XT��'G���DU}�<�.�Ap��/sҎ��7��������הb֜i�S��u��Z����!��u�w���2Ae�e���8k��_U���yf���6i��U�����xd�Od-�/��<�K�(�(�������Ew0���o�v�e\���ڑ�5���(���zywE�&^%�Hb��T��2�;� ��~��a=B� ��/��_B�FF)	���O���o�;���d����!��/��������c�C8Vh�ם�^j�`SF�hB�J���V�h�|�%1��n�x0�W�Zg�'i�q4��mt�$��?�������mآ=6J�����O�~l�ۢ?�'V����
����$~�����"����տ���@SS���WB�+��"�~s���IM�(e��P����0��GSԇ��mJ\�9�H�#���s��l�4� h{�
���4��>�.������]�NtO�QX)�J�M���|��v�B�
N�e��@�`�iq��1P�>Q�-�Ym��h�~#�l�șL�1Ÿ���1ÿ�U8�MN�kd�	1�����pt�=R�\P�<u�ap��h�NJ=	��b�e�#���ض��7\�붨�Ԭ����cF	6�z ��̨��׬j���яj��\��7�$�s�гA�z�*	��oX��[�K7�2���	@Ø$b<w��:5�~�D���u8��(@����)��]���?�ڨ�$��~y�ź5�Ekw2�kW^�	8a>}|��T�b�g��I��(�rb9C�ߌ$�U�w��$Q!|YU�|+��\�!-��I�b�g��������)R�d2>���җ5�k��P/v��?	�0�psp"�+�yz�w�|����rپ�$��� �$k)�p������=�\���-���?���2�K{5�Gg.\�6����oΚL�զ����@-���3Q��](���i�6\���eN)���@
7�+5q��M���2l3�S�/0=j���I���7K4�񁝇��cZV���Ӕ���SB>��C�4�6����~e�1��1/�2sB�f؄�p���a|��F���Qb3&t�N���x��N��'��\S��){v.�ϙ�K�&Yu��������(=j��G/c��ɖ��N5��s��;�Dq�Bȴ7����q�?-,
O���_H��\�>�T��v%5���������x��A���,o��ͪ�0���- "�m닑N73���Q���-�D�涌Dke%荒9�D$a�k����2��i�/:r�?�H{'%�в�w��#�
,$l��n����0�Zљ�^6ʘȚLEݙv�!.��p�*�MJ6zw��ӕ
*=�K�3���\���n���1���
���%�gd� � K�Pd��� ��Ǌm����U��Z��~fݬ(Fd��2�E �������@ҷ/3�9�8�"\s��s���rq�rd�m�R:���� B�?LNGF_�B�(��;&$�. N�	������I�����1�d�Z �EgFw�o�^1�Hd��'�M����(���@sI@�t=4�H�q��;��>�Q�ԮL�1��h�G6I9Z6�ܱF�r8�F����]�H�ظ��������j�9�����
��pB��I;���#w[�ɂ����Md́�(� �,T�����_[Po �@;���hMrN�y���#�Q[�گfl�t�l��n(���m��i��,���0��R�_$���A빂�9�U�F�����/1a�O����9Sc���}EBWk�a���$'Gj��8��>4Yrq�ވlDl���v0
����U��w��X�>K�ϳC���/{����D�V�d?3�3Hi�#��wX�%V��ΈH%I)��NM�z����VRϦ��s��I5IOI;����: �1���d��<[�B}�{U��fOn)�5�ZT+qm�;��EיD��:<��H��E��-r�o�.;��f�h�0Y6�Wķ��$:��`�:t��d��@�ˢD�`�Z�"˜�_��H?q鬫�e:�~�|'G��w�mz�o��s.�>F6�V��B�,�҆�h�p9%���筹Ҥ�%�rs���K�zs�[�Ye����V��.�'
�Y�8ǆUdC�vʑ�����i7[�z��Ѿ��� �& 
4oנs�`%���6?DEv�����$O��N>Cjo1�Cu/�PF���yS�X��1��yb,ۻէ����N�j�|�|����Tcf6��rmj��;(��Rq޴JD��/�2��@S�]V��|x$�Y��*�������d��6�:%��������c[��<"��/��3XɊ�:��&4Ƌrk y�����M��#�Na��"V�D]���C��%U�o����IN�aE��@���qR�.HgF����w�V���ަڧmaWv����?|�9f��zZ�M�hj盿���~}Y��S>���kJWI���8�k{�Y��|��,�k�E͗�za_#��=� ��$�(��_��e(�:f�y~,�)��)��v4X��� ��l{�����lE��_�m2N�Q��c_^".�N>��	�K��u�z���{�Րs,��f�L�YM��Y3u��G}
ˋ$~VM
]E�=�6],�:I&۹��8f`4u;*�<-��h�U�� ��>�~q́�׹���5Y{�W[n���Ik�L�6/�J͝ZD�/�n��V{�Y��O��2܃e٤����@��0��;�p<��c�3��P�m����Yk|(`�8�~lq�?vҦ[H��*e�/�h�X�?�|o�BI7�=��R8�2 ��B|���۟���y����H`�I���{>knOo��#�{���J��*��D�b<Gm�_�%�n�b�?�]�h����a��%ѥ鹂I���k�HM��r���j��\�f����1�\ˌ�+*8�63_l?���&�J�&c���5�U_�f@s[�� �ے��A_���ul3��1�\��
��vA�I�?�$������e=�^G�'��2�2�1�!�>���Z��y�?V>�9͐��;N���W'0���5`3Q9)���1�G��5e��.f@�1�d ��c4�N.ܜc�kk,}4=�}N�v�NqCSM��,~��
�L��W!RR��v]�g#D!�v�/�t��a"���Z�Z_��A �2�0�Ik�㨒�U�fScf��G�Zo��i$��;����<p�uN���|f���x���U�G7|$��v��E��5�lJŭ�7;��4�4�X�-���M򘑬����-�Z ����-����[��(K-�6{�����RzV��*�J�u>	��d�稤���u+KNP�{+�"ǎ����������X�;�M��i:�����V��L�ގ�5�n�q8G������55v���
[0Τ�Z����i��*��eFv�'�;o�G��R���8������3��%=��:��#b�'OpC�f�3��}=�ĻYC��)�s��D������o���4ޯB��;'OП�&�pS
��p@�����#4��R�k�!~��b�#�@��z���~K�)K%߻��V�^�1_Q%�KF@��H̙wk7�D����oe]q�Og[�\ �7�ţn2�8���=+����+BpK]�SڛaL'@�]$W�A\�	�3~i@�]��>�/�ق��~x.�H�ͳ�0��d�I�B�\�מc�N�Ɩ*!K�Q@����D7�kbU��)˃�ݮ�Y���V�xƎCڙ���yl�<�%�^澜ig�S���l�3 ӑwR@�ƭ%����L���m�6���~�YF�;Rg�v"D�,����$�J|'�|�k����Z[��*�,vR�S��s̯�%�����9"K��P>$�c�&�kz���`�HKr8yp���>��gS+y�Ϟ<��(c�	ɜ�Y˘�4��|.��˂xN� �d�_/&Z�	A�h6��R����8��V�f3�����'s��\?�?���^%CE��<R_�,F{���W/H�T��t���������Y.xv	_������.����ޤ9V��) ���I�Я8�
#e
%��+���zz�YRq�p ���k��
F��@� �Ug�+($l
��8{��	��� g�7�km7k�f
Y*?fU��\2v�?<���X�:��?Ի�yt�Gx0�	)����>��ǐG�E���J��\����'nU47@�e �����0���Rl�����ZF_m\��gQ&0���$B8���<T�+]��ۀ*�@��8�zĒ�X'H�'�D��`n;�Yd�8Bb�I�N?L��8zg@,f$�+��]�nsώ��2�뒨9�E̯�I�^��;��x�zD�xIb%�;c}�v�3�b<��^͜�1b��Q�X1L�+ a;]��;�:�~&�8ى���I��$߯��0:���1y�9��U�����7�: �!@bg���}�pE�@1�F}f��t�`!��	�v��n��R���<�'(��fkI'�F�nr���t�(<�雂%+tM�y;2�l������pA�e?4���1���� %٘eK�侊��n��|��@�C2��5"��R�^T�!�P����!�"2���"�H�n���D�R�J&Z��N�i��kw�X��ȕR<7;P됭�OI���5c���å��X=�N-�����m�R�I���n$a�R������q�Y�h���,X>�;���4�hL�9��ƥiN�RN�z�i�~��A�M�����~��D=;%���!y��v
��G]����ĝ�R;�?�A�Z�j�	L�aY���vߴ���8��Mv7�j|�!�̹��o�2<�#kv�D�E�yz��kT�X��@�:(��Zrj7ڻ�������,�9���2WWO"��Ư��͇���Z[�X�FA�<Fj2��N��Y�� ���D_�eİ"*���� zc���ݸ�fzn�n�o~J�kc����zuGl<�=%YϏjoAX0��-��� ��.����ڜ~6x�����);��(C���im$h:j��,W�b�|f�9��󴂧�N��a�r;���+vW@�g���!���I�f���0�қ���/aex�Lf��������Ӥ�f�� �hkwUE"uJ�#c�n�ō>��v`��u}Ľ"#qU�/�&�骘�����.�.Ѕ>Z�R��b��B.�<��N.�P��բ5��Ej5�?�j�p8���i�+Ҏ��o�1?�n�w�b?���YN �+tbB�e >01$.6��3S��Jg����+R�1�i"��U�l�I
.��9u\��ުyr V
[s�!�v�o×���������_��_��]�L�H�A���*#�9PRd����բ
�jT04�ĵg)�.f�Xaώ�j�>m�j�*�=�c�����W�6�HO	����xx)}�N/��-��k ���$z�o�<�
>����0B�Y~�D��q�D��z�RHe�S���Oѽ�;��[�'���:�๹*� ��r�ːn�ِ������9���,d�h��� QPМ��%`�6��z��ȿ¿�!6}U,�U��A������iq���f�� '%�X�D#\Kx���E��\���eX�i�<����j�á�M���� �+����y��,�qI�h&���'	�:��/�<��G��S���CD�z?���pS(s�C���q���s��;��'/�(s���8h&;u�!���k����N#�ӕ �]�fi�t�c z�k�z�^�X��6�h����dݴܦ�ܐ�p�� {&�?[��蒊��q��̵˺���h���K��l7]^o���^w�y÷^�؏ã	�ݡ�*䐂�i�^)�q��- h��;����^]���=y������!l��e��:���R�y��3ų�5��ԫ��H*�+�
��͌h���O�[Q'q�6ש8�U	��
c�B�d]�(^b�:J�+H��#�U�~9��I���a� �l}��UK��$� ر�fF�/ҷ������ϯL���^�fù;��s%]|��M�*F��iĶ��̥K�՛�M��<ic9�_e�։�7C��#�� ��g[J��˳A���G�/��[V&��,��'���o�[Ό�Jy��D��}��{$�oI�UU·�|;s��� k$9a�S��U�]\$_ȘN=ho�*��G}���F�(�9�o6U�]��@��w��Q(��$I�oH�az��u����YH|��Nv��&��:���%�B@W,����s�Њ����z���GP:��k