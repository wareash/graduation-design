��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|�&���ڴzk^�2㨗e�M`Z�_P��xܨGbYe��ɵ���1���i����i�K�?���!ͺ���^k%!'R։F��v^Ҷ+=r�D��ߓ��H��'��p���͋�֯҄�H,���2ӂ�=Qo�5��g���#��{���nS rv@��ArX���-�����҂v���8�n<�C�VT6^z��Otn\MLؖ���;BT*��96���.�g;�����,GI�P5,�f{p��u��:/P~��`�j�'��< �o��O��
��4Ц�����ܭ8�1@Rh+��&�9�첍�܁�f0:{���2Takb�l~������޸Ya>D.�O�PP�DO��Nbj�{��֘N�ss}|���`��p��P 5�_�+m#�	OY����4u�ī^"pJ"�X4��ί�3�4UE��G�nPz@�1�����[�`��T��^�������Iy�j+}�𧧨v�͏+�ʕ3�nq���FSQ
J�g���+�[#�����ɗ!1��u�+����q�o�V/��m��i�Ԛ=y��Vq#
��(|���X��-U�&��hH�8���HJ�pt�_�ti���H|5u,���ȴ�,���:��\�^`���_Z�x���bML��;��*0��XB7��o8SJ�
ՙ�bo�u^Ҝv��n$T�� 9Mc.���|����?�s�-~��W��!����{aI	�ˊ�s^.:_�k�FD�>-��=e՜q$��e�U@Zr�{�������cֿ�ݟ��h�nB����t��X��8r�c�f�_��h�@@jf�vйLV�t�� �٢#:�M!U�%���2�!lʃ���9����'��)<I=ţ����9�ȕ}���5��Wk��"��Y 2'�k�&5b�Q�~\bf���p�.X�^�� |S�R���l.�<*�V%���S��!�7R�U�v}��F��T�{��a�yL���C�^���+ӳ��"��8�8A� �֔��>@K��Iô(�R'�F��;��|Ag��-�\��c�|C 4vU��}�r����X�k`\bx�F"\���T}�Y����� �H�6�W~3� �?,��[��`�I�Ƙ�@�-s�����b:�����I���O��n�767m:zL^�گdҤ����iJ�A����V=��>fw)��E��}��7��A3��o>:����MU;G�1��/�Й�>�`�&I�jac�ǚOa�ʂ�-r����~�J}b�a�K�Z��)-��}jr�o�A�����X5���K<a�	�-ް�0)���(��,N'[r���rp7�h�b�@)8`k��0��S�#��1%�g>{v�%�YE�F<tk���� �WB�o��=W<pS�)��%�Ց�`(lTt��(􁴳g,a����8��ӳT4IXn4qȫK@�1�Q~�a��i&K5�2|�L�^�r�ʠ��ǽgnx]�`r����>}�<��zP��=-����u�x|���Ą
imI��|�/R��y�12�l&&}�d$Ϝ�?��'��G)n���q��^�nZh�`����I1����X�����\m��rU̆^���+�qV�Nr���h�J��~,+��D;2�C8�����CT������C�� �ƚzH���S�5ʮ�⬠X��?x�U�a�ͫ[Q��	p;��"��ܝ6����2%g�?|�)��x�����3�0N��\ԃ����j�&,8��65��xs�(
0'�����&�$R��p*��p����wwi�G�M�e�>;ދ''��vy���Ы���q�ٽ@�����:ȱ�>/td�<�w��lv���	�oߩ��9�kr�
�`�
 �0��{�1@"��ɨFEr��`����M���B{2Q�B���Y㜍R΢��y:�J��p�V1��W�ڋ�D���`Iant�u~�\- {�~k̚W����¡YSǫ�l����y&jLHM�� M��D^�{L?�+Y\`���@�F�� ?�V����}?>e/P�O��-"n�� g�����I����Y6X��n�5j���f�0D=��}Jz�;�U}P�[Q?=��z3�o�N��p�*�K�#�� a���vr�$���i�##%� ��<�f3��(ă�F��/�22�G�,�B)�i9<�:�M�in�I(v�}I;>L�d�q�}Xx�O-	�bB�,l8�$q���\���;��!���d�4�Z^�6����D)���>6��Y] c�� ָ�[�_:��=<�a�)��į���ƽ�������T��!t��v�d�b���	ݬ]<%nF#j�d�l@����.5�����x"��<x�8Ja��E	�������>�H�A	�ӝ��=N^����Ji>������r��E ��<���6h!� �����;"���f_+9A�-	{�'�|g sT�_Ic�m��!�.b��rM�G׏.�Ί��6=�5q�Aӣ:��$bE~`�6[���F�b��Z�@��	J�*��QdˁO�c���?���1�5����^�+Uӟd�k�t�CO$taJ�d��bA��T�G*SW˿x�>����;!%&�{�����e@*��[���//Q��Fy�I���U��1�r�G����Đ_H(r�����Dg{�N��\P���<@4�.(���'�ՊU����h?7�C7(�������)�hZ���뫆稅� [DKf#~�>곎:�
�j?ǂ��b���m�S�e�>}=��%GV��ݯ_H�{��4�S��r0���Ӣ��c\��5�B�'�q�J0���#T�kƕ�)�$�I�zx�qy&rz{*����������_mj�*�䄠}!$�&�	L��������R�z��NIuƹ�mN:��ۧjI�I|��H�hJ|k�-���A���v|�!��K��ȱ)�\4�Ⱦ��(�tre�C�2����d��`������Ӏ�D�B釯B05J�=�j�����o$�U��h����HT)�]U����o�ft�����3�����ɔ�bd�V�F6"�ʥ�ye7��w���C��_$jxע`�~-ӃVCf ��v���׮ݏ����$,�ՒG��J��Wn'O�b3VvD�_�	d��`.Kg�4~��UJޥL5|��ye T�FE�@��KЙ(�4|���$���+ڍuj�q�w��B��t�����v]�=ű���h-�g�}�� +BL1��U���X��5�]�|n��e��yU29}�ۮ����8�DJI�b�nnJ�,	$>���2�)��w��6���Ofe�Zw��3�.z���K��-Xꅾ4���v��=�2f�����o�'�X1�\�0<z��kcm��>�q]O+��bʜ����e].��wc�3����u�Q��m����qJmӦ�f�J@�HvI�m|?�7�r���*�~4崰���F�:���_�*�k���J�~�%���uA=F#Cu��]75Z��!ͱYY>b�OB�=�n�̦�����O�UD���@�&vl�K=���HK�0?}:=�P���u����Y ,��$��졙ȶ�?=�*�����3��m�ĥ(g!a�C}��6c}����%=�-�I�/��J�J��q�X���������րg�_��ӷ2qC/�Y�IYk��ڠ�b�
kN���;��x1nq1��rt3	"o�8�%mѱ�(n&#��mM�!mGB<��)'LT�>˝��w��t�R�am�|=��YzMWV��#_�7�h����%i�[0f���������M�j@��9���2�����%�� cP�D��GeB��OLj�K�X�b��V�����Q#�����U�11�foR&'=�<o$�|d0����,3ọ�ŕk���:X�]�[�?LR�e�U� ��vo���P��)8*>�5"�(F�[��\d�n��Yk����`�eX��B�"�����:�S�~�w`�� �� /oLV�aa`3��]��T�;	����X��q��2��U�����v8�=���>I��OA����gT�p�"52�f����7=�.�ϖ�)Z�3/�
 2�
��\C|L�O�h;���Mt'�^�0â��֜[oݺ�P,�7����������u�:����R��@DD�U6��:����9�i����~���~��N܌����
$M�����s�S�E�ZÁ6�׼,���!�E���l;�x���d>;�i኱pt�[��3��0���W�&"�`<���.)��=��v�r�_�^>�Ď��,�Lv�=-�h�NY�EpN�-� 5��,2�5�`�1��<Hf�3Y��+�~Kǡ���د>������� �?�@�*)>�@�b�#�98C�.�j��ޯ���=��>��	Q��(�����z�:�l`Y�T�����oo�f܂?���7�oB]�?}��u)%��\���ed�*k?HG-hp$���f'��F�SpM���r$1�m��V�v�ա��z��N)l��G¶������k`x���R�����U�QvP�ܱҴ���C*���:�����4����4 a�8��-)�=�|Fo=��ApAt���&)�j��Ey�ؔfK�c�v}�s������0Hu��~��4���3���1:J�HIwϯn�S ګ�!�����ƴ¸=7'���#���E_I�2��	[�O��1�ėU��� �V�'� o��7��>V�����U>��r��y��iI��3I��ޟ�q���w�ʥ��:�-$��t*Քr̰'���zJ>K�m���j48�ޝ �.|�ރ�P�A�$�Q��Q>��Л���:L�2��\�$�;����W�Ӓ��>��'/�f�IK@�!X=7���LW����T��N<���X��HզB8(v#m��B^�rgvS��@g*����T�]E� ��_�$O�w����~�eԯ�2 z�0x�8����[�@ϳ���3 �/�SY;����kB�ArND��b7�`�K�il��	)ښWW���r�����j�v
V
Y���Vr+bH�mIN� ����~ג����.�T5>cl+��JK�b�2.|�P�w&�#�p�,�*Z��Y|XMc�
���J<�aWc�%��(_aYx��|�/�-n�Ԅ*?Ě�º`.o������S5'�s����iC/~Pj��^�Ŧ9����H��O,�B���:ɟ�`����|#�b.7a	�F�h{}��9�o<4��B�Fy��VA�Y�9��O=��%��t�(�3w/F�u��+� �9D��͑�d��:��?wAj���׾�ys�I���X��$}Z���k�f0R[�Q�=�v��bJ�$�l>�����'	TL�� \-�Jb��u1J����"�v��{j�7�
(�|�KF���K�m~>�kT�˫)��=�`����;��G��zo�n�1�{�@� pG/����X���&���V!���M����GV B�/j<�Jʆҝ3��P�M�ջ_X�+,A�^��x�v-�^r ��c�	���{DŃ*M�Y� �#@3L3�A3����.P�j#x���� R�?w�c�VE�Rb�L~��soF/_�H�^����Tu(��y)�.�,�]�*@A&���XMmU�U����T��844H@;�V�a��FD��..t�!.����L��a�Y�+´*)�$����q��Gc�M_�&�[f�d���~.��;Z	��E�X�H�-�ܧ	Si;:T�$�c���[�`i#/�w����Kj�p]�8Z���{�^S�ip�)݃�d?? ɑ5�IG鯎���rq��ݗ��.�q�`+2%�����TH�u��Wʓ��Xś%��͍DȢÅ/�dbq�I4go:�R��44�\F��B�f�פۇ>�}J��,�Hg ��,�4:�uX0 r���������e:� u��B�'�Y�DWJr8��WA�Ŏ��Ճ���B�����/���F�nt���m��V�j ����I�Cp��P�a��R�Z(����A��+S"c{^̉�{�*F̈E�`EH���^&��;q�f)>7�oxE�hM��S���>�hE��9����i�s.9��	�ݪ)C���UJD�:;�9��q�|Q��
�q�7+)�Тu4�D���p�N��.�$�q��*��t�ݝ�MY))���n�c�/h%����?#~aؙؼ�	IfFr,1v�N
������{