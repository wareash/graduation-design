��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jåا{�\�u�?߷�dn@6�zf��r������;�O):�l��f_l�yȆ��CM�̗ZJzc����zF�M��/�b�Я��p�����ǣC$]-�b�0�.C�	�+��RJ��ct�M+/���E�KS^��~%����L��w4�ۄ���3�70�B�6��H�+���N~d���a�V��*$�%���:�#�Fw^F{W@l�&�+F��HC�- %�޺U"�8��8>�j}�@�r�?�t��0$ė����ۧ�����ԉ�2���^��f(H�F��֔`�s�s��=���.�(�P�PT�S���2اJ`!��N,/�@Zډ��[���!ȉ����lj���L��&BW�w@������j1.�Ā~�(�M��G�65��1S�G
L�<F�����Ԥ�B�Q�����4+A���̄���C��qÛ�M 2����rX�a[���%�����m��宥���Oi�dX�I�^�C�	z/8���$s8�`�pŕY���U�R�X���e��~��XPX�y���g��&���O~΍z<Q��OU=�Hd�}���ƃ��Uoԍ1]7��[���>T�zA�LO��zKy���q/@��UX�	A~�풙j�NU˯�LА�\N�c�ϩ�a�¶L@b	a�hS�n�K���X�]�ߩ?�WG
�a,TQ�4����ߊ��AA��#W�|�U�ӝ*�����ts��sw74*��\6�hhߕ�怜�#Lh;F*�����~���&I�6:x�� �6�+;l��p&�8M�TG�N/��k�����r70��䷩��%�(�_t���3���xR�t �:��ʏ�G��;%��\�$e�`AҊ��'ө|Zhm��cG�t�����)úd U���C�Z˂I^G&��l�@Gk�G\1Y�� n�DMp���r)9�*�%��==]��E�������f����	P�[�צ�4�
P�)�QE� v��p��V|���+�Ssb�/w�Cx`��.���k�)r��4>�S���V�����5���X\���|��oC<��[_⽷��,<�/`7.)�d'�pGW�6�vw<��b7�>�\�G&X��� m�C�j��S�b/Ǎ�*(h���ؗ�e=:�Ѕ�H����^;L@���c��f=P�Ig�_b�#�~�8���l���ayQ��mӌ��2c4�*YL��0�N���_ItP���A�nm̀�v��v���(��&�C�)'���:(���CIZJV}J2��{l�in(�0	fy���n�*ڭL�&����Q����B�9���.�
�xD��CE"�e)������v�8�I�2ԶQŠo���'�$�^PI�!#2��������];��	��~Q�Kp���o�xЇ�8X�-�D��j&� �4��'�Y�Y�)�7�B���Mb�o��]R��	���n���?=���>���_�7>��K��Ҹ8[�.�۵��9�3gZ�/�[��)���ؔ�Z��PF���Ln5��w�ao߯ϵ��XH3m�O�O_i�9��@+	֌��� �����6��d�ᛡ��}���[S�d���W��̧$�o*��������|�B�}tH/q́;bm����A���t0�)�N��~K���pE4x3� H�c��3(���o�Tڶ��VX�HQ�1����`Bhᇥ�`|о�r�����2���wg��F�f��P�.�$�#�K�kMz���$���>�Nǰ9�z�L��I,�����LZyt��>�D�@R��ra�i���"�un��, �L�zH���p6� ^���V�:0/
_��'"RM&��Ca!�J9���E�f�'܅�"�z�Z�K���J�֔�O�ُ\\�����"G����E.ƭx&���5��7�^7LB�0�Dڷ��Ũ��Q���{;Ge�"���%̸�b~o����[9��<����:��61����ب�VN�<�0F��w-1���3��Gv����-�(oy.%1	�7�^��$3����ĸ00���?)A_g���Jm�,�ӇQ�~���;)C���rk+n�`�Bƌ�23
�V��=Z���]�R)���q�*�¾|o)�9ۛc�u���@�/M��q��<\�.������{� 'O&M��2���1���c�-�ѺB��A�eǷK�*JJՖx�!�W�
2�dG~RϘ���z;�y?��&�뤫o'��'�}�x
u$�&�~�7u��D��J9)�5/�������Sx�����4�
�9�m�k�� �_��*EI���c������Y^���]B�������b�\cEq?,r�ʹ*9OQ9��<\Qw�����}���Wbu���J����uSߑ�H蟸��X}*�����He{�r�0?�T5" �������)N�4��Pi���n��q��Q_���UG��-�ShN]���O�-=J��9�q�z�y��e��2�-c���Ta��Ҡ:���虒�5hϊ��6��WZ�PnGD8E�K�T��ʐ������pر�I��m���^>���$��^H��\��$�G�5c�T�)N��Zb�N7m�!1���OeČ��"����<���{�N�J�҄��������2{«EIp���(\4��¹X�K1綾���s�D`!�����9�n��{1��dG}Ԟ{��#��۶-\�a?���w-hUsƹ��!�BG7'p��m>�7M�|kO���&��5��B0�R�"/ꆆec A��ÛIRN7���vt�v'�G� �C�G+�ؼm�pr3ݬ�	��z�j��zK \�t�tu/���N*/la�h}�wP�s�6�� ����S1`B��Ո;�XOp6b�U�;�T�?����Y�.3�����=>���Q�Ǥ˟pk�pY}�v���6����5�:̇Q��$ ]����K��4c�Lˡw��%��Deh^B��~E����X@<˱�ZѸ^ט�9V�"q�B���+-��G��yj.k6J.&��5�qB<�F�HD�oYa�B8m2Z��t�Ne%فYĮm�u4��^+����ܟh�ĎV/d;0�4�$�{��9��$�
�zE�]�	)�[�I�Rz�-�+���\����~�%���w�ji�{M}��u���ӥ=�{�POT�a���?�r�b�<w��R̽h���n� 0˜��*�9�N���ΟB�ݣA�����{�~ &��=�Y��鯫�ݘR�`:�ZƸ�x�(�b�<ߞ$0�̓I��#�A�[���ޱ.�g�P��M�>�{D���6<[y�	6�o������ڢ��5YEW�7g�'_P;��x(%{����y8���8��
�w���?Z;J��.4	AI"��(`l�i:�r�&Fo"52��v�-���_�9φ
&�u�����L�k\-��R�ڝ�� ��ƨ�������P��6��H��C&
��q�L��VA��{ e)�]��9s��^:�˲�;���d�,�.�;@�Q�K��]�r/�e؍lb��Վ�Sm��������j�P]<��]��l�}�g��n��2>�&��#���	��˰}vph�`���Y��]�2��M5��+YcV��%�Fː��e�Es8Fף̖����P����C�}����B�0` �v�M)����������{�'�/�$|�y�Q	i?��$��v�
|QBae�������s�y�-���T����b*���ͺOv�"l�q���J��K_�aH61�O��CŃ�'u�$�[KW�=���=��1�`7}ru��M����[�Ǉʅ���^ܡ�j2��0ܭ[R�v�h^L�@K$b�]`��E��ˑ�4���`9�N��е�$6N��������Q����"�)���<�B=�����V��:D�T��SEn��O��_��i����ZN7���2���G)CU���N�̫�v`�2�s%���/�!v�9�!Cݫ,�ᕠK���۱## �ͫ2|[��v�F�3��Ug 0of�ԗU������,�������`SȏJ�����4�q��EW�܃�m8w�>� �.��g��_�"�۞:�����{�GgWT`�kg��1k�JE�@/��c�6�xͭ��U��6��}f&��%�7si�S�C>oy3����8'.��tP+&Qr���so�ST���J�{Z4Cm���PƔ�v:��¦�����B�r�����H�(UY�uh��X&ɾKkhd��I�iiv�ƨ��X�����ܿ�l��m ����;{���Z9���@q��f7m�(z';��"$\�u��R�@4��r�
@���"��48�=G�F'�ڼ�S�)�b{�q2��/�>IM��2�قl��S��,p��?/=!DK�7͹|7=Q�$P���l^�k��(z�%���f0v�H��W�<�%�#�<H�M_{�������)���`�Ra�(�����OK$���tOүٸ�9o;�Uם�<�[�	�����Sg��G�2�0�?2}���������D2t�+���r��;�iD�7�<CВT�{�]YW��-_7^y��.�}7�0�$*�\�P)5�*���+	�[V�^`�ə9 1�\_����p#@�qtdE���O?��&:�5��)}+p�X')䳔���)95�n8i����y�o	P����J�׾�^\��m�-ь\Є�÷�k���!��H���_���4�3rd��=b������4ngc6零|��҂y
df