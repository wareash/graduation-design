��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jåا{�\�u�?߷�dn@6�zf��r������;g��Q�u1�K��+�	��
�\�SF_�%��@Rv��(���wrB@`�~B��7g����64�5P�W�6��>�{~�~���Z �7����m.�Q&-58DK��F
�zf	�rRij��^��[?+G6sf��t]>��r$�c��y:M��2��ܧ����;�5�`d�6�,ퟠ;˾��j��u+�Ν�@��b���G���>U�}.����g4EE����:K$��$S(���ZX�S|(}u�כЅU,�
�?��y����`�ji_
	|G=�U8W��>mo730�	�=�@鴻�	&��'�ؐh�ZTB��<����kԐ���aQ�#��awJ�N��@=�鄥���Bj��;cc�v���O;��)f�i�"�ӁI��,|��FS���z�Lj� �:;wl��u����F+;;θ�o�1Et��P�֜�9=������ ��)QH����,̛��v���9�iI�#v���a������>�r��*��z�BO��U�[��;���̕<}5:��З��?���CQ�L]t p�������Xl�*��Lވ����VOFT${n`@�w"�)�B����J[�d����dkm���,#�;D�䥚�|DV���`į��ڿS뭮Z͘/-�?p��m8������EY9f��j���h�Ф3H\D�gݺ A��`� X�*Rx�?A.].�
|���g ��s��`�����<1@��6���&�tO����(n�;	dP���h͛݇��Ar���;N�&/�<��w���7�S���+d����%�.��F�����=1��}O2/�}[��b�1淴W�lxگK^)�p�I|�^~�B%��Y��G���Nb�@�d?Y����x��\HT������ـ]wFC����1tGx�"����(+��z�r��y~Q�
Ⱦ-PC�l�<:�G٣��T�u�U84���A�qɮ��yt�(I�?h*0����T%� &�hCc2���^$d�mpD6��gd��/L�^`�j��q`)����P�T)Ws�R?�=�𭲾�M��a6T�1!~r��Se<7�d2��"?в'�Q&�D��e8�KVJD��R�v�Ob��qkB��c���vUaU��<&k���_3�.>;�V6-�l�7�hc�6�\����@
�Cy��&������l��vƊ��A�ŉ�e�kmj��'uPq
ϱٴGTI�`�թ�](��/h�����Q0v��Rɓ2�8�ůiϢl�Y�\�DU��5�7')����k��B�3�&&�BRkg��X�����Rh�� �O4F��{!'Ņ�Y�kb��#ÏQ�P/��S0>�Ȍy<]�e�ʃ����7��0���Ge�	��쮐L��Gi�.�ؚD�W^�ܿ��QEf��j��dn:������:�MFD<?ܬ�%�j50U-K��<�ʠx�����hZп0�W:���g 3�`�;�-t��hJr�eŸl1��<���n7eP�Kk���*OC�k�f��%��k�Z���#��#(�am��j_�ξr��O���P�",]ҷ�8��;� &�����XBڜ��=rUO�ĵ�L��TX@ 4�u��A��L����u8i+ro�ZŤB�?��O�q��0c�/�xE�o�G��l����POź�B���]�}�4S�测4��
O-�5�p�מG�8����i��h�3^ţ���ݳ:Q�Q�/N�@��yЁ���>��F���ř��3*��_|��7Au�`vmx�0[�4�f$��95����Oi=�.�)�ꬩ�r��d�3���s�S_�>b��_��}����UwQ�� e��zv#��.v2+K��� �@p.-� �<�
Y�4�F���K��^?��2��O�����,�c�}����c�>���Q<�c�L�^�.)l��*ap�B��'��m��/i�)�+���֑&�<��}����PWK��B�[�6&u;������5[8^�6d7��7@����<+��}�Z ����g^OҷqSy�z��Է7�t�E��رV_hZ�ϧ@����d�����@:s���W����iU:1�Kq7ZL����#˅h����$x��$�����	���8Ψ�r���W(�:�M�my\:Jh2���[r��&BMnTT-O����9U�4���f���tz������'>	E�9�'�f����e�7�b&JU��|��f2��,=�!��;�V���:�}4|w�h���+��;.fcmc%e���5�k�_�G£B'=:K��4J3t��/�W[�y�n�3l�1��w�Ū�&3.s��L4ˠ
Kd}��הG���*��I >�����Ӣ���
��g7�5\�P��a��]��n��c=� 衶Qv���)�DR���rv�� �@;��X���sgǮ�E��H���Q>��nBYxh!]��e�jV9����3j�豌3P��(bþ9����S�� �����]G�͹��0�tzU��l9u�H欞�K�Ѭ�4�&mc�R`�F����z����\>)Wp�(�-��� ��t�:x}��f(0g��kݝm�����ҩ�~�?=i�E�f��q���XԶ���I�]K��+��*�uG/7���Z��!��[�w���	���W��NWHV:�/��)��]I��xj�� d�^cQ�}�_�L���Q���7�#/ �S8����ڤ��k�h[���^͗�3>��qR^;P��Y��䦺�����T~gz�qȘ,�ú��� �I��K�`�^�uX;�4�-�(���q�wԛ�Ud�|�X0Z�i@�8����S��}Q<)2��ۚ%��ٜ��l��,��e���üＹ���t��<�b~P�w?����;Ċ�R"�ŭw�6��֗_#�l�`\B��u,5��4����i�XH���J����z{���<�ǹ��b���`$ƧX|�Blp%�mZMϊp#�p��q̞�u���61���g�U�ð4b��[d�2i.�Z�Y}����8�בxH���Q�����!0�^�������o�����m
/���g*����[� 	���l|օ!�a�Ɩg����GL�C6�B^��q�rX�
�Eegd�.�����p�?���϶��Q�m9\%�КE�`�Tމ�,sp��ی֐��2�NԴ(~�3��؝v����23�O�G��k�������pZ[�c,�vEH�d��t۱��Im>Q�2��b���ş�����Mn��U�*sztږۅ`S�7؈
6kE0�M\�3��j�P̃�8��ڼ�l䫮?��*nfV�����>SS���Y؝�����(s�82��wG��a�J�[���|XH5�9�?l�h8�<�V݂țH��˒�����Q�֖��ׇtP��MsXA�ڢ	�����x�`b"�(�P����!�oV"��W6U��(t7*�U}9�D0�Ὓ~V6�r5�^%���w��Zс��Y��[�rZ1�	�c��F��
�$��J����	�t�H"	)db���]D�7��6.����lf'�W�R�*�]�O�jL9n�M�&Jt�e��N:wS�K�3��"���э�CJ e��5��G���8�`���s�7Yl8G����	��>�ټݼ�n>[.uc]���ʍa~�.�rT��_'�Mm�-#��|��W��� h�O eP�4�Y�lu�\I�񾑴D}�*�Y�L=����+��*��W�&�n�;}^���]dM�������,�v�p�U����CF�1(Ĕ
\�[�	��\}��1iI���'w��\�P���[�.3�s�{��SL��t<8z%m,���~�祦���_�����$�n(��;��
���x�̙����[�1kǟw����
[<�)���Кi��p�(�rJ�9�d�,Q7�g��i�*�AG��es�Gy�r���o�!����������+焄�P�-*�ne $���u���.�׹�I���<XéT���%B�F�hs����)dA�i�V_�~�I�s'�����΂d�̵_Zߗ����ʤ&������luT,z��32���Dг�"�꧍��j����ǬS��Nc�j�[{ۥ�Č)�]0����\���u��8eK�Y[9��JD�� �k�q��J�Q�7-	5#���㮩(m�h�}�'����*�<��������G"$���`P��x,,�s�^|
}f���U�Y�C�^�.����� �(޷�n����m2Cz6!7Mp��C#. ɖ�B��̚����2=��� ��z� p}rW�i�ĶV��%i�E���h�N�Nx��5���Z�ݹ��E�a�@rbp�56Up�/�5��pU��[�pq����d�cVHL�e�]E�������g�<�Yi����*�E�+͍�w��5�I%��&b*��~
d���D(m}ۣ���֪����#�AyS��`z���cZ�tSC@E�y�4\�90�jQ�Q��]����]�Q�䉟YF��/H�0b]�8�=�!)ƞΫL���~@�a��Es1eJ��&ȩ �Hb�/�g�����C��ߖ�..E�`�Itьn��k�I�n�/�ݺ;Mm_�m����qS�IB+�L,���V̖�`����L�no���S��K��H�2�l���%W?'�i���lGȕ�Ԓk[�=�uiq����j:
���}�$��-�4���N�>雲�o�)
��rr�D�TN��2��أ��%"e�Y� Η��^��|I; ��5.�J��\�.E�;N*���>�������(�3(�����o�'/�[�P�����h����{�Մ���Z�0<��D"	��[(�E�
h��	�[��$+_	��V��ڪ��&Q�Y���.w$��W1���y��M7ֶ��Ŝwf�'�_6S ��ͽ�m�S_aP:'�n\o6�!��E���E��9�Yd���^�34Uo�����j�23�DfU+��N��
�^�z
���vk݆��
ה�d��� ������$^'�S���~�������!��x$f�V��!T���g���l�<w⳸��6��2�%�������w׵�'#+a�7zԞ�q��P؋�񽒡ϲ|����y?c�E�Tl��?.R��ք[��C{�s�B�r��]�]n*G�����%j3
��2�9g����	h?��p1s"�,���ȓ�aK-��(���G��I薼v8~��)V�ٗ��)1������*�Y�<zstE��NH��|�Y��m�B��܇��c�o�O�H'�j�U!���N�A�/�i�#�Iɮ��c����l{sC�\�N��ɼF29ı�L�baL����
�-	t�jeݙ�������V�GF�q%e�P�l��S��ם���y!����-�g��}�û�2p�����6�͞Z�� �+�KY:��Vgqt ���9~�T;/׌�4�\�%F{�#�?�Y$[	D��
��j�AٴO�qܵ<�m�|`2Hf�2�Z�O����-�[8x�ss���o��4� G�=ou2$O�s�FĊE�$U��R��)���U�C osÙC���Z�(7@�uYp5�ʢ� �ݢ��G�H�1�.)�#���5E/�w�Άt�~z�,��Kd_{O� �%�=��Q��M�_��P
�Y��%��q��3��t�(2��=%�6T`ږ.r|��a߷��'���]�WS����h����g�O.����*GB�9Vj���5�����<�����B��¸���*N��wFD�g�����m���1Ӛ'��"�_1�a[l���Kk��2����Ԩ�G�L�F�4Y�;@+Q�)�S uM�x��njσ4ܖ�)V`��[�5gҼ�y���I���|qd-���>�wY��ʵތ���s&y�]`%�Lo=%�W��v�����!!)s���h�*�2����j��H�܋�~mKv�ZE��N�9B��������8&S�S`e'����_I��Lsr�hP��bd�������+�vy��	O�"�{�.Q��d�(L��������T���&4~��^eW�b���LDcJ���L�ݏF����F���}���>�����<�Fپ��g��<R�,DՋ�R�S�t��\�J���a85�k}  ��U;�%@����-���N�>%,������9��BGd㋘/nQ�EG�&�SZ*>�ѣ�<&��a,Ƥ5��U��p��S�l�?��ǔ��J�Dm��Zѵp1�A��^2u�´f�R�ErV2��Nf��7��_ 'T��/�=��Eo�f����r�9rn):�A�����IR�Ὑf>2�Չ�\�F{����@��,�s(İÅF"8�g(2����f� �u�|rR�=������r�)��DD	��v�^3��ň�:n�K�;W	���� 1!��\p.�{T���ϴ"�̢���f0��	�*���+Ѓ:�@�5cc�$tW����$/(�a�g�����ZG����A^NN�M���ӻ�i�-��~"B����T�&m-&��g@��>D~,���,M��& ;�vJ�Q	���e��� �DpհX�it������~�"#�>�]	L�{\��3	��I~�[�
���i��|���� ��P��O+�㡗���	���W�zc�5����M�H2B��ũ�cYo�8c[�y#p�Z��%��6������s�{���Ҟ���"*��;��٤�E�2�OY�9���Z��H���0�݃`����S��Yqw�qd�9x�h��`�����^~��$�R�%0�'���,Gw�����+��Z~�XT<�4��q�Nc都��-�^�y^�m�^�Q��2���2��Tn��ⶳ��̦�]�l�~�M3#�	pM�#�sF���`0��F�+�g���~��Pa��|�V�z���)�c���꣋,��Z��|��%*��zK��t/�WX� ��R��Й��2����i��&=β�n��>d��ZeX}���r"WX����r	u@����f�� �������t���Ө�n6���5�!e�F���HO�U�����7��w
�� . vR�
$���{kQpb�{�e�T��mW�Ӈ���ց"�)s���\�#ة;GR��s��42�S&l��en� �Ci���GP��"��f�Pf�A�ik��{��!�����G����ٚ���1W3�|�����	�u!��T�_���>�������~1���z���ⴿ��p ҂�����kKX��#���z��w-��(�qP�K��j��W\o6T���A�Z��u��	ɻ����c��L/���vb&��i���B���T���^���Uz��*㇋y�Y=[S	�+b��	�%V�?V���_%�le�����DcUbX������,�ַ���oZ�B�	�'���4�wo0��,�L]�j��h��P]�j6~�f��{lk[�f=�V�1|�J2Q���.�a�	]��h��ud�
l��(f=Z+���quh������&"[1��z���bό���"d܏֨�|�˦,m��f�՚�~�⬜�r��p�'￬�j�9��y1�,�zI$���¸=�tDj�����.���R3H�d9!����ֹ����bv����m�Qҕ�xW���I�^�\
�|�p���_��ܙ�P!^E���:k��T?�"q�^-�I�2;�f��-��N��ӣ�'���h���.-=����E`�����R����ؔ���[��jqU��|}����K�ŒY�!��+	�b�P��V�"E�tg�Qҧ���Xf��.���(E\��#�TQN�1��������7���r���
Pɭ��ʫԄ���SORȪϑ�*8Z<ۃ9�eT�N/�CF����̿�C�fT�,��,m�2���m#��V�۸�Y4�+k^W�j@�D����DW�r��
[5[��V3O}�;$� u���UY�����F�W#}��rbDi.�51ϯ`���p-ޭ�8B��3�ԗ����{"a�a��d�g0G��q��j���.֨���w��i����Sgg7��֊OP��UV�xϯ��>�~��/��a�	����R`~c�N���+�������T]�֑�˒��=�.RI��<-ݥ����H�̱�?T��cZ9WN��3�g��:��A��p��u��d�O�K����4B�W���f��X׌�w��_L|Q��附p��y�����r���$2:g�c��6�)�D���B��{�%>��|�ٷ����%��eD�㨄?S'Q8ůڝ�('��C{����(�`8�w��,I��7���\\d���]֤�'S��/|z��A���,B�.�#��6Ly)+c�LѬখ�\�6�2�:�"����:Gɛ��=8q�A�9��&ޚ��rr�d�����;J7�D��R~��;yb�W��ï���[�ҺdI��=���������K)���l� �f�r�	�z���;#��h������m{n/
�e~W���r6�Ⱦ�.��C��4�ʃ4����a7��
t���ŗ��  ~��DҦ�D���P����w���SX(�=P�d�T���̅$�[#^��E�n�(�����>�|.�)\^[�+��j�R(�V�zx�1����D��V�>"�=sLo�_^���Q�d˺� �}a�;�0~d@f�沛�GyN=B�R�n�䥸<+���j����
D�+�"t��)��1��J�9�y�����@�ŕ�*)�u�YǾ�q_0]�JG$?<7!�Kͪ1�w�S�|��6��ZG%��Ow)��V6��)��~uy�M;�z�o5�m�������K�I�AH�R(���$���D�e����� �%݋�\�,7���n�
�%�rؕ)cb��l4������"g~��n^uū�|ӂOn�t>�7 ���9���=~L]a�Ȇ�
��-��E�^TЪ����&!��iUZ��]ʀ_���6%,����e^�����BqG�`��֯��Z]���CRb\��tvǿ���C�C�1�޹[�
�SQH��ϲJwZDw��E5�M3���N0��{�2�@���j4\���nt�T�-?�2|pɎeX6[��Ð�o~�Q�5a���ğ���n���)��.(jw��wz]"$��ʲ�@q��y�HB�/�-�Ռ�oV�D	K߃BD2�H�w���_�3\D=������$H�d
_ˬ]T��)QY��o�~����S�����T�^�V��q0���䤕@>�]���d~�P��D>�s�x!�`�:{��31�9��:)�	*E}e��£#��Q��۬���Q�J:f��
��ۯ#�*�<<���A���de��<�]�@���=��g�OV�f�^���5�v������v}>sw�O�{!/�k� mO���/�:��z°9�k̦��bW>��iD0fL�URP%�P��xx�@�1�V�e*��1���_k���8fd�����8���$�_�7�xF�z-ҭ��G��Q�7�)Q�ge/mDobF�}Pޑ��V�(���'{�(���([�)Y��N�%(�6�o;�l��k��F�L�cF�}�����.BZ7.#�7�ߔk�~�.�TO�iF��)�3{d2�$����Օ����-�4��cn�����KP��X`�1����֥��\��+��E��˼���,�ǖW	�-�M���Q̋?"��2*��f����< x���8�ԢK�@���ү~���(;Kx��t�N��F͞�M�O��k�n����w� ������^���P[�`���Í�;,����m���%�`aS��$?�K�}�n�����ԫA� ݑ��d���2���y,�1�{�z*NK��Jo�{y�P�A�Sk�ɻ�G{��3<��-�R2x0����V1�W^7FƏ��i`�k���_2X�`�p�|R�r�/֊�K��� ����
"�3���5�C���X�f7���}q�O�X�6:'�������݊*����ڇ�W�<�s0�H׍U?4y;YI�H}<Ggbe�{2S�!Y*#l����n�������:4mk���]��ߖ�u�`��t2����������0���H|���כ��֤*V) ��i�sgH�}C�D��$����F�t|!��@4?c�E�w7����V�ßv����Ï�G���@�c�p֟1�tLa�+$�"�x-�\W3��%*����[4���{�u�j�ݏ��5�[1���vB6��5O�5�
]��^�,��V��1<_¢�0�����{�P�#H9h؉Ke��?[�-�{�;^��W�v_��XӾ؈f��r8�l��66��
Y9�N��D�$iU(vS���W��ˡ/޽I�VS�����pJ=�Vr:0���^�� ��Y�X�(�H_����n|L�k��l�SC���>9ȩrBIH�����N;�J7����,��M�\T�UTj`�y�0��y��7`�'_�h	��eq��#싪B"	$�[>)n �G	s�ὒO���ir*�a�b��9�A���x�Q{����;USٺ��+��%H��1�E��a=Kvb�Q�ٿ`o�BrLFqg���@���g��� -����rƟb�N2�g�S�"�z D��R����B�o7���k�ј6P}S\�(
�4V�Y��X������ζ
��=%�>&Y�q?����*���7cd��-�-̟?4r�">Z(;zf���k��}�6 �w�����տ&B��)��P�Ib�C��$�������߹����k}�@����I�����4����� ���Y�f�K\{�+����m������1\Ѽ�c`=O��R:�,g:(@�V��
��2��UFǐ
�dۇ�4� �~L�/�{M<�b�^�@G�2U}���9'��ާ
^� �(�	�.��S����cf�h5l�];C��S��Gʻh�v���D�DI���?��U�C��J�u��&�z���P�cf`�(zO�"[/���u�|���R� Z�^`���[���QY���
��?�������_ic]^�	�I��9ߪe�=��@��$L��~c
�IQ��Ȭl�v�D)�a��kfn)Ⱥ����S��dv�/�bKE1ۀ�l�3W8 �z��4�4%Q�8yo�z��uAK�@�x>�Al��J�M_����Yn^Äܐ�LH˟��6�@L7Ϋ45��R���I���i�._o&�eMȢr\?�l�\���Ÿ9���r
��=��VS��45U}i����#3l���mze�G�~���S�r�����Xo��i�����]�j�4)����NZM��?�!�)AhDF���`�,�{Pvl�^����iY�� ��Z9<\�0YB�Ի*�]ttAN6Hr6�M�1D��n�tp�����q��	X��;����t��F�׿(�wd�q�U�l2n�i.�t�zq(��"G2�a��*,2g�����^�O(�m��U�MO<���F�p�� �cmr@O��x��)kq>~�!�	TwL�׆q��J�c���剴�n&�4�"�!�(�3���!(���UUJ�+�Pˌn��~����z�ɼHC9�9��"�����Zt�1��ޟ>tq
���Ig�6ro�=5�͆�g��I� fh���ءcxge y��r��0�b0u7��"O��;N0�PݝS}]�����3�V��������mt�)R0=2j���Z�_[l�	��Q5�B+'-0n��g�����c�y�����
xm_�s)�V�N��o�����V�A���Ә���������oe0��[	�M9}���7s�̠�KXM��ɶ\� �t)��$(O��d��ǲ�~e(����#��kmF�ұ���І���LP������x��χlv��_���O�Ҳ�G��=�ҩ}�v������vw�1h}9n �V�ִ�_Ѫ�|_�>缟�b��Ӕ�tz��6 �^�c���Js��ԯJϏ�,��N�,^�"�n{����Ջ�"Bof]!I6�͑>�b�C��r��l��(�v�}�Z���ٞ�8B�d�<.��KA�<�ZU�ȡ�Q�y,V�w }��%�E8�>��F2A$5�66qCt�ݔ�D��yp+�KEx�߆d
��Zܤ����(�?�C�}��g*������5����Rtm���y���UGD����bp'�z]�6 �ZS�(�Ed����>�y�qL��[f� ?n(R,��"���^,�qN���-U�-�v�(O����Z����5=	A��>���}���N������_P�6�8Ij+�?����V�h��W���-}��#���:,��
�nN2�KK^ W	�	S���B�r��S��֜}�Xr}HLߵȎz���DJ����?�z������X�|>NS�ls����=b%�~��xr_ߌ���z���r�5pyV�t�U��Xw�e�$��Ϊʐ�@3^�_&�X����)� 
�.�nF!!���\'g�5/��W�`�ྜྷd��4���G�,ƭ` �疷�4�6{���fbL��%~����;���$�8��e�x2@m&U��T�_kFɾ�-5@���tSG����z�w��"(��Vt�ٻ��"쒷]8�O	vSX���~{0K�k9&����UИ��󄌄b�����%�5	K{<���vT`�1.��u,�X�IL�� �)h��}��h�=J=���~�+
`'SE[���[�x�9jץ�HB��ha�P偿-؎��k��Ց4�|a,��՝ ������
Z�d8 �@�Il ���L*J��M��<9@O��)���S���\9����8���>2Z4φ	��L%�d�/�k��(�J����T�gL�RހrC�����d��k�󋫒:�#���6ᮊ�n�_�R��:x�s��_y�\��g�s�[���d�^pq�@�%MU#^1�n y=zC~��/Pv��{�i�n��S��?#���8���=}��	��:+* Y����m��9'F��� Osr���0}P���މ�C��o��oj��.t��cvd�4r9|��z�	���%-&�IM�e���{����LXM}����H�d�%�wJY���l�*�%�ڙ4�A]wm�J�fu���j���|�"޺3�7���"�2��1/>k�Kg�$�TKo%�Ę��ܘ�OqWsÈ8Q\Nc@����9�������ƃ��.�h΃2�������Fb��e���*�8K\0��[Cm��W)�:����2����/nz�Hx�W|��Ɇ�UP��_3��\��)�����4/[��O6�Zϼ�ݖ|Aڬ"�ֶ:e��]_�Z�(b)���UK�j��t ����S�ggW�;��_�p�gX�~�N����`�1چ~��g-Wp�'��o�ca�'��$B�_d���ao%W��t٩:��%�I�?�Sö��g����[�쁙I��:�"&�D.aA���EPe�4,�{� x/����V����L䎴��i��V���G?I���R�>�)��I(C,ֈ��Fm�p'R�>�k쎨��80��=�a�3ʲ��s��gR��#�}���tt9�,x&��G�����7+B����3�3��@h;Y�=��O~@դ�S`�%�<ZB�E=Ty	
^�Ԩ��3�aZ*"�F��V�T9}<T���^=[���Z��ggK�z�\YMxڿXG���L�����.V<����=�T�-�P�	�0R��{�3��䮲ԗ�*�LͥFAL�p�l���2d�_Z�_�b�'� �b{qP��$]h�<��yj�g�1E���F�X_e��������H��^�� Q��"�˨��h����L~���]&�Ui�g'�m��Y�L�B�-��z��ɪ;�w��i-�Mk�ĸE�[bS�H�rY��D���k.��r�t�e����m���ޘ�nܽg����ݖ���P�gl��Q�⠜x�������k�� �t�hjX���<w��%�IÇz�R�'�3�љ��3jk����t�Y"��I"ȩwc��Ŧ7F�����$�=�-�Q�Z��;2��l- ,���R�f4��+,�&�A���p��U/i��Jό�8q�.����h[�$�ßBs����Ԋ9|�$4	>�բw�J�~�s�t���W*t�9�6HRf׮�8G��3��x����� �+��c��uEX<��T�´U��D��أ�L��E�BJ�(���6"�Ի*���OP��J\�N a��4����p���ܚN�C��S?�;0<h�<j*Yg��}[�#��^�D�#
SLB3�.u� ~�A� 9�� �{]_�m�a8��F�5_�P����ߗA刦��&����}�*"'��m*��P��U�<���f���YMZ��D��=�"�@��E`W��r��2���[�ؔ���zu�|<4�c=��� .�������yZ(� �ĄM��r`߲~NON���Ln����W��:`�D5�v!��=L+L3bl�G�A�I5�םQ,ee��n�m����H_�Q0�MYq �ь�֤��nG�;t�L�ė�?��P,�]��j�J�z�aS���7��?ێD[+���Tߢ�����$�S�
�Sm��M�s閡�ϙ�q��8}�P�Z'��Z��N����BG��c�/?�w��f>�ạ�N>
��7�h�
4����Ry0��K��H�RTV�c�¸ j�����Ae0����2�ZP�6�X�t��os���t���=j|�~b$[�,�RJx�xgQ񳅞A��r�'�7���֐}��]�����i�Q^���n%�R�-�V)���|rE�
�V�7QK��C��/�� 
R.�`)}�@�?큋=L3
�K�

���������A��i�#��}��[���wz��r+��X���S,������!`NF�G�ɦx��ᙪ�y.�,)��Э*��R��`:3s�h�E��^j9�y�ێZ��v��� ���P�a��^���ҵk�l�l��'�A�޺lg��'W�>�n�?-詵{8�4�s��EL|��8��.%��vJ�ƕ��W�D{�}�r�=֝�azh��K��%��p�
�Ly;2�̷x��+���<d�2��N���G����������Xü�>�$�Z����q���KDnE�b|�;ծ��yE	b���$+Y�m5�;�=$qt����&5B�ʇ�2�uH~ң"��o�Q�]s���Le�8Ŝ��|y��Ɏ�	�pE3}����&�Y,v�itJtʔ����0b2ӕ�IyQ���㤻7'����O�}��o.�(��(OGMf��3��-�Xg���|(z��������C�n��w�Z�l�$i&���V���E;'aL	i���/�(���S\Ҏilv��1%)�I�X�P�%�G#�k��&
ԥ�j
+��j]~���P|���z̢Nπ���8,����(ɰ�h;ʪ���T�L�ۑFį!0�5�n��} �?�p���n�VZ8�1��9$�ec�d	�0����� *`��I���G�G��O}VB:\�i�#9x��F���k��[�v	�,nc�9o21N���-��[V~��ڎ�ܑ�_�xo�����x68��L�)"*�P��l�̹�,Z�@J7%\4 uw�!,(�ڲ�?���prN��Jҩ�����Kazus��'j���`<�����l_^�|gz��Iɥ�,h��J��G�d e�Շ���v�5��H�������.�X�s�߾��d���e�w��(�څm��&��	�;с��H�{\oFv��X�3W�'�8_�$����;�2�^����8;N�e��Ԇ!��t��exh��ܐ��xv.�vIu�#)H�"=ռ���^�J��.5}=+x֓���S�#��]��5;�n��y�����	@����[����W�&���X�lAF��Ts�{�u0��A��W[)�X���j�,�!
Wm���K��>N�������e�~�/�ٰ.�ym�	��`�SYW�01�k;ۛ��p��������t���'�k���ι^���z�YW� %��E���0�S�beR� w��,��qe{���@I�qGki�Vi���Zu��gMv�0��|�����|��юG� ���H�Up��^�	A�l��jHcL)҉��A4.Z1��#G����.�������������Z4a͠]����I��</�e��T��:[&[f@��'���\F��$/ey�}P�Z ө}o�:E��,/� ���2%�+��_h�n� ��e^Vٸ��Sp�omy����ں�2���
�[������e�)a��b�y~;64v�/T�t�	h=kd�8�FӜ�i���b�
����%�9%9�=]+<���|�n2�}���C@���Α�ݯ�I0�ӱ�Ž7�'C������)o�)X���u�_=ΜMpo���&�������d6g��L5���Q\���`��V�+?��` �7���&�%z�'g�s�)>���'�8�8
��Zu�kx�hNB�c��\���u!��}� +����pD�z�#���r�UT��k�z}$��~*D��P����ӿ'�|��5c����8;>��=��N9_}ز�����砷�grx^���E�����Mq]I�dބH�A�4�O<k�}!��GP�V��X5���_�؟���t=��y�7���<k���t��l���i����<�����1��.l�����h)v%*"�t�ݔx�4�B����++��k�Qԉ*＆z��J�YNH��΢���x�R���U�1y��2�t����x��Dq�+���Zg���w��5����j��?��=�:v��9P��$L�?l�(|G��!���a��W��ǂ�ҙ ��2��7�L�ǰ�}Uq�(ꝰL�އ,9pL86�"�m0"v��T���)U�:���C������
�H%�)	�o�W^ 7y�KJz���#�IEQ{�=I�X�^Mk����U`�d.���X�L�u~̍��3�(�?��)���j>�zFg�̩e��r�̬"ޗw�-j�W]��vYa >mw��Q�Q{\���1-�%ɴ�8��:_�y?�� �'Ɍ��i����^���s�o_����,={z�����ܝ2����� ���U��Mڛ!r��1���%(B�Y���sM^Os��*n�b}��Ԝ��2����lqg�p?tB��� 3�pǐ�	�}��;�wK�[��J�Y[b>*:	K���'�'�(�P�B�J��iLH���6�4��=���ġLiN����S�CǶ�*{㍮�m4���|�����G-B(;� �r&y
���C����)����Z�7�r>>FH��FJF��ʤ��cØ���u�+C�m�7�TS���h/��)'|v2R/��-��>�AS���HN�pi��-V�L���Q��<��hEksƀ�dK���@I�gYz��$a�ݿ��{H�Y�9�f���5���j@�o?��~�� [����hk���1�%.ӦB�k-��\閿�P_N B�ql�9$��!��>	ُ�B�C�W��Ky[[�Ф*�ڰ�T����T+�[2L2��)� �+�12$�� ���D#��v����zn�՛�X��w/S?����5�W|O��4pp�I�.�$#�w���M��9bU�p:$~���U�aa�Ɲ��
+FRfg����zMzb*�u�+�
�:2x�욅��]<x�9���
=W�y>�{-��.������V�d1@d�S��2e5_-A��;i3�Τ����"��c�H�&ة�;�r�A������v�_C��½M/�_.gʢMy��F�LL��Ҫ4���N�S�N+I�+f{Q#�j�o�����ɗ���w��&�x\��#Rr�ɦ��X��`&A��ӯ��9q�~Nɭ��"�z�,u��� v�<�)���|y-A+�i���i�U,��	�*quqs���$�ہ�'�AU�8�O[���T$@�zZ����I��)1�����ᕳ({EJ�=t��DC���p�m�lr�p��A��Ҥ���������'�WYV~����x�-��(=�Q2��}� �����ce��;�jz�e�$��___ɯ'�%2�����sE�j�]\oHK�🨂^���&	N>l��%�yUlt��h+���hJ�C�����iB�Xȶ2����jQU�skz������0��f0%�����H��b�s��^<,������2e2�&��cUW���n+�� :�H��yM3b�+Iן� ]��^������,81/�}�[�Br��-ܳ���5ЌVa���[���Ժ7UP���9Z�����	ޒ�8M�Q���ŝuAY�G��MB�N���A@��u�3�p�X��xwod:��� �Gb;�m�ydK�T�co�[d5�qó>u�q����y`���:H��{��/����#����NG���(5;�B!"}�xԃs)�ƿ�����	��@�q�shn!�[��6N˽�͝�BybkV�챩F�:9�����lݩ�:��u�DS��]�-���w� ��tWqB�6���"!�BE�w�����U2�B[H�[툽����
�������/������>�(	��4�ϛ����š��u��B.zι0�=���R7�>��u������IY�R���N�z�#��.��`���[^clw�ǲ^�qX��0�Ũ����8��nYZ�0�4�Л�:��-$S��T�u�-ru]<�]z�*�FC�w���y�7)	�j8q��q���2�k��	g�9��L<�p9g�'wuNh>
���,s�o�w�z�0��4��gj����B�A܇�@�a��
]�3X���e\ۓ����e�W_~��(��p�[�$Χ�C�=�і8N�o�2Q!�G�]���L�����ܧ�@���Y����[�ru2��C$)5����,MϠ���`M�<֣v0 �u���_\���SD
Lb͊��tC�Q7:-���x�� s�nה#����>�]������*.^�7?,)g4�!$�-Ե�5�L�[`��YK��)��%��S�\g�� iᬃ��<%L�+?w���J92���7���Ep+t ������`�ta�n�T6ad%�E���
<V��zc�Kag�	�Z�{(�ej��=L��Pzo�Y�@����Pl�}�diD����zo{2�8�${�(N�p�ɻ2�5�KtˁWc7)K��r@�y��v
��A*����Tm��eA���8���D%�`(�a�_��R�(ՙk�9�>�hϲ=�W��:b�Igb窦�[������V*[�f	�2ώQ��Z��=-��T�Ѷ��@=�C��;��i�wp�č��n!��'r+�6�`K���U�q[�ͲY�?�RtԹ���7�O���S����y�����c^!#c/���.<1���0P�[�{#M+jܴ�ר���2j�k,��OɼO�H�?Gw� �?����=��q�ހ����Y���4
b~��!si�@�3�+�c�Z:�L��z��rxV|T/�� �/R�4ND�����WJ�K�+�á=W���f*u�����-	��e,�L����������@����?
ȉ?��|��/��i=�U��٩��h��}b(3)KJ>q��Y&���ha�ۺ�{k��d�V������:֚܏d�EbU ���7��u���o��?'%T3��o�} �&�BFs����} ��)���73UL=��i�pws�6�'��V)4�3��c�l2�mS�RA�6a���0Yo�+�Xګ���ޓ�̥$y]���фo|���
(1J��]#�!�[s>���0~�둽�|�d��������_sH�0�_�q��i("u��"T���i� ��>�����-�vv٭�)�T$��$�z|[���(&�a;��ùHS�f|d��1�Lw�MTR�i��"�ZbJҿ�=`h�%Ed	�(�}޸AZX�B@`s�����N�3�P�gPI�����J,!�Ab��{kj�TRBF�O��=�pوYz:�?�>Qd8
��ؾc8�VS��Ƃ}R �gC��H���d����4-�0iĞs-��:�-Ib� �7 c[q�
R6�Ox����d�.�@&(߉�����Z�VY7$���CG��M�
�LUx���nV�#&yQ�J'�_K��hX�;k�+�V߈��괪hh��:6�W\A��;?��`��]L��� ґ�I��Z��i�!����j���Y��21��1T�@����V%{��8���77��5n���`1reA ��>��<�c��I3;q�(����i�G�Op$�qA����+ 2��m6n�B�@b�_
Hv��_�נ�[	��x>Pf���V�e1ݮ��H~/�!�jlN�H
I�T�Wk���M ���{�H�(��j<��#l_7�'
�kg&�ӡ`����vg;U�Y$�~֞�hw���u�UNh�<��&��/ O2Ԓ�@=�r���U�ZqB�,f� ���͝�|��1�2�jX��1��T?6@���Q}~�A"輍�	h@|K�A|��=c��E2�>�=9A�,�8f�߽�)���}��7�"��2>�dݥ�3��n�Y�+c'����w%���@+��)����E��;�N�i��皽���.�י�\�sY�M�D]��?+�<����[��w�t"����>����Q� ��ZPG��S��N�f�	b4���K�m2��?+��M1� 䣘T��.%`!$.>M��m�k
$�����ϳh���L��2L;0h�s���Hn�� �1�M��E�59�9�8����[=f��q �n��Ey��2U��g��	7�E�}��\��r���\�� ��t�o~�7����H��ha܁�2���7j<:��	���H:��$%O����Ê¿��T1��B|��H� ��]0����G���&��ߘA�0pb�����@�� 3õAd��)U_�+&Lq�?a��.�����]���@�$��F]���Zx��zI�)�!i��ۙ�����Bb�&n���b��ӛܚ׭t�A��$D�j�|7�T6?�RX�r�֯ͽ�j�B�^W�K\y���da�wB�hr>�����������Lt��c��ȷl �3V3`=�i~�.�''���������͆�� �vTMt�?��]0�*���{��˧��c���V6�}@�*��?�f��C6��M�%ꤢ�gԫ<���l�9?�À�8˩r��y��o	n����*ѡu��e������΀2�<k{�es{?[jgM����T��f��~�F��TGq ���K�q�S�ٮOm�I�mmo��.�x�����-qe��\9�nP�2\�B���Ѭa+�Mޫ��)*9J�f>z�Z�{�
����l����̣���q&��k�:��b7�5�Ns).�`f���=2hX��~��8J��Zi��xvF^��v���4��W�A�a�b�P����Xpã6׺���Q����ݚU#ו��B�d���?p(A�n��5"���c^q�w��B��O�zE�6&�$�G����)���)N���J����v����+[FCA�h���(v]�a�q�8�箭0�
�����J�����<p���~N,��~�I�#�٬��@t�A�8���i[��b��aQ��[nl��G*g���h@��A"M�}E��1R����t.�y �y%A��y�h��m-^���zE>`���(-r���A�}�!Q��+݉��7��	��(�Ѵ3g�6���I�ML���X	H�8G
���.�������u�`"~�-q��U�ޏ���:5���w���$+�0N6+{ҶM)��̠�}��bs�E闕2��$��mBl�l��������q��s��^wQw.�?+��yY��Q�}�Ī�Һ�ڈ ��pJgU�$,��_��كH��E_�{Fk���{�<f�Т)c��J�`�|}�'X`N�����V�Y�"���n���	��F��m��|k�ވ��i�����V���{�%"5t.�w�1qNQ�s�Q*���9�\�C~�����������8�y�$�ɻ;C�i�S�7��ߍ(�pN؜	\�n�0��Z�Qj}3.�|&���Oi
�ʮ����-�9Lv�.Rh@c�۞�E=�d�ӊb���Z��"`L!�ƀ�`��ZpIg�5��mV����A��T&�����k��;Kq	�K9�����s�t�e�^�8J����Hf��W˄Y��GQcb��r��y���B��;7�2#7@��a��f��ކf�M�{F��0/��E2ź<�L�ʼ�k�h@N��<7O�sYT�7g���U#W�����e�DJ�9:�"�.��J@�qZ<�a���?_��啶����y��@D���*%�R<�ʩ� _e.���u.;��%u�*�Tކ�i��Z"ɴ/��t���/]�B��d�t����~d���;d2��#�V���L��@h���Ty�|���]u�O�h���bP���iυ<�+��i[�ڐNe�Ms�qD�O�\�BU3�XY�8�4.\�
=E���K��L��N�F�O�g�^���#�b^�9��Q�n���4xN�)2���P�(�l�m�����{�K&���m5-4�ja���u��a��+�����*��Z�:���l��1I�א�@8�n\7�,�l�:�K�ĀZ�F?��`Hej�wͻ��k�����,"���b-�)�2Q��'|�R�ҝv��do��-�]"kZ���j��s�C+靪_;^�ɝ_��w�~5b������ ���p�k뾶��$��xc;P^`���s���L�F��o�-ddj)�:=+�fb=��c2h^@	t�Z'_�Z�� �6�oT�K�Q�u�Ma���؞�#�h�Dry �ډ�ȟF�W��&����J8g����wq2~#�4�Xe�6���UJ�LP�~.I�����ހ���g3?n�;{�Q/n	�G@7�ے~�1}��UE+%se{��X!F��ȍ���'����1�=�R��+Pv!muc.���ck#�=����g�y�3�3�3V�t�ɂQ���iy�C�Ft�FP���e�C�A���J�	6t���dP��"�>�+ԟ�L?�!h�k�.$�������o�lJ��27ߟ�GE�](32Odjg��4,��ei���w�Jᚉ5r�{QUW0J_����4� 3����O�:����	�g�"]뮟PB���<v�9�����@�3j���#'"�)Kw6l�UB�>j�ւ�HK��§@��
�E�`EI���t���%���Y�0\F ��Y�R� �I���H�����O�C�x�^���$PE������0�@9��	S8$��ޝ'�E���9��ے�3�&?>G��!�G���B�_�aruU~1��Z��5B���*W�e��i~.����O�(���V{Z��ߙ�W��ߵ�rs��U��`�τ]�IK�Ow�]+�����"��
0K�Q��<�>�ӌ����+�2�"^��m�}�jI�G��+B��ɥ�V�.��~�t��+�
Zl��8£�G�Ƅ��*]g	��Vw,Y�e=*�<��(���-$nΔ�ڪ+���P�0u�V�Z�0����x�I6��^�,����8g��i�%�m����~DP��E��a[b����s�Ts�U`�A�E����L�;��3!b��/��xG^NLhS�	q�=��1�v:<D��9��E�`���9��m��\5$�_ (���C$����@�ٰu�P"��K~���"���+c�c�<"yX:n�� ��2����iЭ_K�� �}v�K�ؕ�ϟN�S����~O3;�vauR�Kɕ��t��v��ѓ��o�02�6�/^ɔ���6����"^��bIz7�9��n㡵��ӭ�Puz��Xt��4:+�(�%��R�5��2D���-5h�]�_P9���������v�◸ 5�O�̛��p=2�K�= j��c�F�	�p��ܿ�jŔ� <��ЌĎ�m����=�b�񐝬���������;&�z}���#s�Aԣ!.�uN �Z6������#}��������l�Ԫ��np,Ro��J46��fin��q�0οi��i�,���z�y��3�kʹ��FYZ.�Î��6��)5O^��ě-����d��)Y1�/@�*>�b�ޱ��� �Q�!@&�6����rA���s[ތ&����O�/u�]����UB��ĭ�7!`�C�1œ�56�lQ(4��o#�<�ϯH��}�h{�%�WM����{�����Q���8s@A2����~+Q��u[6ɗ��Z��ގ&~��Fu�1�	W���N-~l�<������O j�U�Ҏ:�gB���ſ8�C���z<0��I��2Y��Cw�JX���\f��*'�h!P/�/��?�Tu3\�B�L|�l��o��.��~��"h]������|"�n��̮H�֥Gp��MӖ]����~R�� ��k��5�CߚΆ��0)ꗾ��?��_ �iY(u���[�]�9F�s���h��f=]�CL���Bu7����"l��g�g���qEA֮��NO7q�%o��x(��
 W�'�*�\.aoPz�/JrM��-� �IF�$k�B�Ԍ��7�Ny���%H�ŝ��	�NU��vF&{�:
��C�v���/�����dYB��  +]>��b�ҿ�m',���O?]*S�3Cc^�ǘ��� ���vQxD��5�vz�uP��K�.��U�юF��L�7h9kg���y�cj�I�4i���o|u��ER
�M�}b���g��q
�BU4���/�7r�_u�\{��Q�Ih�&[��������7D��=>7��$9�>�RAyk<�>0%��C�7���r.�4�[�J�o������޶2�go��p�],@�6���	G��]y�ⷭ��aXw����z%'���O
4����=���5�/>�5V�i� ap��Ay�>�����]q^M�f/q���&ֶ�����Kf�݄Cߑ����t�h�"#T�P[\���u_�Sp�(����
����bo̘�
.=h�e��C
,$��j��K�x��#�`�vAJ��YKd�xO^#��H�<��҆�DA�?c�G��]@L%���e/����- =`�,]��\f��<S�R;?G�(�<R�Dq1m�yq�|6��5p�W�8�D��������czFԇ#��=��E�ZӁ���4�!Bt��4k1삃�[�9���m��z	����0@���0�=c�j�L��K�*7����.IWw$��-�J�l��$�J��1���q��&��̤�k����W/��;��c�$��LkH*��HL��H> )��'C6��1�m�	en��=�]�<_MO�z��0���F�ыK'�?�A"�>�$ߝ���T��@�����'S��=��$�8qL�D��YI��'�S�ސ:����T�pu�����W�V_��k�~�b��v� U��� `�F5o�>�"�+z�i*�U�k.����g�z�z1q�e��0qLɡB�z��^���g~�=�84��h�;���@f4c�T��r`��l��p�f5p`�K�m�~8�>ȓ ��E�T}����t8��~�c�ľ;p�j���o�R|��F��a�
a�zI�h��X䄩`�y�F�U�4��t�
<o
߸u�UMC��w��h$��w7���L���"��RmOSe�|�X�Y�}fjg���A 4��kl-?,�f��d���&����Y��=ǅE�}#��M\��w�{?��jK�gӐfI7�#�&X="'ή�n�íIEJ�������р3�ALi�|��|���mH	ks_B��na	I?Q���;;x`�}�WՂ�-�m�Cʊ��Qs�\����H��8o�&�Ć��9����p�[��Afn6d�%t����1}wLs�B�j b6���YR)�C�ö�8|�I|sl��|�hZ�-��O��$�M������$=�@����QN��.�gH��OLY� �ޞ�T�s֒4���P����޺�i����;��L)�U�hye�J�$��ޛz�������lX����s��@+BFu[��2��O�\�Bk� <��ۈ��1M�nMA���H�<�����.}����L�>\����O>j��ü=�&�nAÐ38�|Z�D�Eu��^��;O;H~�v�=�����P9J;Z���p�z�������(iB~"��o��5m�4����y�X���4"��D�_-$a~�le���(�<�`�D�jA�x9�r�r��9?��p�����Ę~6�Tvꣽ�hP�"_ ����qƔ$���*�"pU4B;�%�Ң�N=��iZE� m�qq�]�IϨ[lA�V����x}ܚG�o����I��}��e,�.B��3̓��1=đ$�̣֣5��}d��~@��`���{�H/^<g�#��A�e�U��y��8ź�Ϫ^��������Ni@�������
梑ޤ|�d�K��*(=�m�L=c( �����^"&��F�ecO�*q(,�	��fE�=�O��^�����e����С1I\���M� ͍m��LQxl�i�� zh 5k�u�.��j�'��m�G�ӱ4��aV�"�R�93�#1��>�s1)G�ˣ�x����q���5���uc�>�l�lQ=�A�!z��������(���rr4�KI��1�dI�Pz���t�YH*}\������:'h��1���q�@.G���}׶/�?�I('�&݇
>L��`.��?�)�l��ݏ�9��5~gњ�u���B�����Tiֲw�����2��_&-lTƙ�o)���싖��R���vN���z}�����r���?jsդI��R�~
�΍�L�"I�p~�e\�_K+'�/�O��BPYb%!�b���+(�rP{�Z�4Ea�WB({���?���Բt�}:z�\&���<$�A#I�A�1�����>����]�(N�|js��2銙����@	�.�[:�t�ZG�a�=~�^�D��\)g2��@l-�������W�g�}��N1�W{��g���UBյ�[��H�jqذBy,�H�ON�,�)��-��l��A�r'����И�xQ���M|�!ER+"��tӫ!o_%#E.�G�ħ��EV��/�;�	(��;�~�[����ݬ��#�<\Х��=��@���� �r��󭆣�Ȏ��O+��ky��>���,Ql��E"����D��W����n#���cM4�8_�GF�;o#)��esЬ���[܏�s�g3Rhr_~�1qzVqvev���RT���"��;n�I_�2��\Y,��j}d�^�C���R0�Lƴޙ����2_���hȻ9�����H*�"�Ӕ�Ľ�Z팘~d|�JU�>@-��|��$��B2�,!�rGF�d;U�H���^�Npx��/��'<�S�BE_Y�'|{�VH�ޥg6L�>���!���)���3<��n� �|٩�W�No`��8��ƶϫt	-����,3�܀H����yY^�R�X�|Q�@����ؾ�"=Xj�h��F[r%�x �(���x���t~H_�\M�S�u)�Ui��K`r��]�]8ئ>�@;�YS����-+;��h5���b����e�F���p#�W0Q�-���QM	ߚP͝��Df���s��cv�!$�#Ye�������n���VJ�+fޒ�����J5��f6��*D�|���)�ػQh�F�n	*�N&G�� lV"GI�n5Q����
�괤��2<���!��������ĸ�}��`��L�{�CJ�!�#�hW8�Yw�g���h|���F�*���
멉x�*&�C����g<#�.f��^Ϙ3����qj���S͎��qھ`�O0�<݌�P��OYv���6���t7��=N!�C	b�/�\gլ�Dc/8o�BG���̪�p� �dyj��L/l��t+%0�LV Zfm� \"�dW���Fb>�4��	�K�K�?��:ď����Y�̷�W���5ԓm3b.�(9�S���'���M�-ɫ����:��9/�����k�ˀE>��T�[��a�����~<�pnY/�W����4��������57��Z��$��e��F�	8p��h6R"�q|�YD�$�C5i6��>nw��\���4�\���<����t�Ҡ�St�BA��#|Ww6:�e�ؿ����v�8��P�6/ꊲ3g"�37����'H1��Dx�\���C_T��9@lԽ�/�-ѽ���<���������0��W����{+���H��^���r�q8�б��!
�f����ƫ[�R�SN!DQ�W��b�(F���p�Y>���f�<�=r^���$��SX�/�
�Vv����g��A��f���] �qo�������'+��;���Ml|]�7���*7�� �[�W#��^��Pza���
��\�� *��$�U#����z�.�鬜y?A�	i�D6ry�u�F*���9�;6�*�9Hju��$L�� -��_�xV��!E�Ĥ<�^�|�'��P�Z�#��_�%��o�S�Nf���03�q2���+6�V����vb���	�xL�6)��$��Z��Tbg}J��~��C�|T�LH?w�)�f��+^�������g����h��	��
�uZ؆c3�.�F�d$6��-u5�k���_ȵMe~���j���f�U��wC�s�9D�,�f�v
���C)�vr ��;�ﺡ ���V�����[��\!d������cC6�O�
�^��ҭ�	��d��)e_ t�*�%�$9�������*����.Ǯޯb���+8"_��x֞'��QI��f�'_�����]�A�k�(�L�������K��e![B�}���:w��-���͏_��:�����RAw�t��z1eCN�pg�S�o�G��J:K�V>�;���E�_����$��k�rZ��w�R�� 
r3 ��q4�t�'�F�}`ꨇ��ty>���:�t��1,R�o�ȼ�Ρ��la"!�rD�1�wc�dƪ���UފFH�Ӑ���֫�$����jt��s�"���G��3u���BR���̸r*�>����+)�^*ꖂ�`:z	We�f/{�P_�"����֦� ,4�޲�ګ���C�K�9N\�M�Θn�j�L��Oh�����M!{�廚��R�U�wT�U��Bz�A���5 �gQ�����:��H;$�f_,Tn���N%;K��p�!���.�ןy�����2�'v��60z�u��I왵��&\:�@����W�uD�\|N�(��	���T���x��Ȣ�|���6��2�!w�'��������P��EW:�m��1�s:�蜢��	�� �t���y�T�mӂ������4��6�3Ss���=��" nq���Nh��"�{����\B��?S���	�ؚn�B �a�p�����:�%��T!+W҉0���8�����(�z�e�vـg
�Q�����H��L�*{��Wo�?p��@bq��q��ВK���J�N��r֥H0�|�i�bX $N�G��K�m�G��������*����&�pg���.�Y��[�3nfoLQk��x�uĠp��`�����M}o�o~������chk�`���-2Q0^��d��Z�p�i�w3Q>����U)��%Q�G#TaU�?��p�x���7͵�HM���3_��.�N�N��f��4+��{�a
�(TA��*C�|C�ƿhN)Y�a�L��Df�����
ӽ2,d�?JIbn��o�f[��7����3v9��o��Rz#�Q0v���
T�w�a5��(r��j�D{�L�VW�(-�����6vʭsѓ��f�M�jk�t�'�����Ѷ��9q�ʰd�t2i*�Vy������ig��.��R�Jfx�Pڲ){~sQ���&(�b�Gc�B�A*'�V��_K)fK�z��J�ނ�����'�t��9DK%�`�ìq��c��;O+�٠�N���Y��_�56čܫ7[�U����O�S1F*e�.~�R����Yhu���Ä$T� +9 ���I>�3�O���h���#�)�u�i�,Upp�g�<��f?�!��� ��l��m'L8�"a�����RHY}�C�=Ei:����c���R�)����@�J��c 03�4c����P��3�qkj��j~qam�8X�x̐�g��+�"U�.F�X����X`���I�h���]ч�f��n��[���.u/���H�8����ؽ4w�D[;Ӟ�����@l@����}���e��������ܟ��� }���Lj�J�5z���_g���'��m@b�`��}��B	C��Sפ�,���^��Q�PU?h��8�����re�뉚���L�'01I�n��c�Ҏ/���f�)������Åx� ҧi;�Ʈ�\m	�x	�(V�z�E��cJ*aa����<?�����d�)k���!�U!nl�)4������UvĚ�ג>b~צ���t>w�RYĭ/�E�'��F��?Z` �V��kk�T~��6QLCS7��OAA]��@�C��@�+��!f{W��]$pp����t��D�C�m��n����l�PJK�5��Y!ʸA�>C���ߤ��-�)�q�tV��a�3�h�&��Cdɂ��=m��%ؒ��$��}�X�B=�s�u���:5�]|�F���Q�ᐋ&��P� �*}p�vP���H7��@�Q<j/uQ@��@��@�B�Q�usF��ZW�"gɭ+'!q*�8�JRĞ�J�r��ė�3�-�][JJg�=��Mz*��i[���z����([{���
�^)���3�BX%A�u��ZǛ�3z^�`��'��.�y�g-���6�d��u���]5(�����~���T�>>����lE���}-mՍ�yc}�Ǵ�����{���� R$�@�w��`���Y�{���!��(�g�S�!L�5���=ޮ^0-�?+.�&﹤>����H��&�z)A;�O��C|@�Eү��^mA�W=���;�O/>��Y�i�F��@0��'s���Sn����2�?��
��_�������$��5�W�H&����y�:A�6��H�o8>u�F��y�ϝ����>[��9�r?3[�&��)S��9D�O���.��H�V%�1�tsZ�fS/��d	*�3B;��H�9��Z����|�Fe�Ţirz�VHQv�g�H�����2ɲ!Mi7y)�����R�Hf�C�i��Lmk��
:��Jզ%��˺w��tBS�ȗ_;�Ӫ	���\'�J�e巖π<��M@J����:s������+���Gm'�m\�jS$��$��f6��	�ME���zq�P}��
�;��m(GCq"+��h����@'�61z����x>!�ǣڃ�	$K��A��������Q�e�iV�g?�(�AEv�N=]#����f��۾�� N��{|$��݅��lm��{��Z�eB6�����B��K���u<mZ}�̠�ҟ.Rr�kX�}fu��o�a�~�HU=�gQ�e}�p�(m�9���s �L��_�+a14v��h
I�D�kt�H�خ!���b�����4���e'���"�AkP~��!��$���j
s�C�}�K��R��7[��{�B�]��2��L:�,��|����^����L�Kxj2ʥ�L�WZ<��/�։~��۹�EOm��sY6l� ʃ~Xd�a @K*�����.�	VpG��������Ѿ@�xק�z���F�*�"$�:+ٳc3�L	jcHjd]�w�w����r�,t�x��7�R�F.@጖����V�*���b!�H���eZ��������	�ų�؇8�4�5�:9n��Xg0:�	f��KZ��u���-����K����M����p�
�0M�8���-�L���h�é�m5>ú�"<���N�jY�&���	�k-��&��!��ED�2&J���߄[�	Ib�o�J�Fkl�#u#v�0m���Z���G*��.�"��<>qjJ��\6�g-GL��tϓ����;�A
�vLGsS�	F�"�m]���1d��gG�+$)�0e��J���,�6|!�s��͠��ޔ��
��`�Cmh��]ճyD�K���Nxq ٹ��"g
ֆ�ySAQ?��+������cn�-��x��E�kCJ������+� l.�=]���1D�m:f6��X�1�p	B����L!��p�t�[����'�^n	]W���xY�����-nvyԺt}�`)Ak���{��+�=����EYd��
�ϊ��8���c����vV�=��6:�g��Y�>�&��A�<�T}a�򕆮�TcI����02���ӥ�|� �&�N�4�K�Ǚ^�z&����M�����G�<��!�p��������~­8^���:������YC�`σgF�L�C?��=Pr�#�V�wY����G4E�L���\���+t
�)3E��{ci�P��UG��^/�=�zТ�R�BNw̹Ҵ0��CM�@��J���!?��B<�����"�����Ru�O~�vF�Kh��\
Ȃ��&F�Y]�Ӓ� �˼)�ܱ�Կ�d�)�X��EҶ9�&<S��.;���:���G�5�?]����@�l=����/p=���Z������O���y�,�6�I�,֐�:��6�w��&��3�ǥBS�C�[��� ߀rS;��WZ��!i6i����x��򓒚:5��̘�ٍ	�G?��3���.���T$M�b(�0��-T8�i����;t:Jղ����ÆU��6�����0nm�CJ��?D�5��O�@�4DI�@���0�L��q��*@�m�Kr�%����� md�ݔi��c�A���`�VTFG)P@+�D��jΑ�J��	�Y�h����W&��d��S��q>A]$W&Xו͝0A�$ݝ�J��5G��w½E�"���F�����Q���4��c��h��
-���l8��<���͓:n��%D��[��*�
,�$��V�n?]񟍆���K8�V
n�0ӗ�Bo*R\�\��}��x��8N�at>-�#Ჯ�F5�p�O�1]�E
���z�U֥}t�gM�����ႪG�Ԑ��q9B����^��q"��=��>�I�r�Ꞧ���݂�R�=Kv��M��<��ϰ���.H���`#�&��"Ƞ W|ǌx�5����
X�G����(�s�h�B����y��8��ͼ4��t��g�G&�����g|�a��[3�~�Ωʿ�{��=��qgܪ��G�{Eoa�<;�"�.w��|�An^�'�~��>��j>&6�	))wE��)�9]�&]�YjI�=�q�\ھ��ǌ���g����p���P�m{�Eٓ��R��ލ�;)��Z��:��_��r�SgI�/e�˟����ۛ|�̀�UE#!��h���ˈ"y�Z�����j��mb�G�5�/�P4/P=����_.�����.�7BN܅��&�&gLhh��z��Y�g(��Ч��=�6�X��^<�n��'�L1�k�R�ۯ��.N�h�Dd��/�
J�/�s���B�LL#A(?v���;o<:��!<&��)Wi5U��,�BƱ��]��>����q�] �E��
��+%��G�H�tWθ�G=.sʈ��fM�˿q�рgA�H�ح�:�ڋ?����D��c�&�����Hs�����9��:�1M�XHH�P{��F�1r`wo	��
,�5ӱ_t�����P�m�5`���O(���f�>��
�"n/G����^��o�Q��r+=5-���܇����]���NB��d�c�����e�4�x���*�fX����-�~ܖn�����>M��&�W{K^�Jcg.JCU������
}�p��c%��Ǿv���-��K:1��5iH��������� ��r��9�P�y�l>�Y�����q����遨M���=vI��L.F�
RB
�Bh�h����^M`�!B\ļ�_�w.�,�wf�"��{%_7,��)N`�?D��݂�X7W���.�B�II�]���J�5���p�w�)�����vc��E�	�}���������C�^hl���AP�I���y~����-|���x��y���q �Dx$���}:	��M�^<a���v�ad�\r�[w��AX�8���B�H���i��xz�A�mrƹ���X��඄�œ�v�(�yZ�!j�+�
��[2��V<=/Mf���i�Cy>sh5o����!��c4nI	9�E��j{���U�"�y�5B�P���	,���Q���7�	I;���I���G���&����b�F� _X��$ 
�O|�ٻ�Zy��d����c�Hq�7D��������D��R>�!�ؑ��Y��Ǣ�B���r�ZF��}O�kؠ���v����W�c}���kǖ�Ӟ��t�%���l�����b�^��/g�q�SPju�Jj���/w�H7����u��ov�V
IZ�F�� �{��) ��� �������	�^D����O���8ƖN��,�d!Ad�D���:�F�؟(�9<�+2EId&�xS�Sr'�`x�!b�Ȱů$��o�KJT�ߢ�*����Qq/s۟.�c���{�8=+�A���b,��5�i���bޕ���>ű�B�u�S�x�Ԯ����	�Bv���}���]5}�$Jx�/B*ܛ�e�ɜ !ZI� ��#~-���PP���s$�F�J	�f�S���y�Z4�v� ;1q�_��[�kR�2wSMZd��k�>!p��|���X��6t����ࠅ��������D��>!o��18XTM̿�1�[y��nП��e������5M�D�/�z�5��j"T3�M�ش��^�G�l��\��օ<��<Yx��as��� ͍��N՝BH�	=p"K�J�o�;��k~��U���� >���yh6H� B�_�[on��@��2g�ad�%�,/��2w�<Y@I"����.w��'�a��"{�$GM�/�z���M�,Y`\$���@�{7�� K'Cؽ�P�������8�C�;ޱԶ�o�+��_/uX!髈����Ϥ��e����,a�g���w��G����ؚ5���̭&�	���f�+����DwfR�	�˘�X,��]��V�֨o����UK޹L:��"�$D�v5����[Yaɳ�|H���~F��U$�OG_��>�A?���x����-�e�e��E��]r7;��J�+��}�*&OӦ�2�J_�Ż�q�A��xաe����S�xRX����Ӌ����v��������0�zR�T:��"�N��!�Ȍ��\q�*'�	�(�8�+֡�IG��Xv��ڇ���m�(���i�W�bSdo��s����Q2S�(
!'X'���Y� ���娌�L���#z��KNK��������V�Gɉ  8�X��g�N�Yr�'�ÞU$^s�����Y��#��O����s'�{;�����K:���q��T����{�5��|��Ĳ�j~�go�[�*8�	[d��ϑ}ը	e}��H;%��5��3�g�s��ּV'�N(Π�Ę+�4`==�����bo#�UO[S�J xF2r��1���f��^
JSY�Ji�t�߱��Ew̢�e���cI���k�B^jɩ��b�X�����\��~������C�|U�A�>t`�^5%�9oz/�s�qz�p�"����Ǧ��P�oKr>Qavc��*��T��y�۵�
ٶV�Ȩ��V1H��`�t�>�lj�������,(g��P�:�4��bܖ�{ڦ���D*�ki5�.@��1�����u���,��H|������"�h���u�/��wE�9SQ��j�k��ڧ������3���� ���Us�s�A�Ǯ�8�5�|��P}��	`�=�ve�z��K��/P`W��ţn�!���T��M���e@��H�[�'�g�`w�C��"REjveJ��2H�,�U�Z�;��b�؇�5XHZ��Z-��C|:��� ./A�ǖBm�Z�U��_(3�_=v�쒼Ge�Ks�,�����.���i/� �t���!����Cq�P�ir�]�R�� h�}J�)�k��&	�\۾9͙�$8J�������+��ۈQ�ӨǱ�g��2]�]^��@�I��?��q!���D��UߧF" b21�]�H)����(9�ضHة"l�F�b���ܔ�t �\8�T5צlj�_��\���!���V�U%�e� ���v�������5�-�O���k2���t/��p@	л��"�\d��q�YaSo@O$�24,&8�.6i�K�T3tB��w�XT�� ���X��o�+��'��_Uw,����d��-�o���Nw�`�ScT�̏cf��V�υ\�y(�"I=M�T��;e��iWG�o���O($�>Sp[���M��
z�&���n:���!�Y���< ��FSi���W���J=�U�����];�%W�S3;���]އ������ v�訕I����O�����ϪQ�ª����4\>�<��$Pw+R0Q�4�E�g9�>��@h���D���F���p ��+�9,kO��1�]�7�(O���h�1�TmV�B�μ�-U4�f��f�����y��̎ٞ	���ۙv_�q��E�Y3W<�1��'�`$��mDC��D���{Nq��M8Q��.���F&8���k^�>���>r�G}뺕���8/���p]T%11�	��9Yf����ٗ}�A)*mzx�)YF_X؟pf�X��Z��W���&��>+�5b5o<I����˳��;%����_?�k�LY��Lh��f\�g&�Q:v�n����D��?R��)�=RO�V�Z�J���EƵ}!������Ջs���'���3_�����
B��/��X��O⹲��qU�De��CEv�h��:���υ�Kb��@��X�a{��@ovA�e!�ƗN���A�B���sQe�+x^ƥ5����a� ��=�4��WjI��������˛1 ��^v���-)��g.���=F�-Q��1�R�g�Ӂy�>˽Z~��\���e�>��T�fhr|h�cS�B��&2U�x�-' �lw� c�t�j�0�e�&��?)�l���g��Q@;���w�����I�������}��۝hQ����(J�@l��I�[W������Li�Rt��嬭����p{�����o�cH/B���_�b
v��\�'�Ny��VW����o=�[*\���������5\o���Q�/����� -���Y����RK�����h�s]� �ݏ�RPb�l���-�3���{��,��Z��+r5��R}�*�E��FQ3c���	�iBx_&Wa�>lq���Fdd&��~]�U���L����]����6���M�XO��-��@��5��Ӄ�*ڨ�:V�ʮ�w�Xq�ƍگ_�m��g��+E����c��:�.N��a��d���D5��T�QC��h�S ��p�g3X6����ofU[�>���	�f�c{��4���yO�pP	�>F��s�CZy�腈�g���M�h�5�k^)9����,m�89!�_Y����g��B��iM�Վ���p�`�W����ݞ���[���Z^���{j�����؇�X�Uh�_+cLv>~�D�&5ճxӾ�b�r�»��a�v���JpGy%M8;���Z�����V�}�< $]�6�h�DaP�>u�����JFd���S����M]��8���lC������D��̅?��ݎ&_@4"��3�������"��\�/����!Sf��@3e�G�W}S������<h��w,:���(��a_�y<P1���-�O�<�(
��Gc؎�]�ǀ��,.�w2a)qt�Ԝ����DD˃��r�����3!&��?4�Z+�տ0џ"e^����u�����m��&.BB`rK��($R�����$�Y&��1�0�o�A|+��;d%�Iˣ�~m�`���3֡�մ�pgCs'�B������L�4�?�0���jXZm��6�p	��B�w�q�@���\�ڔ[L,�"���p �CR�+�-�, �L�4��K�w:�[��C�G���~���GW_�i���;��p��1�zųi�w����+iMH��۱�	��c���<ҡV� ��ԭ�[��z��-@N���S��\�I��ᰴ�S��㼔,w�%�}���=*�:�-�Kr�w�X����E��p���@_��5�'��%�Q&D��=�R�)�|���C�� U�~g�2������=��'��|.�����iw��+`�t�	��!��2�������~��V����1�Pٳ�T�e��R3���ş>]W^�%�Aze�w�����y�E���]�$&��Z�v._�͐�j'�5��u,��U>�j�d8y�r�';ɴdWd��	�<�����䍩|2�����;z�ËDdj`��i)��T~��B�RZ���X����Và�"^�y-��YT���B�S`�xZ��TWW�K_�;�`�y��e�ր�:B?@3���Һ��}w�\����j4p�^�#�5��r��7"o�����~�P4�������.@3y�g7@;��>qݴ!���_�A ����`�{Vc�i��h�Z<[����J���H����u�p�Zݜ�Z��#��^�f���%Z��s`���!��TsXP
$�AY<�W�+�B�^�fw �X�.>�UL#)�����0b�\�/(Ӊҿ�#TU�8����U6<���z7��5�,��b{��rטF��Enx�|!k���!K�E��YX����r��j��y5���((O���J��5�e���GxO��NV�J���!�xچyT��}��d0�����F�sy.���u ��w��j�~1i��}�y�n�ߕu)�]�|Z�pN�x�M��>�� w��k��-��X���<�8���U�ocM�|��GUK��*H^`3��7;�����R�[F�F�6ӝ#�6�!:�E{�V��_|�Z�|���ˁ�)�'֨:$�]�&�]&��8�@0�@�_��d�^��K}���z��N���z�nX���'�gM�F'�w��
��Q������m���{8�;,#�Z���̤�L�F��?��J
�h�����ȪL���8h1��XD)=�?A���:�l�c.\�R5��ڢ�l4ڒח�=��k�I!�·J�-�!	����Td�볻�;�s�Mc��2��s�-��)��T���<$��D��A ��9c�F�4�f+fXf]����;�c��b�nK���Rw3۷���x��l�2u0�eW2�tp~��L�)�em�qxBn��D�>zQ[3�4�*BW�����yZ��+����r�XT����ڙ��1���oLod��-.��,?F*
f3�5̡d%�p�}���V8j���D���N������