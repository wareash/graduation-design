��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ��nͳ�R[�ظ�_����Qq���G�]~��\�^�W.Z��ke��X�?�I\�zA@���Y"���a`MBl��$���X���/~%�cg��OU#,��;o�w�F�~�wy�0�Sa��qC�$�_됲��ݗ� ���D��.����v��C��k���<�$J��3��I
����<[�P�}&ʁ_m3�P{�
A���-X'�H4Eml�}-���i���[�f�c�:Z��� �B=\O$�u�ALߜ��
�ױ�,k� ��lb��X�9��	�X��$SH�}Z��z�Qo|l
}�O;;n��x�C
�ZW �q�	����ǚ��ϳ����d�	M�Q�����y	��Ͳ?��Ia��P��HCz0��?'�h������08V�l�	C�1@5+J"��JA'��n�V����QhJQw$��!���/�����]{�&T���#Qm�.\ǜ�� ޒr\�2]����E��!q1n}Fv-�H��.zX��(�2���!�a7#�qd��j����6Q�����G&���k ��ٟ��2�	�:@i��٪��%y���h�lۭF�s�p��D�pg��i,�b|"A��0G�D)��ޛk�Os��,��jo[59Ӡ�}|�r������W���bY�@���h	��?svw�N܁�ʾzax��У)�ϗ�w��Sk��Ʒ����5�G	|Z�&��3��Oԏ*v�&�O�z�ٜʐ:x���ɱo�N_��(��vy;�Q/%�i�Z�������˂�@��r�����7�1O�Op�p��s��Ϫ��ӿ�a9�+$p�I����T�If��[('2׾_����|�P*ƯnC�'xH1��i��,'M�e���ۇ��B%l���L�Hq�ok��0_Y��)`������}�_�NR
a�I�I�>O9We�Epr�d��!��w]$�AvˀXXU>�Qq���"�� zsT�}&�Nȃ�L[F��R����0��.ο�U��A
»$���=�@+�,m*��1#� ��qX$����=�-b�t������tz36�\����I_t�+�a��e��9��� _�ܵJ�ϥ�� �v���F��5��#�6��<x5q1��	xY�S���e3��?���
��������q�e*&�g�=�Q�S�y�.��M�mR������4�T���X	Q/x�`�� ��?-RN�v̅Wȳ{�C���F���D�5��;%�
;�v1d2����mW��������=����H2���:Ʊ����b�"���x��Ǡ3ץ���Y�/�V�����t��T)#�K�<���#0�x��:�o\��*(8Q��m�A��d�<D)=cugRm���>�aI�y��Z�X�����+�9���d�6�Q���Y�t.)v�Cj�SP]�,�����Me���*ROiT�}쏝�1\�t?l1���g�,n�����5S�0��,S�b=�<��z#�f�[�����#�((�x@�k�:<eW��z��$9����ݵ����.�-�ksq���\^���ڿU��y?z\�A̒�4YK�Bf�F�u;�:��v����j�=�3_̬���̬��ϐ��Pɩ�'~Ř(B������YS�W����_#�(�)�4��O�d~��������.�%Ώ� �� u3�pSW����t�*�ed`޹S��9мuRR�t�}p"����[�Y���8fa���Ba���n�%g ����B��d���W-����B�b�*U�'���b�P<�4^��!0�}��z�-��X�'$�K^/Dg���5�aՌ�c�΃��]� �ݔm�:��=)��(9�P��x{(�5DXxq;�����I��*o���k���͌�������ف��Ud�.м
�����u�������a=s��r�5�<��	��ϣ^Ζ� g��x�,��^��n���D�|^ʐ<�z�����Y-lQ"��R ��v�RV^��u{�Q�(@t��z�~�᠊�ک�NC�^�>�s��X��pb:MLS������������Y�1�Կ�d�r�U��2�
��CHv����� V�h�Tdw< �)V�i�Rȡ��i�~^�]#=��х��,0
�\��X�^6�J�˳j��[�}Z���ld��X$T ga��%+��
�YH	�z��ra�}�1��{���b�D9k���DRy�jH	ܗ&��r�jd�9+q�I�o��㞲�1�>��	������+\� �bڰ�[#j�ݷ�a�n�FI�t�7n�������S��"NS���B@��q�{�d5F3�K@�6�i��5��<���T&-����[�kX$Am��H��%y�1�ȷ�)��L�֮eVˠ�̱{>��O~+D�G1�@j�ѪY	�[�C��:�K�	A�͌�qCe�r�_�#v�?o~瀯�����2��/[�߃���$����j��u�����#�۽� '>�%��s�y/�?ԋ�Z'�lu����3�ӄ'̚+T�Y�h�7���H�2�
5��Z�C��(�J?3���""|H����qtU8z�c�s����ش<!y�ۈ���5�g���3z��-k��bG�� ���p�%���3�Ǭ�>�?�>b��1��Th�Tx���ɪiɽ�_��#��нk�lQ|"y��z�ӳQ��!����ρ���	D%z�躥�R3w�7:�&[�U%	azm���T���?���zbK�{�+q5&@�a@��h�Nɍ�<:�9��t����$*�-Tdx���e���	�8���
�Hz?c&D5�D'�LN������>|��n���Ղ�^�#��\P�u��|�O�1\�*��SA�A��~�~��W�o`�vXֱf�� �M֖��M�1ǂ�;��\�:&�RK�V����'��c��Vl���+�_ �"�@~�Uf���DC���{+�l ��k����"� �k�JH��_���P���dS�F%��^~\�J����βpF��I���!�ߜ�	=Ms��M���T���4��:o��p�QW��8i�٧�y%�s5=�!�҄�@����{��j��L��1w�W��!h_o�zZ#﹐Rd����ތ��l�5K�d��/��I�����+t��(s�/�c�ǲ�_�J��gv��#:�RIuqN�2��%�����%��m��Fq����3��e?½��i�7��`���
HJ�-ãu2-9�(�B��	�����I(!^?L��D�aF�	ݞ�r���T��������(ض����<�w+�����K����� "��{����~܄�pS��i�y�����T��0�{�W�1�$v�PV��6����E0���x2w����J}�
 �#-����|��za+�Xb(�[�ί���X�k_uؾ���ꯨ暼�dZf��}��x/��er"-l(	�ꍌ�R��lX��p�s܅�-��y��T�+#CԻ��I]o��t�ߏ��aAҾs�=G�S�Y������0	�:���R�t�	�&>uj^]mZ_w�R��WQ������^9�O���C�E?��{vЊY$v#gL_+�tMF���Z��<���]���ag���m�A��}�bO�k���ȧED� ��� 2�: -Οa�Y�8�\Z3A	f,�d	-?R"f��]���B
BJ��t��q�~�PF෥"g	��%�W&GDA��U������݁;�m��%�>�oW��>�ݣ�7�hR�}����ZҊ	�h]�����G�W3{"��[K ���E��⥇�������[��>S��#޷W Q�ˤ�W;��g#�����4CdX�\��na\�#�9��Q߿*W�2�E���,�	�x���Xj���)��$��H�"2�y��PϏ��Ad��>ʗ<K
P�<,n���1�ut�8�{<�s\gy��X]�pQ]B�(	?;����H����!B8Z
�-���T�g�|X���������>�����fEN1�����Ǚ�f.�TH��9����Bs��V?��!�4ʎ N`p'b�.����Z>��:V�L��hK�z[���*���z�bw�_�4>H�
���ct�"x�Rgu5���p!�� �lE�=܊��"^q�%�8���6�����k{��RJ��[�2�#��xl���BE��u���VI2�#��	{���gb ���'���_A�:"��]t����'W�J�CAXIh5E�q?�yg���h~?�����vs&