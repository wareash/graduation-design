��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e����d���f{��@����S��>���4{��ת�AO�Q{���cR��G��F��Y8W#å�f�E�KF�������o$�Ni��|�t��>�[���06�������c�S��t�N�G_N"u�DMr'{���=9]j�V\�<��T�p�� z(�t��[OY�>�e���FP�}��f��CUe����gg�U�s8�e�?(NA*���~�Jj�\񤿧�EE@\N�J�MAT1>��p͡��3`p�-��d����7��Ş��C예@)JuJS���bZfO0�tV����+��p�`��h9&����gq�4G��Dm�"V�8���MR�z� x�Oz-�P'/�J?��x\���z��ٲ��I������O���>4�rpeՎq6V��-̪J��R���T�Q���/�M+Ăm�N�揇�aR�W��qoA��Zi�`(�W�����$I�Ama36/�4j��@�A���<^�l'�9\V��a�g�7�Pы����oM��k%�e���}�C��޴��m���.W[�b��.,�dRu�)s�&�\n�U9�-|�@;�P
 U�pnC���Nݰl�/������[;�BV$�7zj�_ܱ	����0���n���.��!�|F`=%�}��H��{��:�~>׊T!���B�+�&0�"�>+S���� ��l@�iu��Rqa�3lb�!���!�'�X/�+���Z�*mC�<��+Sǐ�o.�� ����LV��s*'A�߈!�,�gڳO��z91-p_��z��k}�7�SF�v�F�|�4֤��2�W%�؋��h�-N��}�~ ,����2YŁ�?���v�t}�]8W�3Ml׊��D�D��x��#��9�";2�V���g]�%ǋ��
��W�����pa�N�u����s����=c�  
�|�	b�/o�����[��~��p?��dj\\��vS�xL���5z���:��B@���T	�
e2]���F�ំ���k� ČGrC7TҔ�����k+� #�{d<;�N�9��1�+6�p�1!2?~c�z�t�~�
?����GF���N]�qdw^�#6���"O$��/��:��
k�?QN)��x{I\�"�7G/�g�`)�_'��Q3i"�GY%#j��\�u�f�5qy��#�0���n��H�!�*�&�j�u��:z��>�XT���'�F��Cd�޾&���!��B�I�qMXB��r?�}���a��B^t9�V�*�A������6�=y�i�����-ܡA���h�8�z�׮�~DJ
�Q�f$u���Q��`4���y=+��6����o��#�h�^��"���JH�x�rH��φ�ݒ�3Xn���4C��rF8#Bn�XG�}5�w����e,��"�ʁ���hS�D�Jܓ<�"v�G�De+��凰��׫���3]#6�@���\�ZF��QoUqA:Y
�l���9l���o?�E���
���o���$>&������p���?O�f����v���/�����Gv��+�͵:�1jD=k�=�<7���TUDCaPdr������wŉ!_��dA#�u�A����W3d��>,���s�������|T+�"K��PH޷:���yY�AK1rȔ�0WD���*O�&�z�����J���֫O�hc��?j�e��Ӳ�Q�묌�Ь��x|�T�Z�U��+U���dH�ѵ�����T$&c��Ha6�dk֪���5���G����j�6c���ŖEla�(o��APý�3��U�\5k�a��;>ʁv��+(�-��Ģ���V�@����u�и��B)�yvmq����W�RW�y��q����� ��� ��3�N�J�Aw�={ph<�qp��nV�C�ͤX�=��J4��ʎ�/��w��2@!+}�DN~�$��!BL��L(�+Ґ��Ks��]���ƽP������|�a3F`��D�~��A�@�u�e�<LJ���\B�O��(�!����,�Fg��%�1�^�t�ЬҸ����O�<�b�DR�մ��
\�Z�S���~j2�l�ů+Zf(�/����;����8b;��4*��O�ܦϼ^-�U�uMWF`�L�#2� x.1��0W�ھ~�Ci�w�b�\�.�$�,
�8n�}.$���M��ϒ��H��z�4Ƌ�;���l��(4r_ϒ�]� �����_�9����(�	��Չ.��1W��l�d�]D_��4�zͱ�Mͦĸ���-js�yA��R�]!��۞��+��߯�éAuNo�|����%>�`Gy�d(��Vu��'��M�+�Zɴ�p8��7ry����K[Ъ�E�_���RA�h� S�Z�S��`h���S ��[�<n�3��Ȥ����ԽL�b?E���͎�`�K����vz�g�B� �z����rO�t�'i� �bW����cj��EXp��۫�^��ˏO� �_�@�ҩE�TG_w�ǰd��W�����{#��5�Fg��#�F�u��*���=����&^������7��:��ǪdC"4���zjR�1�\E�H4��H����?:�ߑ�^��0+k�|��� �õ����T{!/7%��ڇu�,�KL(����Z�կ�W�	�H�󺅁*��'��~Ĺ8�"lnO�ȅ�-�Q�d�]O����F12a� >8J��X�P�bF�l
m��]�2���ޱ�{w٤G�:(�Jvd�E�Z�����ߜJy0�Hkۦ涓��P�f�;��}:�& ՄF$$��tk��۩�a��̐����[V��?�ң��6�����"�ANj�Ha���_	�Ȧ�2!�j9��le$�WO?�!ӫ��	 �W�R'�",��s�V����j_4���>�Ce�O��x�ñ���Y����ӫRj��s#"�Se��[����T�^����*l�	/)����v����$�-����Ч{�Wԃ����xŧ�u��ű#t��d^��bz7�oX��[�Kܡ("����e����m�*�}O5#��
T�x
�V#Qn=�ۢ:{����W�>
��6P�3�$�WBxtH�d��I�j���'�[�<�Հ)�sz��8��])~��cѬRā\#|�vG΁߹NI_9C}I��kN��2�A���+��iK���5�躷�;�/�������R1��Pp/cȠ��zGg]B :cI}�4�A�f��B=��+'�Z"x��q�ᐚi&��!]i�A���X��QV�ۍ+7�%���m��Qb��ϊ�aV��DziYD2uu�3���R�fLp�!޷m6r`P�72{�U')�⍰��X���G����W�n A ���5
I�_=��)�}Sr��6VM�Xr��{3v�V�\�ɀMJ�*9���یl���zI�V���4�J���t�|�&�I������xC`D0�਩�g�?{������� �������?��^��n��ؿ��b95\��������f�$�ϺoaS��D\�3������ʺ��ǽ괟~Ȟ LIm��������6^O�@?N��;O(�{Jt�P�ꇰ&�����Y�������N�9�1��[kz@/`����%���Z�`���IK9YPDX���If俁%�ǁ�".�����?�8�l� !c�.x���cC5l�M���ј'V,b���M��ˢo�"-2�HT�1ɔM�Z�>۹����Gim��ܴXq�eKy����κ���#4/�uSČ�m�O���]�Ux��P\��x����g��t[8�h�������.�ƈ4o�7�cRt1Jq{d�2��]MLX���s��+����U�2),�^�������b;mK�`J���1P������E��@��@�/`���8��@B���}�u�A����K�+�*��2����$����;��n�BN�/�ěW�I_��*d{tWr*(�^�!��g��^$�]�6|1	M�3��r�uk��_��rx\���o�-���|BE�W�H@�U�E��G�m}:`q·[�~���G/���9�
A
P������61��%�q7�g
��vИ�{-Uc%q���L�p�$��P�ǵ���G�B���F2I����A�Ow� O��8��5��o_	`0�F3.>�(�; �R�����'�\ya����*��Z�K_�<�^\�G��N:�t|e1�3��H�d���n�Ѡi�ʞ���8��+}����>��䚦Q?O �	��}��aj�qht�g�
~JC�^Ɔ�"��D-k�� ��j��X	���k�hs��y���܌�2��� �-1�y'��N����`�kN<�Qӏ�87��I(����e
ѝ
�,P3������*c��� O��nC�+��E�j�6BD��,��� � �`������� ��}��/����g�v���*�$�}hב���;!�O��[e���<Lx%t~�kV���G�|�g/�o�CN�$F���DWl�ry������Q�W���U���jL����#���$,!I0������>���-3�4��LVe�5�f�-x]��̑���B�:��6��&���]�M�o���:��	�3�/>ч�5U���"VE�E�iu���׽;޺�§�fl;��c�D��S�����T��v$1f%.8�'��š�h���j#x�~�$��:j��c5-g����Q�k�ābs_�w: ��(�Q�Afi���FE�U��捗���|��q{��l�c�2��i�ɻxP[ń�J��o�"��R��9$#�+�蘲,��H���P!�h�%	Ig�,c�b�v��w$�b���I���cjJ���:Z:�R��ͮJ[�f4���#q���,�0�����ӈZ�$C6r��w�L�����I"�6�ِ���'V�}V�։!y�Am �� �����Hu_h�`����G�J0�������&�VL�N�DD�D�O��CH?���gK��}���l��D�����%��g5cZ�@E
��і�j�&ϫ���J Ca��D�9}�߳�Vʋ����V����$#Z�h/���d��b�J�Ψ���4�!���LT;��� ����B�B�U$�q�9q'��g��1��FmW�s�ϭa��H�U�*9��@��"��ZnX?��\�֤��8�m��-�%��D�"}�7 ǿH��4u?���l">����5��a�2g�_Q�Jͳ��׾ �Ȍ�R��J��B�S�������1W�sv�!��ۨͶ��Z-�QJ%���H_H��eǲ5zej��P��ːr �%>}�6�Z˰&0h��N����޹9K��tR���J���-3JG2��p�*��9�녻E���^<{Т��-u�� �	��;M�l�!�d�C*D�Xjq��e��Y@-�0�\D6���x	��9Pf=Ao.Lu)��~ﭚ��0)�5K���H��bik2<P�ԚF����d���^)�ۀ
�(�8^Q fw�u	�1��]%�O�~�&t�w�@��n6(m�S��Ə�ç�����[ƴ�%V&P���'#+��N����|w�"7?IF��I� Ry"�:����m��]2�B��b8�;�.i��z�:����$3�q���2� mF�嫁�!W��eT�n'B΄.�Č�L��e�S���Z)c"�+ۻ�H#�7�VNo'h"a<?��t�;������(k>wy��W��U�fM���M�W���"�sk����1[O��W�)��6F�`���c�.�J؏J�����.���qF�93�Le��_?�y3�Sގ��C�%Ff}(Z�1�i����K�g.Q��Gߩ�#�K*�+n!�4����P�\�ߠ��}eL��0Bm*��Z��i,x�uG{���
z1|���Z`4�)��5i$^D�.��s�p�6����$�����|J�R�D��\C+A�w��̟��Z���������@���5|���2O���Y0�t��q��j-_�b�(���];�/e8[?qT��a~�W���S�'B�����5KMfn�iƞ�F�(�cI�����iU�/����{q�'=u�8U|�Y$kS9�W)㢎	$o�v���n7��Z�=T�<�1'��&'�l�fi��>?�pz'�J)3A&_Cˢ�3~��CW��CM�X��}I��C�v��ha
߲h��]���P��N��1�T�.��^�ɼG��{��.'%����8�^�%�i�ɠ�{HtM�i�.��k��=ϧ�#�����Y�H>���8�5��w�Pf��1(���"�K�_E;�À�������������!�iIհ؜���p��UT�*@�� ����U���\#�"r��[� �wm�ϝ��x�A/}��`L7��4/\�M�'�{���fZx�l�0Bិ�Dy[���hJ�0!��[����\d�i��D��ZS���&�Ǚ�sH�z�-2F�y@���f@_��>�p�)5�����A*�(s/d�~|�:��ُD3-m������ؙ��+	<>��CH�/C2?"���������J,,ۃ	L�ھ!E�D��c�%�"��ɋ�&o�T�<D
1��2�L��U��;�3/�������A�t���<�97z��U����	 �Uԙ�k��Z�6i�i�nۡ�Pq�����S��X���|�=Z�;	�L�vپ�9�`�k���H�9��;5x���`����ÄX�K	+�a5���r�o^�`F�+����2t~���T<2�8љZ���֕�ӓ�i�X�]I��8�)���t�ݵ����l����#F#���Y����m㷰Yj�N"l"L��܅���Ң�s�������	K��n�ݽ���v|�G n�ez���@�BW+J���|�x��@�P?�K�F/��FK���7ʍ45l|Ŗ_�����ٶZ�?&�(@Ԩ
���@�Wj?��+�w�j5
�fkt@>2ȦrOe��v�TTF�E����������V}����l�A	7o�h�;I��3��΅�r��:tيr'"�X9j������،���n�?��̼������ZDa:��`��Ƃi�0N��0F~��o�:���@����i#��`_��D�r]��K���>���$��4wI ,o )�2R�z�e��mଟ`�\0z���m���0���J���,,T4��H���9I$��TB:���W6*��D�����˔�4��A�� ����7]T�Yt���c���7���ήҞ0�B[�&��J�`C�^��F�6�h�Mc�����y��#�s%UTw�Í]�}W�r˺r�g�I�:�������/�h,�si��
QE`��~T�3�Π�ωt�C�ʧ;t���Y��3*�b�!~����x�����VC�Ä��A	��p�	CY��+�޵����?�ť��U hwe�� R��b��<p����A'�0׊Ti- ���z�Ed�kXl��͘ϛEG�r1z������(R���My9!��#>���� �Y*�rQ�cFD���*�ԭ���0�q?-V���	�Uw��� �@ub##a��B��@�]2�%v�9����s/���G|��hnЅ~�^w] �ZX�G��Jюj�����nM�~�M+���?����l_J��Y��dRύ� WV&�ҟ��(3���
�s� E�}��ʊ������j� �X��Oi�,����0'�j�����=����R'Z쉚��Lr�Ԛʕ���aK�c����$�/c�� �k��@%z�����+�UG�r��l�`NJd4�l��wQϷm�!Մ[yd���^|B��\�˕�/������D���?�fn�!,�X�9��b���\�X���793Pm�ݞz���E3� �Y8�Y��kn�v#���V3�j�'����м�^`i*v��N֦8:�k�'��>�)�'���R��;>3;M+P� 	�8�����ī�s�C���R���3q��\ ���sD�}�X�wA.���,�sϳ�e��rxQ��U0�f
�4M��@���p }�{�.8�d��0x�M�J 4�C1.�1p9�c_��}oܕ�ؤzpkO������F��	 �WȾ�{A?@�蕷�dF����w\���G=!P�����ה�몊��ԕg��d'g�<���6)h�$�$�7qf0}.���ʹV��fK=9����w �� �hE�Q�����Yи��;���}���EYź8S�0�y�,F��^���g��A>�&������6r������:A��6�l�,�ʭ�O���Mā����"��7��kbmLRA�/��+�9��V�����7�Z�Cf�R�i�_�:��_F��䯛f�~0��p�$������ّj+��m9��8m���<)l�;fz�._p�����(`�={�wa?�X� ����'�Ot@�,���9+8-�NS�$9K]�uݤ�6�e5��̟��YW,�-9%Z�ӡ��-�;���6e�J�5,���?��/!N�4�O��	����A�ҷT�D�K����``�Q���Xx�o{<6��~�����G���G��;5��4�Ė�9�i~i���e����v�ew�\7�C:���z�����F	���)��d"mR����v�^�~C /a�ʩ�ҕ��3��*iK7l��O�zBw4%��ع�nĠp׿�X���PIa����0�ݐ�®��e��	��.)b��pr��dG�	�=T��t�z?�Q���|c�7d8Bc���=A����xJ��V��:&���ۃ:�!߹
2	T5�5�72�������W��׀�-���%.�0�9�����Y#�|��fk�y���[ص�An�YJ��V}�&<[sbIA�KW&=/��O��Ƴ@�"!���=Ōʛ�
T�܌��!"����aB��d�N�ԧ?uc��#t{�"�xX�UuY�]J��o�8��	�{�5ZQd=;~����g,un<p�Qj3�v���IF�s���W�Z�cY�W:�Hm�Od���h}�kLZu"��4\:I��G߈��;IW����2Uz {�����mk����Ӳ_�������o�]���c�ޮ��i�Ӿ�SՕ'j��h�]�z�~/�8#���] �D�����K��G���y�ɴ�����y ^Cw�/�X.��d�~����<wTwYNtM�&��E�_ڄ0t���n���޹@�u��0#kzM� M��gnD��-N���gE$cO}��@_B 6��GӺ��A�������kT��p �����dv�Y@Ou��� άS�>��V]i�!�WzY���?��'C�w�J��h�B�uw���1p�\h�3D���I>�]��&�mx���!E#d~ڱl];�ɠ҇B]~��`..VQj0!�a�d�Q� T��g=���H��]=�4���Br!���:O$(�&��7�|�v'n�.x������Yw+Yw�S�DP�������ߖh6������A��_C,\�b�w�qt?� u�,H�!g�Q���\�]��L��d�>8�`�QH���A���F��ݢ�dt
�`I��S�O�ɡ��u}gϽkd1�3��O�5J@q��.��|���#S.؎4���٦�?�"�1k,jd۪2-%��z �t�E7@��W`�S��O��q&���e��n1�C,/u$m'�.�Nʧ��a��9�����Pk�$�����(���"I�u�p�D�n2��5�ΦR/�V��;RFWgk,�藽�v��^�)÷/���[���)p�[���)����~� �I'�t�$�&A�m��(�rR/yI��ƛ��O,d���E�݅������P�Q�v�9�4�U�֝ )@��i��T�d�t�5��C��ֆJn8���_�7� ���)�>,����T--��}�&��˱���\zD��%e �q����D`r�s��!������<��I�I��������p&g8��-]�&b~�{,� �L���.W��~��j�7��"����F�7������Ϧ(�?�a�c�����U��8�'��U������~���������{o�짇��UL��ϳ�,�#�h�����FcM�(z�5H�B�v�>Mʛ��nWWi����-.�0���U~	#fJ��Y
�w�RI��Zl�!�^�}�G�k���h o?�Rau/V�[���-���ne�C��4N�o\����|�x3��tݜ�	��a���m�0���~X�&�(G[�r�c+9_x�Fo��`��N`��eZV`]�`����$+ɲ��
�� B,yy�aLO�QsA��ش�z8�K��Ph{S��6�?0poGη�y^
�`�/�m���0/�	6�=Q!�</�7Ea��Iݐ�wr�0S�~6�t�}07��o�u[h�C6S����<`L5$v�x�s�r�L��P��k]�0<ݑ{_�h(S\�:dBa���qV	҉@���g��|bI�$��H�t�]61>,ݰ�5`��-'FtvA7�#��zQ�w�z���T��Ɔ٨� �8p���Y��PT��غ$�(�?�f�Vԍ����^z,��%h��}۝�e2v*���_l����V<h����\��.9B����]���|"z]�*6���j�(�:'�Ӂ�`Rc���!+B&W_���;��� ��D�/R[���
D��{��5��Z��f|�9�y���}�86����ҌJ�S���*�/����ṪK)�ѽ�����x<�Gx�]��n�KS�f���`�c6��|���C�#J5k>Dt���T�A�c�$���� ��$@��!���� ��	2�UbP�>�`��:BzkOP#�~��+�������:m�y2��~/�\�s��GG��kZA�=�c-V�g�C�����?y��Os�5���NQ&�]}?Rx����&R�T����vH|7��!��v -�<:���e�	�h� U��}WqP �tji�<���UΟi�kM!S�<�-��?�+�v5������.���S��@������P�lC��i�8��y�F��z��u�����/\�z�%J�k���i�)��1�ۓ�w�CNF�Y+��5�f_��o̞7���{�D���z`�ːc¿i��HχA�Qn�m�<���'�j����C`^5QC]�+0ل�k�惛��+��������
�H����.C�Fe�LW�S8�|�#}�nA�����H?\��u4���2a�Hkw�3�پTDD�Z�aK��h�����])y	�.�Q"�t�����oc� �V��%xG��g'2�ʌBI@�"�n�HZ��*%��fd6�����f.;*�o��хfY�Y��W4��P���a�:� ��Z)N�pW�2�2�Yl�}~�2���>}^S�!8�.B�FO����ݪr�B��<�9��{5O!s��k�N�,��P�+�����g�m�-\��Q��B�O|�=]Z$�%:L���u�Ҷ-gcݐ)
�M��B�E>���
6#_�H���&i*YD=R�r�-W=����&����h��BW|�����e< 3��['1�q*�����I��Dv3������lb?v@�:�r�쥛�>.�*���k�����5R�b9*k�m(�D�-�7F��ŏ� ��S^=��<B��]K��Ǥ����sC<�,9�lH<�N�cgF	t1���SZ�G��'�n�wI������A]�����d�YN|7�yV��A����'����jj1�Y�y�.QZr��c�[z�V�$iR0��JB��S�~t��+a���&$�ZX������T����S$� ��N7��qF *�jTe�/�zL}"+Ǡ��x��_��2y�!���
�;B���o5�B�zRuჄ�>��?�n�ԻJe��/��4��NҚ�*��|
|m����u�n��I��p	/s�G���K�Y�MQ��1���\ȴ���Vkn9�xr�V��L��h[j���� wW��.O̩���کh� Zm��>��NJ;A8��Nڼ'w�9O�}|T܁֮�����c�rt�wnG�_�i�����A�Z��8���k0z���~�C�vP�K��tK&�P��zS1Vh��� z�+�x`�������S�����U�L��1HT�?:�$�ٰ	<�q� ݍ�B �ĻΊa�x��q%����R~MRY�aŊ�Oix�=��4�fvZ~����2�Bǉ���q��>+�c`\�!���������
I�Dw�x��1�ۭ6 �~�i)�-'��!>���Di$��%V��l<�5������K�n�o�l6j"Nx�_C,?M���=yP�d��M��_*�'�n�!�_�ի��eR8�����A�X ���'d�#*%�@�J���|�U1�#�ȓ��ī	��0���O�05�S�J�=�Ԕ�2��z��E�V6qh0|s.\p�t�����(�z^zA���H ���8&.�oep���NBA�祢8y�Xt
�Ck�+�ZTz�F�o���_���9_�%�^�h����z�����*��o7��������O %�ۺ�{z=
��`K��X��K.�E��e�`���w���(R�8�qĒ\��΍���v(����h�I�Hjn��/�G����y{��4jB�rc:X��,7,�=������}�Bp@�B��"�gl���*	4�P�*��*�Ng�@�c������l�UΩ��T�CO��Eð����J�X��`�ne�2g�"�_��Z)��v�4��'�O�$���*}�(3w,�qG�|�Wa��6�VD�Π�U�#�5)c��ir�F	fؓ�>�i*��S	,��E'���nz�R[�D��YڜпJ�4@��Da�Qd�JU^n��!�ΧzpV|��
U��	�x�*����sNE�66x��*j,���`��Pb�b���#�Y�RMܾtJ�#+:�a5� 9vQ�W�ɩFQ������d�Ż'<V6L���K���~��� �i������w4<Ç�����w ��k�<�n�Az����O�h������q��ݚf�Q�sg��B5�+���"�7��L�ȫ�uULƗEcE�^&���AI�L�T(꨻r���[y�R�$�uh�!�}7ya�
�/pp���h"(����>�6n��zRĵ��� ����� ��aI8����`��y;�1�;�RP3��t�{[͕ �-����0�At,x�%<+N������<L��}[Y�ل��uɠb� ���
�������f!��Y�<�J���NXW4wba�f*����[n��g�K@=�4dd,�Z�D5�Xp�s�;S<�"x�4̝�x��$��=ׅ˕��L�F��}!t~�&NA��K:�fyI�3�]g5V�8�°��Y1q�FGO��x6�yI���J�&cn�-�4oM�KV{(��j���j�*#�o��wC������FR��U'�zl�j��P$�[=�l�����K%�B����l�K\��I?CvVL3��)�6�,ιp	&*zv�(,�I��Omք\�K���+乺��;��ס8 �yK�O�x?�<�~+<�VϩG��BBAG��(ї�Uj�o��ȕ�˿�:t�9Mn ��ͤU#�������(�ްA�T��7����E��<C��2�"��G&ǿS4�y+�.��{yś��3��E�>f4�r���6"M��Q��ڝ�4�~���� ���q�_�g��=6����H0�	�yC�,C����t6<%4*.D�=�[�ԑ��/C����u��jvU}_�x8&3�X��	%��8�8<r_�_��>S����O"���P"�]��/��!O�S�4x2�빦��%�`�&���|s����O"e-!�Id=�5M[�N4.�m!���f��OufTZ����.ݧ<��r�~�rdz�^���`0�_��u
4P��e�nE�/v[����o�lٮ0�P��8Ƈ�r䩄�!x��%yI`�N@�?�}���U�����f#���+E
_��vJ|�	�[�O�/Ar~,�TWL~Q�,�0�L�ˎ)���ѝ���C���*�7�T��Îpv#��L��e�!�Q�҃P�Pb�%Q�.:44w?lW���"��������<�8�J�(j�kJ�vI�LS����nh�dqD��n��៪ˆgo�}
RX9 �)�W�G��7�0��٢G[�^9�\{R!�>}� @�5x�/a�]qH��������ќ��e�������Yj�
7��7L��k �~cI������x�C	C��o2��3�(K��C8���=�qߗ������Srʄ2��33��?���]>�K}Or`�zc爪y4&CBH���h(0��^_�<,$+5"���*/ipl��k0Z��>
X����8�ڲ�(�ܻNҾ�Kňۺ��_Cjhk����$�f<������n�|�q�Aͭ�  ZV���������V=.���Ӳ�0Ϲ������}FK�o�Cn[��ѫ�q]�dXG��"�p���t�x���ד/(;ϑ��.g�ә��\:6���7[P'�4!/�m�la_����/��M�J�6!�����~xaE<�����+��S�m��1���R�D����9�D�|9�p�� �$�=��c��-�<e���M���$��l^�F݀���A�璸���
�9�Li+�x��϶�x�Ѭ�u*���L�-]f#�zT�>ǡs�I�߁���uq{�f�7ߥ���lΑ#)�G����wyyAQ��<ғ��lw���
���Js1c����7�w�������jl�Z��95�%�;Ѡ�>���(%�<� kకT��_a���+�����b1�hI+b^��gB2����pU��G�s[r�k�ߤ���9b^�Uf1�M7�?-��~�.�<VPM�ϳ�r�V.*�b�2#/�=z��c�0��Ⴔu7�kX��� ���B�pפ�ZJ�j�y�h���	s}��'��E&���@�~��y�C��j���CKc���G�Ø�gQ�����$o}bt��f�vr��do=+\+Hb���ĕ�䣚?H���R+n�-׼�}v!Ym (B܇�p���!�҃9@ؠ/[<�f�g��׸�D�#�
U�ŏ7��F�0�<�T�ג:�^�$�������c0zK�
xy�y����(���^��1��*=��\ .̙Մ�Jx��T#ܯ�?�b\�q$pίCÕ	����]���x�����B�\�_�9�(�;�$OD6#�R�d
[�##�H@}�ŎxcU�B�&��1�l�R�sߕ
��ˊ��ԋ�<i~���E���C٫P�$�y�0��h��a��6��z�Q*��$=��O'g#'� j���D�e�R�k����UX[�ҋ<|q��g"\J�8%�`���Q݇ ���)�� 0�Q�q
+���b.�{a(%��N�(]�%ρ��>��~�[Y��x���}������`u51"�Ťf3Nؿ~A$q,��M�')ֳ粪|$|ը�d�?d펡�9�"��ũք��߶d�[����<��R��GǧhF�R�gb������9���]�M�[X��L�KqJƜ��qrdܔ{Y�v%xͱ �EF���o��2��7t�V��/� 7�H	���a2��F����A�"�|�����75��w���I���yu��,�p�ru�.������9�ci9�Gt���3�Hc�M$�p����߄w�����Q���5zO	�=�=ݸ��^GO����Qp �p�#�'������WN���)��Q�e@���\�����w-AJ71�Qo	�瑉yr{y�!}��y%�����������#� |4Qs�D�u�ƌ=,�[r�)'q&��x�x���s���kr���/G��$��k[$ľ��>ۈ��%GŃ����{DQbC<I2R/�qk9���}z>م0���:���d�mO)x����0{����-n�m��f����O������)p��/��B�����g���%%g������qQf[첰�Z#��[������Ǹ+��ԋ�G�N����S���*����g'������uW[U0�e�.��x9���M3���?WCU�md=>��e)�h4L<�K������q.j=�Ʀ�j;4Q�7�o�D�2e3�����j�Z��a�rL��e����Y�����{?%��T��^�y��8�*Ù��gA�߽{a��xb���!*�ǜp<��#n���,8�~R20x�f�)�C�YG�	�׳�Y���T��4��i˥�� (~\
,��.W��q>x ����
{PחTm��GQ#rT>hv��H	�����S?�
�Jj�_'6�v���Gwݵ8��o1�"`�Б!��8XC�փ�5���n����	�P&�r��	�;�26P�-)yByN�7Q~R� y��{�7MF���9K��`ʇ䍦BjẺ���VX4��u�i;��i߻�>�X�6^Y�����-����{��a����?b�g=@$�΋b9��<�`tT���B%�EE�f�o��Җ��/���ЂC �0 �|'S^�h�QQ/�6�>���'=��/��@�jz:�hZ�q�zhdE��o1����A�G3�U
_έ'L;� [h#�T�ޔc9m���ɂ|�3��4���K�ߝ�<F{��}p<[3sVY׫������b��A2������Gv�8C�w�슩7w$6K�J+��r�-\�w�5l}� �A<5| t��g+��'#�3���r*�މ���*���^����L��F��&'�e���ӫ����ݼ�lk���#�K�ٴ!tnf��C !9����b�b�Z����%�bu�Z�����P�����c�o�*�+ւh�S9�Ck�q��I��8O-}�J�f������(�~em8�8~�/�����W�`���v
-�U?�?�mO�/�8r�a��#"�*���	y�eR��A��h�a;��I2��a#��&"W�x���Z(�Nui�|@J�F6:@���AQ���6��#�$;/�C)�����΂��n�����&�I��t�ɤl���B��<Qd 3Zt��o��6s��L h	\o���I���3h}t2�ݹ�^"!����B��Ҏ��~^��Z��[��}@/�<�b ��{��R�>#Y�B}��tUb"��u������e�������@���u�2�H
,�pA�����R�/]�,����i
�U����|w�E�7��ݦ�L�H�	ڶq|���p�Nz�`NL�������>� Sp#�X�AZ��� naB��rO�Ax���ԠM�t�e�S�]p>r�o�KC����0�[iZl����-ֲ	����ޤP:��p��Bګ-f���({|t�E�+�hT�^i��X�ӻQ�I�m$�x�����$2��ȕ~�Iϣ!�i�ȍ���z3��M�������1V����J_�H������!2����ɾ��uvo�[p��^��D&�|�Ð�y����� ��%_�� ��e���>�_&�K��?���c���f��(�V�Q =s�H�v�	��R#�i/�m��hg
d�J�Q\���"zz��4B_�0�Xm��CҺ��/)��X�|ȗ���F�H_~L�܇������Q։nA��^���G�=�[�Y�̇y�P>�V���G�����#Н�9�
�A�mѢ������>)�����&�GO��*4ʱ
y�N#�S���8�p��_����ޣ�a��.'T������Ln���!��V+bY	=��&�2�ƻ�҂���)B-���������|t��P�lA��x��m0W��[M��>�ܖ �<2hK��_�e���4�0W}�kof��p5�ȗe�\o�B`�Sn�Z�J�w%�O�T��3=bXtC{r��$�M*�vA9�����W����a�q�H�~�A�>JС�<�X�F�X�)($!���8��/c �3*�עL3[+		+����-7��q�v|��}��yJ��ʢ��^�7y��u+"�La��/;���͆�e�"=mb+�����u�P�٬��GQ�K�ف���,�G�٧3N�t��[a_��ǝ��oT���D�'=��c���Y�Z�.��E�<O��{���6���-��I^,�}N�W1$K
OeO`%�35t�����	*R\���O��p��>j{��
Y�F>����T��z�g"����yϺ	%o0h0@w��Dq�A��������\��\X˳V��ϐ�s�Y�{`��.^�l�Frb�T�P~�ePuj=�#u3�ݫ	�O�w���N�^���zJB�6 ���x{i~N�r�(�r���`�GL���4�����	c*f���m&Rg��5���Ag��Mϕ�&�E۽Լ�I� �tE!m Α�iՈ�<��8��ÏV��\��Pl� �4c��0���M,/��.\FS�6P2J���̏{m�s&Xh�� �=�$;cу5��tY�fc�_�X��o����ӿ��Yu�D��J�z�Vq���>�su�R8>�uKt/Kg�l�ɶ�⿋$�"MB}�A_�m�l�=dy(Q�>X���$8��\�ʦ�#+&�~��ꑮo9��~R���(QJb^��%�~z�}\�^]��=�Y�7`2h?d�Đ���~�~$�#��NM�24�w]0�b��hs	���M����0�D��t�ܙf�@AC�s��Vr{�bl��qZ�D=��fY�r��{���՟ �����.�ݏ�V�ep<I�QF�