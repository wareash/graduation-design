��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� ��5���5dδ���KdXyݕ�2�j����B�}��AlU=w��m�C�}�S�[U ���c��6��u�������K���ֵZ$�<���?�ޒO 	��ȿk�Ƽ�o���n� �����4D�������;����l�{6d�0
�Z�^�^�2�;�D�
�UjR!�1�2>��Lb�`�D�l�W�?��9�J�ס�Y�u�kK$�ɓ�#�NA��Y�o�~8g�!'Q�Qd���1��+j�i��|Dσ:���x4����j���g��6��� n�벙s���c� v�f�GMcˎ�����0���6�R��$́r���E�^vq8g�O�jl\	��ч9ݢ���/�p-Zo;i�c�at��zb��M�պ@
�G{���CM��0Gm��w3���Q��ɛr�v�^7�<��cq��Z{ۙ��]l���gw��Eh��v|ۻ��&�xN�I��X�eъ�_�PB ��'%xRWh���e}��w��X�ə*J�Q7�j+#�1Q"���E/n3L�r�~��(>�,^�"O <r�b�?��cN2}�8��[�sA����+k2��\�8�YҐ	��~��@�D@�|��u	T�IU���|L��Ms���<��ˊ��U��F�5КkvП=5Ǩ���-�a���ow���I�@нr���\��.C��JxNV��IO�,�{�F�\��kR�[$t�c[��ܘ:^�� ߐ5��nV��m�H�p�m�:��y!o�k*y��P����P��U
���܂��BQ���,�O�/a������2B��1�f��oĜe7�拙���{� &���"�G1����E0Ja�>��񻺼�\�z�aA�=a��2Oq��VG��6�H���c�1��`^��uKr��Q�p�Fj>�ZJ.�~�:�4F�eV7�^�q��M���td_����a����Ji��՟�����	��ZXD�`:�Z��>��6�z�H9�ώ�.��M���[�R_qL<U�t����i�gIo����b�x�g�����8��7X�|4��R��c�t?2
��t��D�r�=��`� �]m��p���.8������K����DQ�Vz������!#�B��"�y���I;�j�$v��+KY�T�KFt=Q����z�#����_[1m���U�+��*��ȗ�?���뤳�ݭV�����A���%1a�HW�`�C�s	P��`���VDp�,E�@�.R����m^0���_�|��&��k�E�0e������l3����F�~��BiF]Q<7��|q��TO��6�!�~�B-
Q9�}!]�;>�g�چ�����^��Uń�S�_|�Ќ�'x=��G܈!|�	��}��y�+�M0�i)���,8�4I�SR_=��$��:i�)j=�yMB(�c�u�gs֘EE��2*��JP���&�{h���EL֒^��%'XI���M�vM�#�yu:\���
w�a�+��k���P��[v���,�t���x�Uʆ���������Q�����+�PZ�A�������k����3r��a��@��"|���`'�v���*ɈE�m󐑟�g���A+�/ZpF����y�$�œ.D�]�i����,	KO����Z� �!B.��hg}�Vp�@�fX�D�t�㛦y�mY�\>��h������$���ߏN�%�X >p�R���o�
�_#���h����A��z�y촦�%��+\��O�,gօ]/P9~ALs�;�@秵�PEZ�u���#�F�u��| ��5Y�X�>�Px"��#q�$/�.�;`=�Jxa�ln�i���x��B@����m�eIJ�J��L(�ۜ:9�7^�es��� 	�?�����j���(k,ER7І8l#��{�h�ve�d�����l#.���]��Ñ��=a$���<҆��1��Ű0�eM�5.��tU�鱻Vk���S���[K��k��[�Yc 3�:�5�a��ыZ�4CPL��
����rh �$�ɴ�յ�R|�ɗF���4�:IUS�_
�oQ��t�-Rc���ͧ�U��j�כG"6Y�V�)'\�Qx�a`��u)篏�G����&G�0��xM�J�3s���X]�k����LY���w]�l���30�(}9rYd�u�8 �[�t�|�:���w�>�27����d{�h������U�5���NX�cd,�;'JK��ZS�vĵ��M�v'��"Y�\x���I���(����Ю�8��Z���~	����ii
�!�96�xx�#\��]����O/ q�U�y��ӿ�EM&WL��D���s7����M�(����Z@�P���uΚ�S���U��
Þ��%/V�����5��W�:����)\A�q�۴���;z4{�c��I-���Hm�8W���[�s^�fT�3J�������*�8�[��XyO]3�x�W��@�[�j�꣱��Io���5$�gBp/y]�uIG�p�9�\���o����vE�9� _?�*=��� cG����Qo|���J�]`R�T���a��z���
U�\��ĥ����E?�d��m�W�}�$���+Q:\$�	������氡���5$&p��hC/��U����H
�,D����9���A\ T'*k�(Lp3{w' �.� �#����<�t��q��2�͌$=�����ln�^{�+����#~��r�b�#��հ����)�U��yQqT��?��y1"m^M�
&e�fu�?�Xֲ��"�˘��h�̬�ad�B��jG�gqn'�W�%�m[�x�c*�vRW཰Qi�X��� ��;�i<w�b��!c�X������~z��Z�_'Z�����0|��w`u!���)v����"U��OKS�}̍�t���pH��``��fg��&˔LĂ�i��J�&��Or�r�������.�<�+c'��Qo�k���٥�(7�y�޹����bܑq5���Ͱ���Z��M�Z��M/��x�	Č֕��z`(�i[�i���R�-���