��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e����d���f{��@����S��>���4{��ת�AO�Q{���=���n�P_i:}g�ջNy9�<���*Q�k�~� ���"�Ncd��0cǢY3�F&�{$�~������^}��{�*�D*���g+���au�wZC���y�B7��N��w�YP"qʢ"�u��Ҵⶥ����$Ԅ�������Ur( �K��G�SϬG�/)�5�.>{�7:�֎c�����<���D�F��Vv6{�-���&2�@�&^U�)ʂ)�=:M�:���=���y��u�:��y:�{h�d!OYF��q���e*~ň��%�sD�V
�7Q�q��)��_�θ�*��|ڜ�]��->Vm��N5~�Z�.���i-������x5���2$m�%���3ȝֱ%�mf9�$����* ����=�4ñM��}?��`�s�9�Q����XԪU2�ޠ�[.aCT���٠[����)U�0�gR�# ݖ�|+���=W��f�j)aﳫ�j� ƈ�ߚ/h��cIey��F;�� P�zS�vh���1�8�33nGy��ǁudf�GQ�Om�Y��q���d+�<�C?�p_a�l�0�/36�b�kR��*��r[�F��I�g����Lt�
B��E�s(��� *,������0
�h$A���ZX��3ї:A�jDS5Ú)�Y�&��������Ǿ�-m����(I�F�B�����Ii�� ���]�[%[B�b���XO��H(�oA�
'��
Bew�����uN��i�3�	�~2���^���%9q�v���fj�뎉���慑�ڷ�fv�=��B��zv3o��1c��.x�N[�={�H�~]&�ʨ��*\0y1d���'P�y�i���,��h�U����\.u1x���(r��B����"�u�eO�p�<FlT�F�b�.�Y���š��M�Ј��JJ#�|U�?W[sG����2(e�#��v�XU�煬B _k�H�XG��f(�A9L���?;�Tش�R���mt������J�_xOzK��Ã��f;��%|���us\fA���ݼ�TǛ]�]e��(�`�x�y�rGf\/3Y���o�ph^ a�Ebd-��Y��A��hpL�\�d)9����Trzg��__,����ڜ?�*t���kĐw@�a��1UU���aw���R�!��ꔤF�#��e�l�k5��C�qq����5J��MS���%3������������I��.����_}�!�",]�Qs���T�3�*-16L��?��E퇔����ǀ����ȑ{��2�ͼ��i��e��^����2#�d��P0/�Sl��}$쐄�����8�����$���P�P�D�NTM��{H�*%��ny_U�`�{bZ����<Ni��V6H���U.d�3��xLXx#��df�>�_'6���������R\Ѣ��%��ptE*����f�Ǌ�Ӣ���`G�B� >Dhd;�yjV�k�ӥ��������:����f�/�臿��8C �(�<�2X!�eGmt���*�Ǽ�贈dSm: TC�,8x�#��I��2Ȍ����(L'g.�j��JI�a�ҝ�{1��y8�}x�t�g�[B��0���S:�zV�L��s<X�La�0�"���;0���Rp2
Is��O@bQ��~��Ջ�_��2d��Ģ!<M��V�5�΢���t6��M�H�_Ne�&��5׶�0Eq^�>J�q�� .�0$5ނ|�b�k!��"@���Oň+�J�ٳ���hE^Z~BP�IP=�$R􃨿h�\�~�P'�Q��a����Fhhu8~��Rui�Xs��q]��7Y�τ:|���|�+ȋTcmT,0���|d�{�b�Z���WĦ���GhWԕ�v�N3`��!�$8"1�S����O�Q�Q?�4���s��ǚ
�h�gl�|w���dcl29�� )�V8QPv,����j�p�l%d�GM7*��ċB��s��Q�]dڻ�P��2^����jTg���8@0׀L .u��h���ͬ��2�M�rgd�X�$�O�����O���{1���L�{���A��6Z �	q�d�<͎J��=�Ubơ��D?�s3>���X""���ȵ��lD�5�
9�VXj�笊�S��=�;�>�i�VKB}E�Ǻۙ�bx���nPy��a�����X�����O�Bp���*�}�S	��bad����/p:Q�ֆN6gv#������E=)zO�u�'�eTC
� aJ����Q���;
}������/Q��SD��B��Ǩ)!e�˨W/p�ɘ��Fs�)��f�����TL9�ejT�6=%C�tR�K�~82�j�V���+�@�����7k��O�
/Q�ʓ��D��T�k���%P����"8+g�3qz��l�M�6��LKE}{[ump ����u��堃z��~�����:�PUVmG�����#��qz�5���m�(�Vj)�,�I�<�OMm��Q{̒�V�Msw��%a�>���ŷy���QLQX�;��Z�'�O��E� �}JͩAٶbM�h	 �aX[��gF��4�6}�}����Uޘ䠝�E�(b-���;w�=TlC�*�%��0[GX��6�f��n�,�GЋ�uZ�6O���:��\�ɔ�(2����,� �nWM;�Gs��-�p�P��{�Pj&��>2�Ԅ�tU�ˋ9�lg�J��w�����	�� ��KN%ϥ�j�{SK [H��|�y��q��A���х/'jj�?�2E�݅����µ̸�K���l��.=�l�e}�!V�߉��S��}�\.���7��b�Vu��Oc�w�th����f��"���ت�\Y]�"y��MS+=6Gw/$�u3��9��{t�1�I&�V���c�`_��V��\�">���?��^�#vl�MR�ɱ����Y�B	O�;%d�N½�SGށ�EZ���k�����c���̦���}�z�2F$�]e�Hw���=�'i��b/q0-d�Q�d����?��"O@�,�.�5��L)�J7����U^n�̾h����n^mE�I�t��#h-TWc�����`b�y�� �G
RW���;P�yCF�VJ�_� xJx�N7����1E�5�6�� пv'�E�}�
��p�����h#D�-��G�������<�ރˎ�Z=���G\z�_�؉
T�[�CxI,���7�����r�AN��at͚x>�c��&&����o��?�ݾ��Ҵ�r���Hl���F�<s+�V�­l>�/�hHL�y��;?���Kb�F�l�OA�|�ˮ�}���K���t�����G`�IB�Ma`F�?�u�3U�hㆤ��:m�T؆��/�3?<�ؽ����'��u�P�Ї���KǞw���*����L`�y�֎x�%�E�qҴ�-�c��vq�֪�/d��^7��V�`�J�M��Lus/�N���Y�9�~^�>C�t��!Vό�N[�ƲЅMu���ĩ"�.��c? �1�q�َ�|�3gwe���$`�R-��.��"-x��AKPb�Rf��-�{R�DYt�\�X��R�`��>_���0���u?�]���j"
,4ex�H���|�a�8C
},|����'s����Z�&�>�����A܀="LM^Z�T؄
�&Y��P�5�~��y�Ϡ݄�i���x؍�W���0
�n{?�۟���~��C? ;!}���%F-1�NX���˿ 2a2m�AK|2r-��}�YR9ʊ�kM�o������䮜����A;�"����`0@��-�Ś�Rd�C@[_��N��I����|R{Cq�:�i�9����3W�=P6���jOY3ǋ�?�m.-��)��T�m�- ��nF����Yo:�ݱm�`����>egU�M�n��q	���l}�!���[��oj[*�/����m>����P�����z�c.T��+�i�,����}�r�2"B~�Mv�2^jp��ԡ�G!Χg#kX�+}�s�/�M4'�����k�O�	�̴E0(��V^Ӆ@�W}�(�hM��P�Z"��[��!
|r��{�K��!dce���$�{g���۳�y+�dN?o�7M�SՍ*N7����K6*�JM�Sڧ�)�u��[�־����̴q#z��Q��3���٨Ƚ�f�xu������/�EZ,�C�\�ވme+::��c�,lz�6����5��6��ID���e��_l�ӝ�Be��+�?*B���Z�D��y���pg�ѪW/�p�a�x�	P�:;�q��m�(�5	��>iFF�ګ_~��6pS[9�?k���]�~�����u��e�
dz�0�B�A�沚�_�}"nh^������z�}7���Q�>ҧ��zȜ_:Vą/�	9o������des�oQ[����%�����ˡUKe��'10HQE���u�0׷:�	6��.SBR0����g�y?Azmk��`�aR�|��A�<��x�������1�|�vJpMY�#p促BF�.�m��;ِ<�)u�y��,l����2p}���c��1kV1���S]� �V����ҳ��j�W�����[f}{��i�0��m7ב�����~��Z�>�䯁&Wo�T�Uޝ�`� C�5[����+�N���0�N�[�6c5����^SIP�?	W4̩-�<�h�)�A�ǙK�=�c����,�[�d�6��w`��� 10�]r�ɪ�/;�"P~𙨣�g_�Id��Fǧ�o���˹�p���ul,a�H��w9o�Dl
���':ݸ���Oj�ץ;z�I��rE���{@�J� � � 6
���:ep�YY��b�F�G��P�Ě��Mm3�����'���w��ժ���X���r����FUAC�y�E8�iN)0����^cS�Q�r�#���ƵY�������#å�`���X�"��磯�fuf��>F&�Ǫ�.�N���K-�ݨ<;��$��|��VVE�"��Rq��|1�l�{�a�<��F~%0� �ЙK.�A�M�[���M�<�]��)Eti��9�J#Y�E$#���L��d	�RBR�@|h3H �zf�����4����< |E���ʙ	����� .a-���&�����վ�Yz�"��α���~F/����P<M�������X����+���A;�!�W�^+��+_�nhc�JD���r"�*b6�p���D%jUھl�K�wv,L�v��
)e_�`�/�1dd,�<�s�-Jq��X�U�$ڇ.�R�ܴ�Z`��#o~���BS�z�B�՛��������1��	 �i;1Y�D���o�Oܒ��q{ʖDNc[�������pFyUu��l���!�
�ܦ������z�*���3O�r��מ���o���g��=F5��=b�D��y�]|i��bR��^��]f�ޢ�JV�q6�*�RL�߅���:�8�/ZP8�>��/Ӫk��1���U�8s�vOZO��0���������6�^ţù������Z�>�aT\��|5�}�� 8�5������~�N��7V6��W�;V:�W�"�I���ݪ�r�K��`�TL_,iqu^ ��DOc�q��^�}޿��������IbM]����5�;2��m��oP���?H�R��t�����Ι~	q)�*��i�2���W��e�`A��dA"M.l&�x�����9,�5^��+ڊ򉹔(��l����N��Mzh]7��Z`�[g	"::�U��G������T�����١����7�q䩪�q�p��|��h�M�O���M����DzK��m���f	��/� ���V+��>J�eZ�'�C�������`4J�n`�O��l�3n��0RM(�Un`�h�\�\�h.�@�B<mpi����4 �;0;y�7U�)rk�����+�3yi��$�rJ�0a��ȷr�W �-�
�t�xZ�9���"��.�Q#�;>�l��7b jyqZ����=��֗�8�w�4d�1�B0KԎ�u���%�8oo�,������R�D��-��H��ʂƺd�If0U�ME������	�M�]��e�ț6~�>.SkKg�q�_�I�?���w�:Zo��y̐����Y(����0���\�FCM̊NI�⛏��)��K�q�������va���b�9/�ގdDv��M�KM7PK3@�rDWp��el��Q5���?/���w�	+�Al��s��z�&e�r��ف����4�5P]`W�H-d�hFw��ςqS�C�P�_p�=�k��I��k,�yI�Ld�8 K���ܽ|F�.�P���#���v�}ј%˔���J��|T<��Ҕp����arc
<�+�!,<&���$�����+�5Y�(4(�uU�b�b0x܀�VD֘�N��/>�=v���#�3����b
ga�i��Q�����X}��K눖`j��ך���%gFpL���(q{'�q��i�z�(O&��´�"<}�m��\�:x��?CD�*MS���DH`eBzQ��Z ��
H�U݁��<��u��k��쐏1��ob��R��W�5R�;�['�|*K��;�2<Or�_=�V��*n=6W>�T���?H .�z�}3�Q�!�EG����_��n �+���J|���Ӝ��>h �>���0����Y3�����[��$o�6�D�Ҫ$��~�}��wu��|<3�װ�.�-�e*Pô�1���rB��c<"�T�,Q��%���)A���D-ݔ�߮��ʝ	r��m�ȸd�f�����K�6F���ˡ���Q�vQ-q�S(��Bz��(�oX��%�)Jw�F �T��3�&;��n~��~;�q.[�_C7��
�3�f�j�^��WEP#�[�x��9ēj�V^���P�*_���;=n��A�l}�`����<�I���"�"��A�H;.@d������G!�_#�PQ����D�����Nۼ��'�Z+炯�(�z`�'^��K��We��I����*D�B������	��F�F��&�sB�Pr��"9����
C���G���+���\s����O�N��v�@BU��a��{J���`+��U&8	!��"r���q���n�����%���a����C�a>�����j&ߙB���y3��65�0� ��֛WM���H3����rg�k9�#�������Eb�Zm<��d�a��D*�:9�����#�����wB��I�=�þ�����(�F��Y�#�TA�n* ���)�.�vJR����=���H�)���䲃�p0��K��c��|�B�ؚ~H�{Xi�gd:\00���G�%��LQ`��kс��DK�����`)��5K,��o0
�W��'��FM<�W�+�ʰ��ъ��{� ӊ!���Y8�Y���n9��J�LPr���-w��#��%9w�����;���`y���)vv`#��kE��Ǆ�́D�l�p�Ӂ6��f>o?��	P����9K���E-!#��i��.�_&Nid�`�U6U�Q��KP�㽛AĮ�m!���
��(�-��ǌ�m�QWi�⑗S��#�q�{�8�XEӃra�0x��]3BT��K�##$M�B �෠t���"#��
f��y㇘E5Vڳ2	��4������՘�л#d�xd�m�$F��y�ʎ�{cv%��%T��l�;�	Cs6�j�,��olc�BK6`�!s�a����xN���r'ޯ�&g4[;q��E��s]��`_�K����۱��k����2(J<�+�`0%tTq��A��Y�U˘��K2ͩ�i�צ�|9Mi�)z�P<�'�
b95���#�����/p��.� ��vr��E[a����;��w`�&r�b*��
��}�/e�C�Ʊ�6DX_��D�UǁՑ�nҢ����m��q�������֠��������/O{���%c{(�y�-�>�~;��a��(�_Ӟ��Tj>
MTysD���1���`��~/��x|ް/��G�,^����!5�H��3/JF6W|�n���'�ぃP���z�wI�MQk�A�~:rC�0!���%$�e�*@X���e+�<ŪL��ex���v�1�:5���mG+�qR-��wOc����aj���9N&��ҵ���x�w��b��O�����o�����2�.ϡo�[j��Cm�~B$��)��;<�)F, t�)5�,�hҵ�tbߞ�w'��I yzL�r�[�Z��S����!��e� ���_�����U9����f�i���p�R�kެ���?��G�9���s�M\��v�#��U�^���h\w�\԰�v��|M��q��|D0VZ��8�Ҵ.��,�	���g,�x�D�����!��C$uu��l�{x�f�!��X%�R.Y�( UE����D:���j�m�g@ExL����u�p��	��g,�}qն2h��&�V2�����m��wEj�^/�1Ӯ/��FԠ�<��a�K�+�X��z$e��i�������K��Һ��QfJ� q�X�l,լ� ���L�MFB��{C�W&������p���"R�@U�$�g^gY�� �����>sa���F��O���)�� �iz
׈U��_�g�����g"	~� �)S19���������c21K����.����W����l�~(t�����g�'Z��|��l.�v&9����	e�r(��6 oQ/U�����"y��E��M�5l�dǌ[��FB 0�0�	V`�'~�8�m��ë uh%}7糁*q��KU��}�8�����8��?�.�2>�8��eF�M�f��âXЍ�P��. +�߾=�b���z�?�`V�DN�D�����D|��|��c%�����MN7���i���M�Xh��&�4���#F�K���@V/ƅڭ\���1�D�`+v�,��`�@����TM���/�/캡U1	#�����|hk�lZ���WG�p�^�����f�{R�o�mah�zxgmT�|��A�;��*K�I��������"�Ps"ڲ�4��4q���=8A�aD�K���᝷��c����׈Pn͛>���<�L�(�Xp�����7��R}z��/4e��
1հ3�#��d�{Ȑ�ϙ�̺��7P�V�v�R���é�`���:�r4z����Fa5�J5~�ݱ���[c�(����F��r]�y�������e���?��.r�	��{ICS$[Im Ao�ŁH���@('��8��ٜ�o>����
M�0����Ee�0<^��KW��-�����=v4�79��j�͛=>�����4p#Y������D�j��pYXњ��0A���CC�[Rk��8Cu��p�ӻ��:Wet.���9�� �$�ɉ{@(N����*���h���4Vג��mO7˧:<����J��_~� gzˁY�*�m[@8�Gܽ��nI�U��<ʙ��~�y��?���I/2��J�;��̽90���1��*�F�*�O��Rr-�}�(�u	v���MS�ZL1z�1G�GC0�-q�N�P+�l�\+��z9�k �%D�q)�^je��\JB�L�Ԭ��;?MȨ��2��Q�	�m�R�t{���hA~AL�7h�_�@��w:�m���Y�O��@G(������H0�K����_�����zM����r<��.0H��fq�N&��X~R��a*~a���$ʶ�iI�@��K���5�&���x�S�)]���,�	PrW��lo�L�<���;��w0��h�)�:*5�<�d�T��)Zo+���B�h�6�E$�J�0��U��%=�߀% ���|�2=��@�����(-S�8����Ő�'�Y�I�Jt��|�v�>z`����r�t�>>�20�5D�Y0i�I�"�����Q7�����cu.���(��n��+�����uYB�����N�p��&���nZ��2c����@|Ҏ9��yb�L&P��7(�x���6-��ݵ왿㥊@�4ׅO|2z�2D�Jm�?���`�`��r�M`�]�~V�����'�u;Du�ӛ�/au�l�<N����#<��:jN�j:\u��Mc��3�Ca���jNt����l&�o�����w2)�8_f����I� �B԰lڄ�+�yyW���:�kp$U�0�76�� ��C(���@S� �UV�\pg}�&���>�b=!"�L�Y��>Z�q�h��H�-)D��U�8��P�O��U�L,��EIzH�����y�[:z"����c��Ŗ�ռ�j��j5�D�1&�0.�x��
+��
 _R�[�t<���I+6��+T��a{���ˍ~]2�����}��vR�U��ło��2�l���� x]�b�s^㥣l鎢�w"m=��e��'�("�T@���09rVlPg$��t���C�����}c�!�=5��;,|;k���\�6�@�,:�����A�ّ�����S�OD1�YXm�T��/+��(_"��������n�ϻ�ʱ�����X!�$��j��/��:2+��-��,73>�7����;W�R���D6^��N�"U�u߰���m�zq��>��5E�?me�M��K�2O��ש^^�n��3��>A#w����H4#}֛e�����9lE_�L,���t�=�
@u/GB�e7��a:]_3�����4��f�<�U_���~���W����B|6�,�Py��Ԫ�'�R�;�}5:�#��ګZ��Uu���m�uhh<�4�,d�4�;mV��XNqs�a�Q��E_���%%�Wyz���zh g�&��ʝ�̓�u����� ���;�ʚ�W�s|�#��SY1C���Gp�Z9�������n�\�Q��שhGR�êь��X;$��J$^�L��I���P�̊�{K�ħ[�;�lk6�����02�����W^z����k�:�eI�!0�]
~˩��/VY�
����/����T��9V�t�r�t,�l4B���NJ�8�����0�}���e��=�7�牢W�R_�)��]�ލ'�����o�@1���ӵד2�=���^j�H���������
GJN����l�S�Z���[�Mv�
Cڐ��\IZ�:�D	W"�4����MH��ߏN���X����s�xW�;$�x�Q5o8��zpG��ܴ4�������֓|���Ag�q��5ː����މQ�Y�P�ʄ�H���w�'�՗y�)`��,1�˿a�a�s_��v�	ˀ��Y��	_����L���B� Įa�u^J���o_<� �����!���R����xT&�SM�<��N�wo��1B.W�P&Y��lU`�c�$NW��A�����4c
Z�����p{�C�ۈDa�(BQ;l/xO��u���{	���2������-C���+NTp֌�H�X	@*�����\�$և��E�����u����� �&4��r;�2��j��l�I.:h''�m ��tn/&2��-�	���b!��d(��įiLS����ЛC<�V!��S���BF@?��(6��M�I(�/�j���e�ĵPFz�Kz�%e.-V��jrߙ�mt�R����s�\����DܟЄz��|��W�O#�ySr�V�+��M�e�n��gsh����Jn��=xm��,ͼU���^��#,�=|`�L�2���q 9�k���Q������Ȝ}��P����a<л%=��c���0�<��B�1?�?�L�g�S9AɻZ`�ڇ�1�k�ky��]A;5��x�d]�ֵ�-�$ e�ᩫ�P��Hy���hH�3��?�,0��Uњ�v�`dL	�r*�5N�˛�&�>������E���:�J'g(����#re5�u�Q,�g����������;���4� ^U=��/K��G��ʉ'A�����������j����GA���Ad�#U��{��u�i
CP��Y<,�G�#����ۮ�E��u���)��dg�J;��t��]҉�	w0�΀v�������)G'�P��3�wt7���\D�gW��EG����V�2�{�u1Pp��c� Rct��Q�Iި��1�2�/���-����c:J� <���V��v�Q��
R�:�(/���vb,N�$��#�!uS�W� 쵮P��g��URa/<�	�x��/���g�7�G��qϽ���pY�)�ْce��������E���˽hv��g��֥��#<6��/��$�C��Pc�s�a�߸�(i����:�o�i� m�82��?"l%����Θ�ĸ�?)�Ћ�zٲ��L��EL��	6�d�5aҖ>9��Q���2ry�=j���1��%Vf;G�#�Y&��zGF���r(��[��oD$�2��Y;���Ǣ*!�j"a��	~b	X��އ4d���RNɕL���!�MX�f�efW�K��*��'튲h>O���;��/%/lE��N������R�#���w^1{xN���o�\���n��o}WH���MLs��H����4;�x�� �66S������Fď�H{�vv�N�sɟ��M��W,{o��*��Y�Oe�?s%,����>w敻K�0��<�!oyA��i��F�kb"�*�kc�ӟ�dsE�����L`������������GM�Rh/��}�Y�ℂ�ߴa��YB4�5�����hc��A�fT���@8JvN��)�q�{�1�"N�0Q������"��M;�ѐ�4�\9 ����੮�1l�vn��ؐq�����/A�qo�Cm��m1O��e��+��=�:q��a_�T��c0�*�ep�S�_��
�,�Z���7�`�ͧ��[�G��hd�sԝ�p=*ñ|�����1����u`2��w�hnW���8����9��~��dt�x�.͡�yw��7!���p�}>k�^}L�6�W����ܺ扌:�h�s����&UxB֐�`�$w�?J�A�G���*�8^�7�J�ע�z��'k.{�����~fa��K���7��׉<�d,ް��g+L���jUty��j�p��MLڥ�V�djMm�iqD�nG
�rv����a��Jg� }!3i�I�=�RnyQ	�n��EC�}���>i�l|T�K
=���y���,��R��z@;\kP�yU6�;��̭��y�qU��]�X1��q�̨x�OdR�qJ8����'�	Z���"q�~ݰ|�/8��V��m>0��{�VT�M�5es=�����2Հ��;dsI���]$%1�cT�%�A��/s5�FS l�?�Q8��A��}�#']jː��B�R�wEUj��M	��7	k���ZpL]�
�#a�%�T�/�x�
1�V*�&��d�f�v�V�0-(f7�'f�PH���'\��`3?�j��6c0��h|�����MK�j?�omơ�u�5Z���tf���(�=Rm��W��VH�EG�#����b�:X���6B��7&���B'w�9?�5��\�8bd�È?Tǋ/�ko/Q�*�?E�c#�G]�5������!I�㝓�L�H�"j�+)@u1��]�@f?�L̪�ⴲq�D�Q�i��,A{>��w�d�
0����7�D���;�Y�_�_�a����&_�ܛ�M�6�hQ��
F�L8fvL�Ry�F�NS��Ѯ9�Z��b���䃅�=�8(G\	\X$4(�c�tP~q>)'{.����.ʬc|������;��7R��a2���v��pv��X�����a��E�W�w�~�19Ԍ�U�Bm�֘�\��K��":WJ��6�|p2���O0�����qp/׼L��"Y�0}��.'�������t^��q*.��V�VQ�}:��'����t�v3Ƒ����tI�l�u��%�u<.��
�������� �g�
f��ݏ�Ү(�fA���j�sגL#���Ff`ȡژ�?�oK�4SH�`�
7:��B`�{��%k?���xS8� ,%���݆b������}�ʁ~o�lZ�%�NR�o���E�����(D-q]3�	��̼:�;��K�c��,����*y)�'Ԧ'M�4=X݅`. Ԕp+2������H�I��Brp:�\:��[�]����s�R�f��K>$�0���@��,��(�r̉]Qt�U�.Z�Q��Y�(��z���u{ۉR�T$�K^��q���;!O<:������!U�X���n��N)B]�Iz�V�Ơ�G5�"&���C�>;_,Y	�Tk�xxw�y {�+׎���p�i��=.��J�Ξ�K�(H=��Z�+ ���ȟ��|�V%�M/j>4���l&QΙ9e�8�H�B��9��T.�g�U_D��D��l+V�>�ꖬ���@M����.R�fhb~C��8��$���b��$��c���:`O�n�l�5��M�Ji]�3l/��k»-a6l��v�X\�/8�AԪ�~����E�ƛjsުA	���	��觐���Y9�o	��''�b������ �V�ӷמ,�t�2J�E�)&UK,��]�Uf!LOA��_Q���)�We�5A����0yz�T�<��,5�GLs�S�M��aK���[DK?�b��ji�����jU6�����M��S����V2��@�F_�רj�K�MЄ��;���u"��͑���c6c��r6��7�^b�;��g	*��q����I�A���q�sВj�@m���OKM�~w�]֜�9W��������X�����Y}gg���a��?�(j��7*�`A %aɸ�EA�D,yC���1^FJ�b��>�����z�ME:�Y1���˫�_sGS�n!L����u^���o�:h�S0 �jJ�E׏Eg@
]'�xK�3)9/m��J"�/�h^o�)�1g;�F梐Mˍ*>m�x��;ab���䌫��͏��@d>"f+I��׀<5����a�z���O|���6Au��B���س�5C�b�t���^$�dV��|<���]�aN�#͟c�������Z��^I�C_�6	~-�f��[l�Y|D1b!P�x���u��=��#���l=�k�Ec~=�a�Q��sEn�ng��RW^zٮ��X���R�{�Wu����D� *l%k�M��;�;��!3�}-M	�����e�d��DDe�E�?�k%Y��4k��+��_İ��n-���K�!'K���^A���@:�1V!t�
~�wK9���S�r�Sh����Q��ޯ"��|�h�;M>��ƅvD͓���)Ak�a��k:�C癁xӢ��R�g�t���ә���f�D�=aG��W羅N��¢T��$���Yf��Į�����E�$�hRf�n�EhW���n������;3��@�D�U�~���i��#�x
��.�1�!+@�K�����}�#���Q:�9�Uҡs�E5����lKϯc���9y�\����o	�^�_l+D0�A;���]!4C�"�;���	j� �.�K�5��7pg��6��H���Bz'΋&��71���. l5���i	�%���^�'��iC��T��/B�sT_�`�֜c�l˳>)ȞG�?OB�ϯ�4�?-�YP��:�2���"&>211
u,OҶ{��
\Q8J�uH,��k��~��Iƛ�Jtc�6�P���a�	WL���k[�\b��z�n#�^�8��X(�`�Y�C�ƭ��f��WV�����^���cU��y���	+>�P5�jфkS˒_-��í�,��u�+�@�.ȶ5my�2�ģ�Vl��uy��_�������{�U��%�_�6�B�Q:���!�<�L�`,}��A�KӦ����,ޗi�r���RiT�����*{(�q���W��I�l3/*'�u���>���e�����4���n�jQ�� �Zy[�{)_VS�4{d�Pd͋�K0�ag�*��'�Vl����M�5����Elw�
�7��`_�;YU��)�H0�*.�y
2�eq-Y��ٶ�K45�(���M�%KW��s��j.֚w����!��>���i���!9Z3�d�P���z��J%�lA �.Ň���$��ҷʅ{�0"�A?��N╤��~�W��6]!��9�Je���雯v��ˡ C>|S�7�D7c�Hǁ���/���/g�/'���Y�<�=޶�*�o�Y��~lA���
FK�]P��K���3yB!�<&���n~b�89�4$O{��A����V�(4l5���e�;�k���N�q���qj�o��������e��#rV���
��<�ι�E�ꈲ\���� 3��`�����<�Qx��퍱V�ZK�{b�.�)I����''E���D��g=�))+e����x`��9z�ݮ ���Ss����j���7�cՉ��� �Oi�����&�Ld���5�W\`iZ�AUU�4���>�A@����Ŵ��xey6bc������G7�3*���"�]@�;�T���Ywi�`~�f	�I��I��XQ�K��tB:h�;�{X �\3�đr�;;�K�W{+/��nLz&u6�eh�J�I��n��®�����"����V���璓�n�.�)aN������#������ƭ�
�@;U�%_b���}�4�X�J�'%b�Ǽ��]�0[��?i���vR`6�ą\�<0��8l4�ow��6|��O�����\�l��-�����E��h_�0����bUr��M�'[1l�0J�.�A�߫��|�ݾx;�����Zc�h�jК�S�X}s�i;p�v�̛�fc)o/fږ��i^o�%�����i{r�ax�%�ӡy\�7k/mh��'��s�#���Z�Һ~�����	E�/)N��-�����Z��)�\�@4���ra��IdѬ�19�H(�Ej3�I�H�բ:(7W���3��I�;0l����Ŀ��R⟭d��?�rB�4���}��.�i*��������(>�N�컚g.��*��)I#18�ks����4'py.V϶j��;\�	��sN�9j$��E�)�*S��H�e���q��3��  ��Gv^�iaI�Rۉ�	g���"��)�R�Օ_��z�r�AO�:�/�EWR9�-sf/��|�iq$dz�k��Һ�{{�x��- �����|����{�5DBF- �3lo�P
���"S�g̈́�t�6/I�ŧM���T����.�F��}9�[��h�\*�9B�'�!�4���}�����JzcA��\s�ťK���BNn?)L�]���5�a-���m�q�Ao����q%�8{�V�[��
�D�NH\^�LtQ�.��b3�rE��J>x���p�]�e�_y�!r��
��QH��^��J��Sq��bw�53!No��B���U� �P������:Eu�\�߆��T�]#md�c�硄j\q�4cP�K�x������@���e������5�s �B��o#��g��*7��Hl��i�,}],���zԬ�(�*��[�)��ؽ
��iXyGjt>YF'.�;�׽a�j�/cn�b�����|�\��j}���#�"���^kA�A��t��I;&�.��'�T��a#��Ýĥ��	�St��憦����GOI�JJ�����S�n���ϫzSf��,���.Y�'l��*�y�TœiZ�e��qh/H.MmA�$S<w�ƽJJ˅<j�~�ꆫvs�<���ΑbX�.��u�R���pB,&��̻-""֥,��������yV=��Cr���(���O����[�Kuv�h�⚞i�m��9B-��4I- �ɜڢ`2ElD�7A�QL���c���Xx�'��E"/E_���sE�+V*�`�!��Z�X��ۿ��>�O�V�.��bΫ:�Y�.���z~;��$�8��4�W�:����K�K�$9TPtq<�����
�1��mI���uD[�pI�����{��F�H�� o�P����c��Z(px8
���Ļ���g���3P��G�S��zx���M���8�p��\&A����K|�����8���3��q�/�gǮ���/�%i?"�(�����s� {��7Ueߤo��9j�dN���5NM2���G�&1����O�=s��;9���E��u�����,��4��~�o����l�u��P��) B���hA;`�8t$�Hmu���2ؠ-�m��{��O���X�'ŐcY2��� P7������5k:���i�1fd�=n�>i|�MZ��.�q�辰ﺸ'��]`!%A.aMC�#��>�ғ����Фo�(�}��(�!��t5�)1�U�q�m̭�QKi��3�vWi-	]�����㠱b=i�R��S/U��iW/�i��1I���V��̊2��YP �A�5#n
k�{�|��*���P�S9=���Ӛ;"�T P�I�xo�h&�O�_-�V�¥Y��(����̈���gtT7Hl_�sOKر�x�,�8�
-p�
8�
B�;k��?�9X�A⒊P�?6�$����\�u� ��sZ�O���v��\Xx�8wO��d����j¿�0�{�
V{��gʙ����*2�b2��Kg�/OxE�,.������nGj܇<�U���f
=Ng�������h�$z.t�8��bӏ)��Q�3�fZ��������3f���cQ�i�,I����c���b������j�8�mtd�ŝ��!�<�^pߺ+�����󶪫���=��&s����,oi��$��lPB�q��=c� ���f5����C	��oP�1�x�$q�c��4�`e"D[>{�Fw��f�so[D�rSk�C��b15��Ʒo��ám�P�����K��+�����G�+Z��)�  ۞��
�'��s��\X�q=�og����T�(��ob�ĕi[;t;r�7l8�~T5Cz�J��@��T6��E P����F?X[��lD��i����23�"憏���[����(j�Z��Bf�t[@��Ng�y�ݡ�b�A*���;�=_,��#�pWQ�I�6��`�kn�#~:��x296���%�
�����[��$�����Q�#a��4a�G�`��F�w�M���<"P�Rmi�M��D9���|,7�{|7_��7�����^�i��S���_�|��e�I�"+2_>nS˔zc���ڰ����M2� �;�1+�N��0�\e�E���D� <u�����k��Gٗ�`+	U4ō���z���YV$�,�/�Z���z��J�%[�.��{��Iu8�I��.�V2��ŵ���DF�:"���Eo`r4����{�e��j&FIhie��Qq�U�X����&V�Z7n.*[p~�m��V����}&�$.�_?��q7{�'~��� /r�[`.��<�ߛ�ǋ� 6��l�?H0!m�h��I�q2a���Ӎ�J����4��4�/׵�|�٢�M����H�k�|��v�37'ɭ3`��x��`��J��Z��C-����#5��w�N�Xìv������珒(�Z�JE������Ȅ^hJ���d�7�=>I�u�u53,:ZEJ�E�K���U��U�
�
N�E� [���L7�2��Ù���<C���1�����X�� ����V�s&0�w�:D������ �{3���r��G�Z����Z^B T֔S4�>�����;�4�ӈ���d�H��y�:�1��
�ֆ����pj��d^8�	���֢W�ףvPŢ^���(]���0ǻ�'�J�B%��ܭGi�&1�!GHe�߄�ӳZ.,�8U������G��ҭݖ�'�C6a�/��S�ģp��JZ��R��)��^��$��'�l�"V�O��䁞D{�.ا����_�Mp�t�!�_j��B��=�h�hPM%�A�BT���"[��g_%�n�u�~�*����dWA� �ߧb����s3��ȉKzZE���q+��nj-f�$��ӅQO�v�OU����I���j�n�PO�)��e�Q$2���i+hd(�0�ߺ:�
�ϲ���m{V��c	:�B�������wyuޜM^�B�Ⱦ�=6 9n�BQ}�a�w�fO���('��Pa���u����ڄ03�>�{�?�
�|�h��D6��=]�-�
�0nܫ�ƣ���a���ڞ�v������xS���-�4��3y�],J���BmZ~�7��qg��c�+Y�7�WǗY>eԒS�T�)-0t�-�nUrJ.�ɺ�h���;9���-�F��W�3N��Wc���߬��f3BnW'�T������)��y��xL?l~?�9�z�L��W����
�r �17�0Q� l訆W��hGD\���;N|QHh��'��t�mh�G>��R/$�2P	�����46bB;A�*jw��]Pm'7�⮋J��4Ǌx�����5	�I���*��������+�k�� ���}�L��#���
'蛌�p���E.j�%�8�P�f~���ԳP\�8U��g��)�o�͏�f4tfv!�&b:@�8p "���<��P�RΈa,�gS�l�C����Tm�����J��
������? �UϜ�b�B�Jfn�$�bz��@�x�`p�O-DC����ӟ���y�l�=��^=u�Ϡa��s�Ѣ�I��.�X
D���>�Sb����l�lnx�v�h��B>/G��[��4�d�WE����%Q���9#	���]�׏�a]V��t�:پ�E���$j�mU6�׮��C;��j�2�����>�bɒJ�*�"��F���#j�R�$��YN)B�
coy�q���L��5���ƿ�n �e(�-�'��f��Y�Ua�;�f�G��~ r��^�����N�*uI�4���
���a2(0"UM�ц.	��U0�U<=�vh��(-5 .�>c��YE�ڦ)�J� ���0����pl�_X��շ�ю�%RQ�ܱ��S��
_���"�SPU�ɿ����X�[�d��&���OƱg�sg:SP1�c��=����w����-���=WN4���j�e�ړ8�_R���v����"��[����j_��2Gý��0���%�������Z�j��t9��=�w�L�mW�Jo�+� ��<ka���v�	|_L�7���j�h�U��rjw!&:���僔Y!��J9���u����>0
��X�WsQ�6� �>�Mڢ�ЬP���a�	~i/I��z��b�;�;n��PGxo�ݨɠ�t���8�̳� 6n?M���prҟ�8��y^aڬ�hSXf�l��&�<��Q�F6�jب0c��ώ�_�I4��4�.~}Aeme2p�XA;��S�i�g����%n<�e��D(��M������$���v�!E�����T����>�<��u�[��P�`7F �m�C�q���fl�ǳ�m�.��X kH푕|0�ѷ����>�ӽ�BSmfwb1]��fz%l�E�I��9`)գ¢Bv-'��j� �KG����%�H#˱���5��Z�sb������M��]�]7�d���1�:Qz�رv�~Ƥ����Z�y��=с>�--�����x����F�.��+��gO[��E汬6���J/6�a	0@�_(���կmk1Zq΢�s����QZ��9Wp2�M�u� ��1��gr��|�)"�c�����H�m���\k����� )�9�き4Ч��R��_Ͼo�؆���8�7�{�<M�N���.��=#(�`k8��ws3u[8X&r}s�}��p�pf`�.��fbhځ��M����������{#$6��0�ͳ�[��!��X��`5Wi��@������`�5�x�� ���׽jh�:�-�Ԭ��`o	&���{(����y��P&��!�+H>�jʟ��໳�Q��%�=��xS?���.�F$�;�s����<B��v�&I!�ʿ�^B@����
x��A*9q<,X���NZ��X�wDR���%VQ�������zBP�56Ł߀ްd��,�^��e���?k��.W>�?��\�5t��i������Y,X|�u��p�V%�J�Ƭ+.XU�W���}->���K朄������"�G�?����%G�o��[�tIK:�������c�!i9C���,����%x��{��C��W�C�ý��ݜ`A��dg bS��B�BV���X�9����8�~��g�(�/��)ič\�L�D��Ǥ*c0����4��fG�sg����'��(�������O�v��v����1�y�����9�N�'��T�]�9���lrn�;9��Wޭ�e�J?7��Y�k6s�U��N�c^:�n���*��ɺ i2�%�䐡}�l���g�U������(?��D}����o�c�?���u4Jl���"��l�}�uOʼy��5�=��5����q>�#���R�"+2^s�6���7�D��WH?�#�Ɂv�Ğ1Dz�ݓ��V�tZ����ݲ��Òi(%�Qw��_�m�� WhcE7Bmm�#qGe�9�����Y��ė{�`���t����9!�Ǌ��̦jz���s��Sqh�U��-d}�1ʎ�v1���ġ��������<¹��C�K��~cE~�.�+�5�s���WDd�))����~�G���j'8g!��M�T��
�zQҢ�*\���UJ)�{�ﯳNkR���|�'����4�<�ē6<���Fw���YeԢ�V��o�f�+\�B>���̨�ݝҵ���������{*aP�Nν�=0ҨnT��'"��y�y��顋�������M�j����Y,�H:O�,�!��a��k�*vE��O=L�����{����BR����2�������K����ށ�ۀ�^%Q���X���q'���h�'	_��e�}��t;��v�H���h4nr���; �0��;jy�q���18E�@�S
,���<�/z�z��!�͜�� x����<Wޛ��5^��K��b�-�%�6�O�Y�OoS�Z��$�4@}�s�sv@�,w��e�om�����lM�cj	��nq����������V�*��@��!��޳g��v��ҹ{��
.{M��\�\	�@_%o�X�&��T�K�	�����QՊRgK��U���`�+'d�X&��o#K��&&�2�T<��T�3k�
�i"�|���ښ�\*K�g�j8At��@OAYK��[�پL���ST�FG�p¸@\�U���y�^�� tQ��M���*LtV��bqϱ/`"���O���cB��A�5����U�$��`�QnČ��NIq���	cc����7b�c	�W�("�37kݫp�9a�=�4B�Zn>���o�
^f��K�j�3���������Ԯ��3�0�'B�$��{�*YO�H�6��;$~����k������J+�R*�����f���"_׋)Oϻ^S,���b�$��++[prc�-#��7����MM����8n�8�+a�˅ǩ)��Î�/�qZ� ̈́=ME���-Xr;��q�{�F"_��Hj�ɩȀ��բ�@Я%�Q|Y��2�yܾ��uW�Xo,W>!�Zr
��ǘ:�����+���IvoY�q��&W1^�Q+n���	��f�k�s&�D�E��&]����2��*zצ�n�	ܚ�Y������+�?���y�RG`Q�T�]=1
�����U�'��g��� 49�溺���0���ps\"�"Ό��ծ����"�Ci�4��@������bTl�s�6b�lPI�)�M��8�<�l�����0èd/3kGs:�p�9� "�G=�$��*p�i�IH�;oh�iD��4���A�DH��ܓL%��\���ʣ���\�/Z(RG���D��X�e+~+�g_f��O�S�zL���FҨ�6���q�$��g���qK�CW�6�2�y!�k�E$�`����l�'ux��WK7�J��È�*�h)����$��z�Tu�4=]��t�FOd��Z�t�&*�;a�G�)�{���<�Q�y�&��gܺs��Z�\"����Iz�؉ݚX/>�E�NeԼ5j�;!�pB�ŋݎ������na�T�iE@�m��Ϯ����4��M���ra��)ei���`�ld1�o�A0�� �[G����	��| �zn���&t����~wD��0�p��~�ܯ��r�)��QF&	�X'���%�����)
�Q;j�C�bP��f��&�B��G�A�4]Frh��Ը}S=�w ����9��i�σ�,PZ�7�+/��	y�8?�dl�42�y�P�XU����������X�QGl�"W�a��AC�Z�;��`81P7���Vi_w��ñ�d��\#$a�P����ߥd���������[�@k���0��̍�4�כ3�Oc��SN������_?Zy��<��0�P��]�w��G���o
�<��3Lvݥ��u������F$���*�E�ͭQ��A|v,��q��C<��N��S�ݱ&+j�n~D����y����6��ᯅq���xQ�dA���;7V���Q|ݩSP��Y��t��n��}�%�	a��#�,�`>����T6�T�G�MҚ3�,�kע��ɻM�6��[1◓U� B����R,��7�v�2�l�(���LPb���7L��?�CHp<#6A�<Z%��\��ї�J�9����Q�v	5���M|���[$�ސ�!u��I�J���t�Y�M6U��5~C�T�A�!8�n�XwڐE����� 9��T��巐������)�ߑV �7C�h�P��x+S�g�@tx:�lc��F`�y�]�ƾO���3�/sZ��s����K��Է��I�X��}��?����I���@���0o�+]�Oz)kU_�n����l,!�qC���if�e4���Ս�m������җIŚ�и�r��/}��S�:�)�Ԁ�8��gI9QP�9�0�t���L�NG����p#�S5��L��K���<��U^ϱ~��m:�7���l�uW�:uo~|W"�v��
K8�����F3X��������j��5Ge�(��F��Q����'R�dO���U{I��~Jf`>~���~hU��VL����u�
�w�i��Vb����>B�h���_umgX�Q���49wT��N�s~�cX�C7v�5��Z$Zs���ǃ�K�ip��8��8 Bh9��R~V�s�c�z��;��J"�1�}+�]P�q��\� �j�m�&�|9V(,#�;��4I�(��̔�d�/�5�Y���T}W/�N&S��Fg{̖�"	�
[����C`�P�� FR�$9�T�P�#�f��:�`�D�uu�'ɚ�� ���Jlc�iR6�ǈ���'�8���ʊ��4�yn�\+#UHm�q�t�i����r�Q�HƵ�������sq�g�Xd��f�`53�2�	D�n�a�溰���dUp���7, k}b�:�/2	?�kG�7�a��t�gM����e����O�Ѹ���a������yō�E���y���U�$�G��q�"}0=1�{QN�8ߕ�@U�j(Rw���)��HF�%w/����2T��2�'Rv����'�N�R�=5�)#+��FFxx�'K���g�zt���Sg����P$��UI���\�c��h�K����I3�bI�����~��+�([�� qJQ��Nm>�W�QrZζ��v��^�^Z�E��É�����
=҂f�j,�6e���G+�������#r�q�V��N~�V.��r��T��rA��"I��e�x�tj�Ò�Do�MML���i�CZ #�H��baȄ�l
�i��Z���]��%��o�O��)[Q���Þ���]8Y;~r3\�)[�kEX(c��{2�z$�FE���`$q4y�^�(��(W&{W�(��lG2�.gr@��N"9=2,c�X�H�,�6�Ĕt����?T|zC�R���i���%�i�iYք}�g�J�A���dGP&<��wE�^Q��r�[ �0���Lg�Dd��
 �� �O�h��h�d����Y�f%>
Hq���S�J�66��0-F�=���	���N�SH���FÅ/e9�j�*ܧ|`ިKq�0z���af���䓳h����ZMO"EO-�>�	��dD2��o�ψ����=5&�5O�Ik��z�O�c����߯�������I
M|p˧s��]T�&�M�1E�ש[�N~J�f�X/� >5c�?�\�s�"5L7�W_�ӊ"e*@�{�UW�/8ck�J�az�^�	���&�׉�\8ln�1��,����� ��mP?����H�^z��)�F6�Ƈ�}O�o��0Qe]|B��~�j'G���.�5w/pP �u��G"��Y�b��7��s`��]��6\�PM�)�8w]}�>^��d��2`��i�0��ߗ(�_U�PJ��}��xL�lW���\sX��U��\(~�+���O��yX��cAR��ܟ�G���k|�,
@;A����d�;f�JM� i�z�!���!;�q�۞�χfU5O�E&O����.�:�Ow^���m_t�pv��1��	l������L7[��4�O:��sX�rT�d%�z��l��J�n[-2�^>�m-ȇ�L�c�
�/X��n,t�d��!��0s5�d�ڧѽ��K�~g�#����!B�\��k:�}�A�N0J$��>v�Cw�t^���(I�^OG�J��+������Ũ��`�L�iG	�2*G^# �7@��)���\��
�l��E�W��hB�;����W��m �*�f}+�<^E���P�!��h������R�[����M�.2�h������[����"�B�g��
E��@�y��F"���"�"xy�
��Tx;�n�U-�x���x�]��Q��?~P����e/��U���6��X�,� %�Ur����OL+[Q�v_&�P�Ց�x�z?���f��U�@�LD\N#�å�9�|7�V�N ��]��p���Y>Ѯrj�_���Ig �nJ<�v����3P'K٫;w�ٙ]���v;�A�=�>�PaD2pP�Hc50P6��zv�'�>^�ϕ������g�l���I�N��I9V���i��B���<��^\��̍��}*����z�ㆼ�8q�����g�b�c.IG⌶��Nx�&���Io͔�@I�=���|Q��>���$p���X���qZ�<ê��t�չ��@�w�Kd�F�C��;8E��]��d�ZU�^C�áͽ,Z&5���� �! �� �K�j�.��@�p�"�e��A7���{=E]��k&f&ͬ�-w*z�C��s��X��;�4B���v`�s��㬏qOo��|%Q��*y��xZt�Ą�7�T� �}c��QIֵ��~�����_��=��v�C���z�IM���\����D�u���+ <h���)��*�F�7�GQ��M�Q
'J�����R$.}T��Y�j	����IW�c����R(`3F���{;�A�VA�Ri��m�1{Ne\��,�1�*��^"�B�-"����9���b3Ȓc4�'q����D������r��d1!�aGb ©��Kշ0������&|�2�������Ҷ3�@H�p��M�~�����N-M�3�'`�P�0Ѧ�4��Nvm�a\H���-�R}RҢ��*������U�q�@�x e�Em����zʔ�'}~��ëe�[fm'jN���u^2��'���:����x':�c��?���M���N9S�X��Q�+�#ث���)z����@Tq���m����!U�]���BB�&[ڌ_�5& ��2A��d�op��x��-{(SO�?�V4�D]��Y����bI� ��'On�7F\�fUy�%+�ݱ�*����	%�D.�;r:2�?0�Wf�8�'�z�Sq����,�*���E�58\�=\`Ej3�����VX<t�M�Gص[�|�z��}�W�>P�Qfz��� ��`��;��_���9��,!��z�"[i�*u��!�*ȉlqá�y☽j���ȃ[�*A�3�7`�c�/�쩥څ$�"���E���1;�^U6�.��M��ZV����<�8�w�1�V�z,���*�n(�|�	�+ 7������C�ő�v�ڊ�
�;[��(�x�mWiɹ=�1�U�������"�ހ���wl�N��2b�Z|ٲ{�G-Rhܹ ]^�dM���,%�W(���r�����A����6�	��d��=��]�>nC���[�>8I�
����o̓���Oޫ]�[��6��Z�	C=�c�3�#B c7��M)k-(tT%m�!���m��LQ���F��N��_7���.-�_lކ��Zc3�Z�����p�r��ϕ���s�2�'ןE���{�HєCUW��U~�0�B\�*c��I@�
D��
>��=?�2��ϭ�%x�a@M��{�a���F���l@�e�w�F�o��>��+����2;�k���'�|���1S���K4��k�R�!㜓I�)�f�
]vp���K��]�����M�&�����4��j��]����x�>�-X0!X. m��ݝ�&BJ�ld��Q�o��D�up������V�>�6�]W�S��l�F�Ҷ,�CPK&݁���<joJ-�-F<�M�W�6�|�$�~�ݶ;�*��+�@-F���8ݶ-����#P���#���Xىxp#)�d7b��srkSL�E�Z@��po��Α�p�\X��$�L85t�C����;ص�Sm�e�lZ�����������OOC�����N1=߇��3��=+^�j�V���Ȩ$�k�p�y!��c4l8�ռ7m�q�
�KȰk�'&�5�~�+�EҮiC<�/6����:��W�_��ݬۓ[�r+�L8h����c�����4�� z��3(^�a�	"�e�t�D�WW���ͅaa�P��n��W�2����;VL���G�� ��6�5z�4"��Y� ��Q�n�*�}�֪50�f}���	�1�3ƴ�JzU.��>i����o��9\�`�d�߻}�-}Ʀ�P�-;^3���7���҃_r�/%\6�շ7��vO�����-�d�p߶�JZ�QYf�c�Q�*�������^#1좍�U
�I���,�Q�AԒE�L]͇�G[�J��m�bB�Οи�gYΨ��wNB��;���Apڜ�K=���پ.
�ZF���ܯW�*W����B�3�!q�ѷ�B^iS�n6�lѡ����B���k�e�K��3��>�߹y.&% rN�|�|���gh�u�W��������4*'lr�:����C�,I��w�.��u�E���yA	o�9/?�kl̟����z���5v�*h@�e�Q��j/R��cQ]{�&�,��7��{�L����fAR�oa\�I[�o	L�r�1��T��pn��陦.�F��y+OD�����n%���y���#B����!�ƣX��ޟ?�����^��9����B��j �vDa������*�< �M�U5-��+z�4�|9VU1Qy͝��(aS�9�x��3�9)���l�*@,�DQ�t���c^�>��-;��]S^�q��خ&�Mlx�����)I�Ԩ]o\�F�}4}v��,v'%��e !�.-�䚑�R09���S�ց�/
='x����2�Ƀ`�6�ov�g�����/\�O�p;k�m��-��	����L�z�I�b�F�jG����A�}"��I��S��{$�n�c\��(F�b�S����ݔv�fv����R�Eѿy9���p����ڡ�DdZ�L��m�[T�.F�B�rr��ɵ"U��s��8T?aT�U���A��"�x�Z�ú��X��4Wp���� g�g�鐧vW�$'�����t'e/���%&��n<<�?$��7�oF�����]K��j�\�����m�K\�j��{fs@a9&��-D�l ������ߢc�7\ӌX�˩����|S�Dj�Մ%�f�(����'I/��:�K#/����j֢����j!$qeu'���Y��	o�ذ��)�H@�c;�2��i0��~O���~W�&K����f:�?p���op��Z͆U%*V��{؃�.}��;/���k�}�p�K}c ���[�AYԹ����)��I��S�X�46D��~�Q|���̏��/9�Ց~cPzu<<咺!��{�᱄�0�@^�_�
Ҥ��Oy[��L`��jFB�7����}�ԫ�h��(Rk��iLw��>��RS�r�v�1�z�w�-�U����)[ �Q�����X������/R��= S!��lэh n�LmE�oD7�O�c:��y5�VRP#ڀ��l;�a���TJ�i{��/�wy�=*]-���=z��Ñ�9CB���Co�#!5xd�Ƭ�W�@�B��H-W��<*�� ZDF��_xU����[�숓��Կ���l��SO���S��b\�z�4���r�<�D�ɘ$&�X��A����;�l�d��D<M��9�v��{fR�"��D�<��K��Ō���Tl�DU��呵h`g�z^�.�T!I6?��y��.�Ui����P8���5	��p��ur�*���G9�p�s�� ����$4�����s��4����~�M$Sm$�^)�7�1dAp.����.�<�'��0��z�E�mr�?z�^�*r���J�}�]R#Ȯ����F�������_g9���M�X���<a�\ۭssS��]x��rd���+C��n���Nk`�����#����d2��FG��؈�2'�5�8C6�:#�9�
���a�[E��Ȯw��ǻ}P�c��oX#��"��'���N�����æ���Y��X��i���Z���戚��oZ��6�-��	'o"����ޡ��-�o�[h܀�����u
5����)�y5��bCuƙ��13%9��x\�� *aQ����� ���^Ļ�-T�M�J��e�A/�L$�_-E����2������\����,w]�aO�'w&d����,屙Y0��bܥ�Jy�`}!˰c���w�I�M�X�tML(_���f&V������5��=z���ML擗�{���7�Q	�OεW�	I�/KI�&�؆��,�4�4 5s���P�Aq��؟��0�U��ZnUq�=�zp�2em������;�OI}p�>��ܐ~��q�p@��v���qY�ƿ;~Lޘ&;�c=�u��
&�m�O|�X0�ՂYZg+�r���YҮW�3�k��Z�3o=�e?�~W�DV���y�ZmW��>��
)1�u�Ⱦ~y5���Kj�_Y	�$� �+v{{}���V,�����hoY��먫-�7�����hBC����:��'������@Sl��n�?[Y�n�4���}��1��Ҳ6Lm�æ~�I���n>~!���-= ���f_���d(��S �Sl�R�Ǜ�S�����*��7����?���I �Q7ժm0d�RS���Kǆ#�@���K|�|���֙"[�p�E{?�n(�9�H��rȈ��c��㸷N������"��"�m9��6��rL��f��;U&.�fvu{�<�A��x!4����kp�����|�a�P5�sOs5J�g���%��~[�%?~ C���!ObS��KF��r��{�?������'���[�����
75P��Z��_�߄�=�U�S�z1bf2�o�(�Kq������Hpy��
�:��`�̪l�uxd�_��).W>"�T��g�1U�%+�Y����?� �p�&�RT��7�����p3�,�Ŵ[=�w'��~��,r-�b��o�������*�#�����Z�$��ȅ�'rw��&6�?b\�VRm�riQ��D���d2�N�ի)�-`Y_,R"x�Ūu�o�����ܡ�w �˾�{�����#0ُE�wP#��Of�����`h�C�K��}����&-P�����_�Q�7��m�!�$�m�g��J�'M�:�'y;q���w��t(E+�U,jV�Uc�Ѻ� 
��C�',��\o�S�}����`kk%u����v񚍍N�k��6�9A�L�e^ZS����% >o�>4��|dZsC��-�`��z��[��ĉU�V	�H_�K�W���]*�)���$������F�b�T��q�ΈT��e��z���p%�{�3�׌A��w*��ӎ��
}I=KH*�	-5�H����f�φ^i��F���K���c��&֑՞7�z7!����7�3hƛh�+#!���e
�Ax�m�ƶ�=΀a{�3(�=[��>r|?�5�2������~o���i,�n0g����$�Ř!�H�h (	Z�"��y=��:S.��qX�@�F��ޛ.�-}��Y̷���"��,
6�Ԟx��O�q ��(0i�{��R�����G�y�T�*܀�p��$�z[�ENL;=��-���L�b����>.�&�̄G;��
�-��s�\o��,��X2 �뜝�Ʌ��!e"�����I0x�ibr�5�!���q�:����P0�5C��ݵu��"C/�&!�m� 1[94�R��`<�8�P��'�=���y�Xɫ��}��Hj�25\oS��B�4��V�G>��7���p�?}�z���D���pz��,�;�X�s*z7�<~Bv�vÇp�_4Hs+��M�m�W">
M�7ُ���~+,=]����Q}9@vy�X*���1XM�L֙��ܩ����W����ڮF�w#��u���5�TdA=
�f1SR90��]פ�h�H���W=Q�5�=���@�RI�M��%�qj�%��x���g��
}����g��A�b�OLM8W3d�v�a�"�3���UlO��zPǅ�;���U�����x`��
���'Q�Ԋ��y4���E�3a'FL��X��,qNC/
�ʹ�̙�c�f�=%Jmb�]�>��ܚU�h��%g���Q]\���(�jg$����FX�9Fl���Ç�5. �(Tr��It=�'�ݩÚ����	5��8=��lX���$B3��s2)t���Q��n�.몮��L��d`�D��N�8	�y�qJ�7Ғ�Qb�� ����d.��7��*��Vͷ���dB��o��d���c�s��b|�+�o�C�]Ա����_��v�TD�o��i�5��U3\��O�\gF'�#��w;ƓS�hL6�+9I�6M�]�"�[W�F��Af��-(�۬�oӊ2*Wiw�<%	�����?�V�ٜ�#NF�GªT=@���0�ٶ�o�Ȼ��j.����d;t87kB��tL4�$
��1��%ס륁)T��g�I�t*F�����gu6n`���`���  ݩf�@��ve*�y�H�j���n�F2[���
`���;����9%7a3�NQs%azm�wP�?��1��^��x�>�a���l�W��R�kd��ɰMUV�s{AI�{R�m����G_�ư{����� ���%�J�-�Uƙ�$���]����Mr�qw�-�;�`j;�LH���ݙ�����R�t���1��h���86s�8����4 �6��c�2
`X�i�%��ZeY*��b3���)�XkE���4���ëĐ�mJ>g�yJ�i�����W�����cq�C�{f���A|��8&L\�w^��Vx�p��\F����=1.q�Ab�GQs��3JI��uM&�LH*�Ou{����}ͿvM���(���R�h�{>r-���9Z��;A�b~Zj���5mz��|������w��0d�$��o�+���@c�:���$&x�3��a"]*��9��X��&W��.�t�k+6��>���VL�5�]�7��nbfgz�+]���`��:�~��Y��Y���(F���@ݳtԪ���2.�)���.ky�$�`Zl��x)n��K��~�fg��1���Y� �M ��z:A�}<�R#�������H�ޱ�G�@���&��⍿�����<�!������b�#�2wjs�hU��6��cXx�T��dz~��t]q�����3��4.�\d�u�l�C}wy�w�/�OLK��If5�GJ4�X����"󯧁A ;�Z��
����0y(#�V��(�_P��ت�Q��l_���
&Wk�Y�a6�ք|]�uY��_D�v��a�%�Ĕt�F���w�6�A��������myh�|��>9��l�6�N�ʙ[��)�\���+��lo:��)S��l����8������ϤL����K����҂�&)��t�{�|Ĭ��G�s'h�g���$
-�9}���4��1&	8a�!�^��݂��<�ū�p�`�(��L�@��)%S�{��K=�����88ԭ�8~�C���:K �`gIV��B�۳��|]�ԧ�99XbE:o�������啒M\��.+�dkaե����h3�����_���\��tXAhK����hsW����wj���iC�9
��Du���h���'cI_4�������UČd貯��
U)A�x�	���Wۉ��k��F
�%�wA�v���������]�ǊcM���/|�D�kl˨��O�Ŏ��]^U��]���B�}ù�Ĵ�gY�𻽐d)�=#�T�@֜�����t�}�$��"^�]��	��V���־5��o�$�a܇U��.f��Z�N4(o��ĄS��~��c�p�k�c�t�1}K�����t}>����A��Hܪ-t��M�OvBm^B'H��A� �����[���I׊O$W��� �^��_ci��a�w�.���j^�M�=oe58��`(��6ݞ��:�y0]�w�GHL�e>�3hk:�Ч�-GpUn�%�{��Eȳ�h�/.�xc5����1�1�j����KS��m�X�3�S>92AIC�+Үh��m�
]/W��,f^�3؈�/p@"�b��J�G>�+�Ĩ��f���ڝ��P�G� 4a��
i8.��H5�*�&tGڀ���T��<��;G��Xd���7
��=	�K��b���p�Vvn�����xs��+Zgg]M��q܏݃׈��@˪����F�~�'T|��ƗF'�߶��켶@�rM�-�$�bgh����~2�9
Ļ�ߚ����������.�"��]ƭ���u�.��A\IP�c"i�:�8�ł�{X#�6�d��옒>S�T~����5�����%`������e�2�3iX���,Af�+Ћ����^�o3�/ϻ3�(w���4B.� Ȉ4,�����|�λ���^=�$�%��O���D*9��Mf���U�
�Z�~�Հ�;�P��A�D���5��U1~�RL��<.;�.,�R�Vt� uC�0�����R�:����G�w���^xk���.(���2��o�f��ߒ&�����.��� ]�B�pX���	=j���o��c6#P�ఇZ���#�%�n�Z,���'ώNI|Un�"�Z�� �����	d�?嬑��lV
���;lo6�@ �b�hM"�n��"���<�P�`�&2$}�T9�'���CD�4����]=�b-��$��u_���t����.6΢�e_��]C�,Q@�	��X����d���1z��U�l�X�n�'�1ϕ���y�Ţ�+A����k��/c(���+�x���!�D#^fqU�]��@�V� Ꮶ���9��;�@¿Q��!��P�^��u�4���|�O�����f�]R��U��K�����]C�q��p��%o]��1��lƯZbN5�v��:�J��ľᇩ��O2 Q��5D�bٓ����(��z���{3O�P&��o����g����E�Y2~^I�k�ݼ�o_/Un=DN��0ו3�坈0�(9���&��~�7���YZ�0E1���q�Bp熝���x+����~-ZM��a�C�e�2�3������ybV
Ǵ++*��O;�@�b�]j̠jxԗ��#B7mϫ����B��T� ��A���՝�F���A��E��^3.��]#_zx�:\>�,�<M��Ʊ�����"Q[}m��֔�Q�ݍ=�9K[�Qbqj�˕��}��a�~vit�O�w�s�3��>]C�M�PO�kb4��F�s�s@��1�y'fL��);�eG�+��m���z{�'��s�����8�+���9q�r�p2�z>������mi)�����Id�ZA*�ǞvQ�x�$Ut��bM<�֥��j����*�O�%,Z�����8���T�riT���Y
�9Cr9�N�Ѭ��g)3�/�;@�9�P}j��'?%P�t���m
1{�>�b������#9,a`,�3_�( bSZ�!��_u@�.����o�K��!4<=E���'�JӰ/"�W�ub����e�=�K��i#؋�t M}q) ��QU3]R���̑�md��znb�z�����g �������Z��� 
�����VN���ū�G������+Z(���7Y��o�w�Oȴa�o�f�{��:-Lx^�h��Z#|�a;�emjg�АLnz�f��}�3�a���I좝b�cf�u�W!^������"!�A\,�I�ǐ�ppS3u�HS�~0�66	�N����[ͦF�&�h��g��-�������nYI/��Cړ[k� ������ٽX�n߫�i3k[�k'�}7�%�X�XNG��1zЌO;!�9�"DQcӯ���L�r�P~�X���Q�z�7o����l�����)�_0H��C��)l�)��:�D8i� ]�|ߔR�}G��?�x��G�c^�_ظ�C���F%�l7Z�{��+��]��Л�L��Ө����)�,+�gȄ�R��N����l�y�n�yca,b�Q�]��-�����c�����1��[ˣ�(rta� �Ŗ��B͹����zΖ���!(}��.//u=����[��hKP.�oo1B�VM�N��m��8�oG�p-���x2AOO�/�Bg�8��K��4���24��e<3��wz��%J���ILȫ+/7�Q�%���וî_^�'���RQl���*���1�~�Fi�����gWY���J�4WT�{+{�ǉn�*0�W�c S��ȗ��~�} *�i��xY5��F3�D�/u�L�ӳqØ�cC����NEY��A X^��o6�5�e����x����|�S󪄊��Ym�D;�F�̽ �ɴ�8�
3�����\�e�]��Ǻs�}����7���g�����b���HBĞ	9k�v�G���0%|*e�vŚ������<��!IUs��#L�'Xc�{�s**!�k2��F`T�5�5O�ћ� ��1�B�$�i�^%8��.([�� �:{ϳa�A�S'���6@�JE����/�.y��9�;�ެ�J� ��V�q�Q��P�lQ7���$0��0��r} �E�,.	��;��H�2�z͙���,O#��M���QG� w�'��s�����>�VMI�8a��(�IS��0�q&�0~��Ư���-[�\���1Q�֕�L"�+W-k�������'�*` ;q�.�`FC����U��opu�Ѐ.#�f��8ŕՆ޹���������U<}�b,x{��������*�U��e���sw\+�>���mO�e�c�����X o ��|�
�)�B��V�V�1۟�����+Vu�B]�y8��Z�Z�N,��=��b�� �$�'�-�d�:�A��ϥ�-B4��{Ҁ*uX��uz��H�i�j��l'��H;&ad`p\�NB�7�ƞ�d�7�1�|&��Q�c۲6�!��@Q�֝n�zZmX�A(Q<�EYP@��`G����H'4� \��N\%Iߛi���w��}��"~�W��j�J�K+Y�����d�~�-��p��N8�w��軚�Z� �m�>��>��&͠�R�1y�����W��4�_�7U���&|^����i_��aOL�N�A��
u�ˠ��֜p�v�	�NT
���8�L��Qo�sȭqH8�y�ɕ��D/Ɠf��y�TsMQ�����Y��.�E��M�&I[gڼ��SC��{�:��J�[w�Y;�F͕��fA����>E(��Ȏ�E�9��������ʼ�z�x�E� ��X S�T�YG�g�V�ܰU����0�3!W֖��c�ь(6=d�>F����^?�I���V�"S��x	k;G���a���۲���<N�I�	g��JXՇOrg"
?񧿦-�_��Z�+q�z�;,D�:)��ܻ���\Vٝ�h���A
�
��~7#'B���0㩁Sg���P� D���?Ts�<H,�,��c(sT��t��|�$���)���Ŕm>�f��C�Dɳ@,#>�\3d'ٿ���CL�`dx�~�
�G�%�Ob��e�����n\�'��[z��?_hn��Q�!?�|~�f,��Iy�)	�������M�dl�QV	|Iڡ�x�j���c�ҩ5�������b=Ʋ�Y��B�M�2MN�����0�)��Zt���WP��d�R��-v��ՀB��)8s�L���6��ݳ}ł}`�Rm��ǥ�?���S	�!{�,TEUˮJ9�,D�M���������u �͚�sk���ج�g_2&.����I�lx*�TT�(Q����}����*,��]Oϴ³7b���Q@��fK���,�MmH�m�U��X�D��ՠ����Ǒ.���-?O[=��s�7� �'G_�P��?���@>������� ��/���76���=�����?�@x�`X�,�e��&���m��3ZY7���3v�H�`��;�}
!n`����+�13]�R�UlP����Z��[+�-���xe��W����,&
�f予7��$�dvdt �ʪ't'�B�㰗"�.���;�����V	k�AY!�f�P@5C>i��b�,�p&��-�Y������.�{�,/L>,���즹�V�F�z]��)��I��@��k�*^AgP;�#^EX���h֎^˄\����X��y�e��5�ҿ1�Ͱr��y��0��C���Up����aju_�+E��� �)T3�AM:��/(�\�6�/;�:A�΁�e��RV�z�����+V��Sॠ�+��
��H^H.�n�����P9�T~!雞[�	�mLC�����%���#bR�	�Je�,M�$��5!T�l$h��{G��Qr� �[���v��I���|�+��?��) �O���1��~-�7�L$�b-�%�������;�w���S�ݻ�|�`1& ߕ���Bse�H�tY+翾O��_*��H�~��u���ۨnd��r^�#�� ��-�3��� ��c��:k�87������1Dl���+=@��&�H��лc���b����#~�j! zU��d
��!n�ڈ�A:�h�S�hϙ�A���f{T^�J�Y��.3L\��h�#Ҕ��C��;����Ƹn�6I/�B4Md�X�(z	����da����H��a�
�b���Rt덋�bW�y�,N]�p;���מ�(]Uk��Y�>!�^0L�[�7������ӷ�ĞX @��g6��E$��X
����%�6�����Zڱ9Q�x�|�^5!�R`H�M<�e��:��~A`���8?wz�}PD�	�G3�r���zq����VJ�}�ę#���٠�Q��0��:�K�ϯ����i�>Oc }?���=�~�c�3*�4��iZo<��d���1/�25hB�f�7Q��T1��&,��Ѐ��[�{r��I����'t�X�|��+t�{	�y��wm_� ����
_3+�� ��(Q�p�J�	9����z+>^�iT�cú<��ݍ��(.#tj��'�\���^d��TN{�3G�w����w�Ǐ.�B���F��9.���tg�G�*�����3�� @6�%ˋ�3O`��^~2�ɑuQ�I�K�5��b5u�a$�c���^���A骐@Uh(����~Z��VM��r��=��s�L�~���h�&�H΃&�����:L��Ӹ2�7vZ��'��($�G����[��F/���3�m�]?t�莦K�H\߹���\�:�~������bl�߉'I4�\ld�Q��jA��0	d��M�+��3CaS|O��̢�2��9�mܧc*`@�-;����J�d5��J��
6���XWǏ��j�sd�*���2���0���Bw��G���Ŋt�7���3�~�Τ��rɪo7�g� �VO*@��Tѭf�JNϧ�m�
�9Sq<e���	բ3ÚX��p%��1K��Z��X"����(�j��*t��ϵѵH���[n&+F�����n�XH4�� �=ˬ��@1ٝT�,W�)��]�����=�1�a�/��ƃ��E-�i��z\�|*�A`�������ܢ/������e��.��"���y^g֘ሇ��ȓ �2x���稢����Ţ����\3`T�]n��M�����g���|�B����c6(dS_Y����0EY�_yr�YJ}�ֳ6�fL��Yа��%�D��J�-s��������6�h��s��GdH��V\O�f2�� Z�����J'[@�}`���&��(�5M��4��z�'��ߙ����s{�b_��,���H�����-�	��6+!�rGǬ@��`����o��X&X�K����	T��$|Vx�WNT;�_�꽞Td�s #���EװF�|�xp�I����>[e5��\��{W�Y�G̭[�Hs��z���p�u��¤�?p���T���s��!Pm�.{����k�0����[%7�n��b��&n���h�<។6�S�ٔ�㈘��k
��xȾ�>�.�iv5�ynU��S�X�JF��4�s�pz2_OL>m���nJ�7b�\`f'�=�?�*���c�3<�6Ĺ~��0��4����yϤ���v��>��@�CCC���,��L�N7P�JE�uBŇ0F��ZL'��tf��$C擄�:��/�>B�N*��ҵ�ݫ�EqS���~N]�M���؃~��~#�{�9I^ܹy��Y¦)$�I�	�2:�����P	��w��^�w��&��pN0}�Ҙ?u�ou�j��Z�$�����p厅��E
��C,FRFe�\c�#��߯��nr��׶��j�qz����Z�2���f��c�]���,O�9������[qf��dN��$�)�r��SRI!��↫)��������#��Oq{�ì)Aʱ1�L�fkv����X�m�ȇ��3>q ��W{h�xR�řzɻ,-�w�1��CO�r���C����c�,��sC���QÅ��u��nb-���5�K��#8�=h�E��C�&C�Y�yAA� )}3Oap�x�^P�d��jv���Q%�G�MJ���� �JVv<P�O��3�C��x��4Ar��y�� �� ���᪛�	y=��}N�K@���}���M�(�Gd"�������.@�ꍑt'8o����
�;"/�!���;1�E�J-
��F}:�������K?t���@ۚ*yg���5\=����.n+�^�ӷ�ud~&��P�4V�ꬪ�����eW�G}�.��Z|�>�c<X����Z���H1��CP��-X/���]>�]R+�J�8�^Q�*^)�O,�:��s�Ver?i�g^V�6H`���G��IMl����6��9v^'zZ�x���w�N_��.#�&4� k�����/���B+�/���ݴC�.�b�Z��>�a�;�7y�O��	)�|'��6�'V�����~�y�!���+�L�O**ߪ��̊a)�S���`�<��A �Q�l}���}�I(4A����&asI�Xή�Fa��֠ ��5f ��B��n�,�R(�c����Q8Np����)�|��YX��uy�#̱ۛ��MQ�~���W��Z�o��峬��#R�΋;M=
�z=�w*c�K:��>zS\+��;!*}� �
��v��Ly/oBWI�I�=�}֦��BP�NY2u�!56�d�@��	�P�9�^%��a%p�:�D�&�v��c��c��B�#m�k  ���1O�C�F���rPSo������X��}~X��q�O]ٛq�`L5��Cn����-��#�s���^/�d�s�1�����*0Xn!D���T�?�i,W�o�릃O���uY�M#��?�{�M�(�*�8��>�g0�_���n�K����CB�Ao�pըz��L�G|��݁�i{�)�9:�^��A�F���	:7��
`҅���Bzcٱt�H2���EJ9C^_V�����
��'G\Of�\��.�-I��lH\�����݀fW�t�ͼo6���*���t2w�٬T����s�������[W<�u&C�{rr^;2ܻ�#WR,GWع�(C�^Z���;���~�ne�]{�v`Ϳ��\TR���nA�z���o�,�Y�vVZG�����IE�}��2�e՛J�85y���8�V A.~����D�n�t�\�Wi�}B;��+,3��rԔ��o�x]����� ,�w�D���@����6i\�}X���X&i �$�\~u��S�MK�nbC�����j_���*3���H���f�pM�y�-�����0��Y��r|i;��	��Aj�d���Ϥ��0�)��@A�y�9o}���2X�x1��+��a��N�:f���gxR�"�I#�#�%޾^jpt@��:�։�zǖ2/DI�Y�{C����EE��zLj��2�Jv��ۮ1���z��),��:�t�T\o־��z�!pH0�a�g�T�>q�TZ�>�^������jg<i�V��KUq�[�.��[�Q���.{G���GOLŦ���^�XC���X�qn�}���7�m��wiP�ϕ0����w��}�q�}X�c,��I�����=�іXܠ-C�Suh�{!'��T7y�g��X� L�+�|���-]��x�$�t�əT�,�cD�T����Rc[Cj�[׀�<b�[	�W��شAY���p]�� �PV�'��q�����Ǝ�^nT�Ǝ���r[[�Y��J.E�0�o[o�y!����;((b�� �#&*H
�h�f�Yg��ش��Z$�+c<]��?��Eh���TI�H�&xh�U%!��<y�^;����V:�=S���L�}A���㾔>�9U�4ug�a�~M��.�lc��ټ��.c�E6��]:�!yH��� >�l&����nC�H��*�z�1���'*�D2���
�;��-y� N̠��k�{{�,��zCݚߠ���n�{5�9A��-Ej�u������h�sy�A����&_8��8��w������BΖ�ex�`޴�R��!FZ.���/����OY���hP�{����@��n-�F��3�(J��/�S���[�[OTlNM�k����HN�9A>�E��N���}��?��1;$��H��-�&�l��zէ�)��4�L1"�'\���\��s^4��G�Fˊ�,��(jk~�}���@v��Hn%J���ˊ��[2��N�� ��@?�����4��#��7Q]�թE����$���y���,�s/9�)��ad�3k^���ITN�/�l��&6~�$���<��Ù�U �P#@��h�`���oo�ĢQnmTC��rw17�CN�s��ELNj����P WR�Ulc:�V�~F�}�4��������4R*���h%��SA@!>?xf�1��+R�"�c�%?��^g��O���:����.�p�l�悾F+{��J��PU��~�b�-���4��_L�1p�2�5��8ΪJ1�r��R�k�N9'�D���`v�^+�n4�"t�g��9u�Y,��U�|`��"�\sC�N�oM��`y�FI<���8�Wʼ�����	<)�H2��<�v��8�`E�@��0�Q>a�%������aC}ۼ-�	6ٗk,�wb�
]���� |K����XS.s������Li5���%?U
Z��d;S��;UCk7^�Ɣi��}H�za�o�:��C��̙�F�e��#O�u�{i����d�<m�O���[��ĖhԍmN� �\��v���MC�P>��c)�q�g Ą>�=�,�����M�a\�<��\8��b-׸lp��VdhG �϶<���}�Ț�MN�my�lާ�O�/�*W�7Q�z�i1ޟV�1�ƂIq�H���0�3�s�ݬ8�pB*
�#!Mb�����V����չ�WD�v�Gb�]+'���Y��0�;�mSA��ĝ��mjC޺�aL��Ҿ��e�h�K��S���N��*s�EW�z�ʿv�rm��	�0��޼����e8e�~g�<?���M���(hd��C~��Q������
��gͦ� ؕ5#�Ǉ�;�}��vY�8�ZC�m��s����L|����%x�?�6 /�#����fp$�EՏ��73���Ioj&NI+F��:#��WzB�)��+lnl�p;`5I�P�dg�NL���=��"�B�J�^Ib'������-���l�甐Z�*ߊ�HN\�f�j����;
$.�+��?��q~k��u>�&�iR�Δ�(m��I������="�#�l��ֆ℮m�8{�:�C��Mj�2���o�M0��t	
��:ϻ�D���(�&`����W�a2?_#qxBU��1{<��m�r�]6����s�>��g�D����
�����h��2�>E���҄����O7cK=&N��e�
��>M?W�f�v����Pna�-�p�Ϥ1�װn_)+ϡ��{(�_�i�%�/�;�W����3\6�W4�
$_(�Ǵ
�y��u�FwSVe���;?������7I%u��z`���� ��OFQ�>,I#+�7�^��nL�S�;xI�a�X��j�(pl��CT�^�p�-cX*;X�����Z5s�4Xp4�W�R ��%?'i�d$h��g=�D�)�����\eW�f쨍_+<�f	�#��<K�������ojDE�Dqm�O��#�N�Iϳ��S��Z{�e��w�L=<[x��mL8�x�W��)�y�m��T��ȷdHuLh�+6V͵<hg�p�(lza����S��O�;�������,2^́��I
�� 6�n#�hΉ��gWEd�5���?�0*�;�����Gtiz���:pB���0��#v�o��<K�s�],��=�OB�����Ͷ�ױ�<����Q�^�E�^P�ݦ��?�<��-
����gg��3u��ď�
\w7��k~KH��ո������.���ݢkw��<�/ ���rB�M��
|�ބ�8��7/O�	oDL&�Q;�c������y�g
x�>=������=cIy�l~TG�d5r8g�ˉ��Pv�/��$X� �l����|mC�	$�� ��K]�Dl��Ny�a �
"��sm[\�J��%�j-t����,�{[F��`���H�0����w6)��E�f#I����9��z��Se�q�솄��;:�S@�<�H�f���㰠�aH�.6ME\��"�����묒)����پ7�[z/c{�{%h!�#��z��#�[/���L�ԗ��~	��0�@�E��"%!��8˴�$h�zE�|���"l�@g�B'�¢񵗄3�M?2/���g�@E��%h�����B��\���l�&�
��8�b��<�R^�㫰ѪJ��:���B6&Q
�V%7��@���1��ܐ�ܵe��$� s�U�J��z��d<ٌ	���K��B�JM'��ΊU;����φ/�2�x�8��ܮ���8,!�������Pr�LV]��bk�T��(���g��]�?aa� s���O��ܲ��� �<�o�ԅ3��V�*�˩�/�s�ɢ�� ��h��'�H�ʩ���15�6^�v�L��r�Y��;�6���l��o{l�Q�f~>�J��.���uR=""�_.��t�jCDս�M	T�t�a�E�2SW�R�s����ˊ�z�1���!o�f��ǆ�@���13d���,=�|�{E1/����:�;�2`@�c��N�޺s�D���J6�w�B�%{_I���.TTf��e̍�{�7���"q���r�t���u,f�2�R?����y��7��e
�WM�?M�����UYL�ń���� / �@���F:u��Zx�Yc���m9�2�{�m誳^T?f��ZTGy7��ƽ$��&c��;�������MB>@��B�8�\#�i�-ɢQV�U��R�h��6sԫuR�q=I9+���E��P�(�C������D%=��t��>_<�Neӿ N�G�Y�rT�hH�TQ1�73��z��O^��C�
�B+�@�v��#CYS��MU?HJ���+~;�t4���K��){g��!�-����U�
���y<(�Q0!n���?ي���&Yф"��~�nɨ}i��:e��SB%���i$��f���X=?�+Xx����?*�h]��������_��B�XUC�S�],�g�ӏ��e��
��Q��R�xqCy6p�o��uk��/�|P��ДV�C8�j�����Beo"/��צь�Wy��7"����@(~���� ���6�B�i�J�#ʌ��1 �&�]��UI��<� ��q?��e>~�*������ܡ�@h�5��Wl�t�뽽��]uT�>��-

{�����v	�!.�ܷt�ZT��I/(U"�WŅlM�-��~�R�'�&2��+�6��5���8�ߋ���=�N6k�f���)�PbSM_i����`��eaMY,�7[�p<��������H��d�� 7�L�i��W���Z�a�9�.޹'|�V�h��-�x��P_(�li����[6u���Π�/yv�r�QVre�v��F��#be�w�?��}�����na�NyP�>�\����~hR��֭Y2Nj�/?Y^���r[U��L�t�M�	hz�3�=�k:��"�=�)M��ĄL'�#4�e�҈��Ў�q㰘�y݇�X�]�^v^+`�ȵ~�N퀊[�u���H����@N���8p����~�e(aA�A�.�K Jnx^N�(9�qgܜ(��SCnD�4{���M��̈́GHx�:_VQ�p���$�A *bR���_1��U5�0V�DAM�?�E��w���;x�ͩ�W����s��2Pg�0�;�I�p5펙6�?CKI�������e����?ѭ>�����U�����h��H���2���!~`R_����4s#&��2�:�__Ҫ諬�	Y���nx�f�n`���;�H�1c�d���@��QYY��a�y�*�qt���SqNߓ=��#�):��8v1�hјؑ�w��	���+��R-ՆGLyPؼD棢����vʶ|
�3�)@1��Z����t~��gf�5�pÚu���7`�5j�d�윻�׌�Tm�$��h@R���á��><�X��K.ǘH��P5L��K�A%��j��4���G𳬑��
-���f=r��-`�%;�U�@��\f�[�s�Aсﰙ�Z+�@�Ra��ǒ,��~:��P"ty�Ⱦ�;�����#����?�8:����V�
��&��� ���L�~�$�Q ��܍��/T���_'|�P8	T{�����:^C^&33zds}w���]�������f���7�Ӄ�D�k���/m��m���ī��3���p��vi�	����}/��&|��۽���֢�f%ʧc�=0�ao�pi[bң?~�Gr+aM��tN��4��A���Ҩd���l��[�Hb����9�#FW �A�7���k�-;ȓ̔Xh߆�aD��t./6y8�'*?�yR�nU��r'�B��_c�ݵ�p�+0���-CٚL� 7L����XMJ�^xѓ9�8�liҒ_��o:R�O�R_���Jr�)�D���?������v��MYy,�&2?u�m��-�ȇ��0�*�+f{Čr�� .m��"�WVB2M�]@���ؠ�<����"��ƒ��fc^<9�`6��K1�4c�t+{�w\g�o&X���MA�R�c���H����N��rt/���3�-6�
@ ���y!i�:TW7ܗ�hш!�N�03c�
b{�toO�����p��a�~I���y�.ԙ7�g\q�i�r�'F��\���_9�u��W�h�TI��~��9��?��'c��qS��Қ��wc&�栨�ntRRhO�h��5r"�,�'�p�x0�D���N���RON�Z��ڎh}�:S��@�
$���8+�L�t��`�m,\_�~�ӣ�����+���$���㦐�	�H���+?������n~�����oZ�E��q:omJ��>�֭xп����T��άf2��}+��S�'P���5��N��F�i���ڐ�7"x�r�:�0����}����8�'��@�j�IS6���x�x:v�a=��k��nF^XfQ�#�#θp�H���&�~�]���@.�όv�.��)��v�j	����XBd��5b�۟�����p^�2��A# ;\v�Y�����DcJYf�$������]�φ�?G�6�������"x�Ac���"���iem�-�DmZI��v�E�u˾l�nF�W���SC���(Za+�r6&#�L�a��߉���n������&����
*	�1�t'�H&ᤝ�)������2��^n����v^�_~V�o��/�Ń_tYz6�����]��X�f�@�!�%�7ds
K��ˋk���|ͺ:�y�^1���
�	e�N��/0́���p̞(���kU��u��m�m���+V�����i��ei�=��_�C±����ִ��	گ�E�@p
S^�� ����|�L6.�M�<��7�����+� ��L
k�3wQ���m�o�oRm��AD��^���J!����7���q�p?�{Ăx�ђ
�y�=����޲��77S}$XS��Ȁ~�m���d
�T�>9�+����&�^z��c�Er���f�t#�\RSȸ�Q�Z�[��k5W�Lg*�m�'m�+��*W�up�oz�7��WL�GS݌�BFHC�֣�唧3W�c6R�����m����Q�z�ܔ��,�&N��n��R�Ô�[?��G�_�������8:Mo�N
���.y ̙c]�E�����@�[�]R��ǻ���� �z��?��7��5w�-+D>� >;(�	ε ��.c��.����E��E��c	
 oǾ��EL�l8}��,�cBlʂ��(��у� ��0����tlD�{�0y/n���V��+a�,�����ӌ�F�0)oˈ9����JY�Q�<Oˀ��Li�B�kFc�4^noq��dwz�F#��E�}��H�b�S��9Y��AXLkV����t�m�pt17>ǒc)��T�`0b0?��;�Ώ0~��VR�i�z8�	���7�RT�Y���@��^��7��7������i�8{��,3�`,xs?\�����)�>H������a%�$c��(n����e�ś��կ:�"��w^�}�oNެ>9�>��5��&�m�������������h�K�ǉ�%�Y��������;@2떆2b�-t<��!�YF�]��<��[�|.��]�'8?V�{M������;�����;8n�\�n�l$��R���Ls�xO�����X��g�1�͏���o�G�~��,�p��O���!�ޯ��8��i)��).�kt������<����4�V"��aZGN�z7�  ��|(K��L����#m���s%=�=S��MV�KOް��(��g��`�`C���dMUhx322�b�a�Y�?�Ĥ@z^g>���C��:��30�E=����Z2�F�N*1xls�G+%H�mG�c�eP�ݹ�u�7���Dݟ��Z������9���=R'�~)��R�m�q���T�̵	v�4t0�c�Wi[��ϔ0��k�BR�U?�CMm�t`�a�0? ��V��4IK��lBId�eH.��P]���^5�Z��Լ<ր��?}�X��<��qsY��30�<��5���sN���<׻�����?»N騑���큢�آ"v����$?	��D�W�7�>8a�bn��ٚ9���-;awivoSnH��w~:�=!(?�,#Y�$^
kW`H�5��^��Dx 38�����ۼǤ,J��뵮��#�	��|H�ѡ�q%�&�i��;��3�L#�q�P��p�e�^r3j�N�,�F����g��h�Þl�}�K�ٞ�76+Јi�:�����Z]w�\�bҦ�)�Q�ߗc*z`��$�\N]U#V��}��E�A	�̍6�y5܉� "��.k(d�ת�_�3�n�=K�ʈ)h)�Q�l���Lf=���v��1/��S\���w�jg�����r/�O�^�X�-��gE�P�bOޕ�j:h��9xo�㙂�=e�"��I�d� C�������V%!����C�'%��H��Ƀg�"�1.R�u	U�	��Wav��&��Ɲ��9�|>����?_G�$i�r�v3�r�ҝ�=%��"9��)���Hw &��ugu��Z"�*V��ws.�彷dV��m�M��>%�Fv�n�
�Ip�X{�9u��c9y|�M˞����c��x�7�"m����?��'g�!/3gOGx�W�M�����V`�鎑H��P!�^�`>�e��n����P��!����]����`F��M��:��\����!<X�����k�;��ǽ�Zt���!��=��F��!&�?:d��.�\�Y��*x��$}�e�����������ܛ��.��{~Ny�D�uF��R�}���}UL��y�Ψ �dV�C�H������>�7�i�\熤���B�M��;?�J�]A�7;7X��ÉSr8�h`P%R�zT[��"�ѥ����@��$j\=5M�4)4.�`x��bK���G�V�Ft�rA=KV:AWQ�a '���s(�h�X�j5�7=�xz6���~�D���b �)ٿ2w��
V��^�AsC�^H�ݗ��=}X'�'.v��"xN:��ޕ������v��M��2�n��7B+/� ��'}��.B�(E؃����{xh}�2�����,�*�z�-Oϸ�"F��r���2s�ؿ�c:�.�QqN��4�--��YrCe�H?@N�%+Q��G�OF;���!�]�cpN L���}���}�.M�e����S�}�����m�)�dc�p_������љW-�1��&��E!�0��ս�a^|��mno�d%)���t��~{�JT�����c�oyq��ڑ�� 垘Fsc�Kr�L�c�nh5D��K�^� Z�s� �&P�ɇ��&w8���}�\!@�������I��	�y[(�U�k�c�20,
>��WK����� �&���(��.s��a�A�Х��q�������X��N����I!urbk͍��� p��G�U��i��6�Ff�t�?߮�'n�ęgyb��{.���f�S-�����;�L�������~)�m�N����Ń0��+�ɔ����vҌs�a�q����`3v�=)S�:��o	�|�z��1)㱟����l|�d��;�:�j��Rz�y�f�n�|��<z
��t=?势p�S�b�
��d,����r'�$�y�@5B�@Xì+N�,q��zr�8��~7�򙽭:�����`|'/�)dQ�Y��M�b�*��7u�K)d1?8�a[9�2��a��/ ���;\&l��\�OY��L�[��Y^I_�L��bg�~	@#�%���3Cn-@�7�+���OO��$3���vd��!C`z�eD1iK%�y�-���0,2/�X�a����}�t�������O���D5~%8P�������)t/G'pJ3����;��9ϥ���<ќRj�{]���&�#B���_S �	�.=�@�{����H,�3ע�H��y�Iˬ�&FSŗB�N�&����"���Õ������g���v��5.fZ�Fz��г�.�\#�Q���6�Wۇ�GڄQ�h����W�E��x��/�&����/��޸/��2�g@�"������%�Qcy�4���)d��_D�oX�-rnC�����H_d��T_��i�u�9 �V��jPL:J1;|rq��qC�-���h�Y�[����Ɗ�5Q)$J��I�s���CrOfM\�8��~V����äY��Jcy���1Ly��n�4<�Z���p^C�;�5����L�u�M�h�Q%��Y�ǏOu��-S���CN��.GQ����u���+��ST���,��ht�̑��OA����%��N-��Kp�b�l�K!��*�x�FϪ��?���y���e�+�#B!�����@�6F�]ܾr�l��Y@�mzs��M�h��-�j!2#�!���-b!�]����;���;����X;q�G�Oǁ�c.as�<����Q��DZ4�$m�ǟg .@���_x��׀��V�ٕ��,�YoRv�����l�`%l����)�	�C�Ff�������I�c�䲎���	rE�rF#�[��
WY=R�1����*6BE��q�T�H�W�y��J^��G;��u�ҩ�Y�x���*j�4�
F�5�O'bu���V���ָ�d�ޖ�R3��K�ڷ�<ݹ��H�,��-��������[_�c��gwd)H`Tw���ʦIl���x��=؃R�͌B����������3��vQ��4�sO��\Dn�< 5zBF���ٖ�&���\��3>�׮!�`5{
��žF�OL�	�ˍLlZ����s�6�[s�E�:s����"��a��g6�
��~1��f
|�݆�I�]��j���?�݆�(�{`���cu� g�%�J�|����+���3����k}ŕԛ�P�Qڈ~<`�`��х��zs�dt�d����,�BQP-�%0�g@����B�����o��hܔaQ}��,��hnQ�_&������	�?0RE���q��4��)��`��I@j.*���������Z5�����ꍬ8�/bI'M���ViD�b�Ca��-��M�8�o���������h�n�d�C�g.������ے�s�,L'�MB�ݶr �ü6���?��2.ޜ�3h�y�|ɦ�z�(�y6���'(عP�����Ы�2�nA����V�4�i[��O���1�E\�1CJf�b4��#Y�؆�)�z87BJi]�݀۾z��T��R 5 3$����G�W��4��t���,���eg��)5�`��L ���.%Sڟ�`ބ��5�85RT��m�n&z8�������q�S/��`�CQc3����|T��L~eb�q��M��	�i4�d�E�'���݈��
e�$CP��S�N�rfE,�4͝ +4V	P��2�!�{�B�1�������{Y����s5}�8_\ ��Ye���5(_�j�/ez"�*��F�ɿ`G��j!-E:�[����G��HOׅ,e�V�IM�у�/���z�i�1D������E����BؓMϵC���Eͧ8wx�6��,����t��YS���*���/�S:�B^��,��F�2���C���_�%�q����{LO�K;��!?�fm��s���K��j�n�+����9t{W�u�x���Q7��J��e4wN]���Ӧ9A���E�O]P�:�?(����4~W)jDI0�	��f{KO S��,��@٠�q��(W�ڞ�b���Sv�]��P�x�4����o�/d�d�_����T��ˊ�Ӭ���<uxC��c��)\��W�-�/P��z��+�+LR�7�ħ�6�	�d�.U
�"����w��R�F�z�} �~5az�<<��Ziw�����6
���N.C������$�2��t�A{@�o�ձ���S�k>@
1�jgJ�'1[���[�)�
���f/v�n�_y�l����c��}��3!j�}uhָ�1���ї�}	�k��Z5���*{�p�D�����WݷZ�}"*�H�v�~5�8�OH���-�)D���5�ҿ;�"����B"��'�� "Ɯ�����_U_���	���P�q.fY���Rg�ӭV��{o���0SE<;�W�4oo���g(��+�o��>w�,�>a �[���f��eY)z��|,vЭ��Ћ�v�Ck�)���h
��09
B�I��0Q��),#��s��tyF���֭�.F��3����l�QCy3k�.�a�����nP 3�7}l�7��A���?p+B-�� ɪ�	Q5���F��9��^G�^i���C��I�e�ËN7"� �����l���ŗ�%�R��;��i�?�׍�
G��tڬ	֦�gn��eg�Ǵ�,?�R�<z=[�<*�M<��Dy�l�6�D�u�i�\u�����e"	����D�YE>���`VEؾ�@&�?�FƤ7+�Spw��u�a���}��Q�����q��/�<�	߽���C��ޤv;2!>��S��`�ʞH*�$a�{Ě@��#(0n��Uz��U|U�� �Ζ��<������`�Lpn�do5>�Oz�J�uS�ge��|C�5n��L�k�4xm<�|��6,�7�^���G!�1��j������Pq�:�i����y�K�!'<�
��=V��Z�͛A�.�zd�+��ϼ�cU�\��;�B�x��ӫ%J���)�l����Z_�O�b�{M]mP�@�	>Ż���[q!~��"��ҽ�
n|=	hc|e	�پ2��*n㴙$W�Rqih�_ҷX��i9*���ϟL1�#Ig�;��NGO;
��J�j5�a���ֳ���k���̺J7J0X�!��4~y��>�B�	��z'���Qa:�J�d�Ƣ�z���sh������`3'�xK�%����c^ֳ��/�CY6��\=0���%p򚙞Ct��Ӊ�r&��}b�����'LZ�޼���<b?n��D�tЕ
.�&ٱ��u�Pq�SJ��#�˒px	!o��!�d�H�8��+-H�*-���Ͳ^qIE�x�t���Ŝ膮�/i��^��T�;���Z5�Sl�PZ��QV�h����0G�E��S��6;૊/�*���b{!�����C ��><;�CG��h����]Pg3{��IM�z� s]���So籨=2��T�l�Ibb�?e�+BI�]�K�9�v�<C��s�}��KW�n��f�W�.>����ݔ`ڦ�*�����L@�d_q����,5㤭�-�~�F�̿m�ę+�E�o�"65 �S\F�L��[�=�;̠w�ez��5Qiv��< ��i��]��O5"��ާ_��Z	=ʽ�eH5�[QE���;fm��o<!L����}�\-���IŊ���K�w77�ߵ��Y�!8h��~�ڬ�g[�\.�ݎ�Aͥrގ�C�o� *��NQ*���K]e�ۤ�~�k;��u�G6;�>��Ɩ2 ߛ�߼�,s��_��H��dڙ���qÀQ�Ea��yC�����I��������S�މS$B�B3�1������N3��,!�==���,�:&����5|,d��i!�̫�/H���,������i�c~�L;:�f����)hӹr%� �0���e y�98^��9�Қ_���x��)Y6<�q;N�Y���c���ڤfmk���A��pZ�X_��C�l��aua��oζѕ�����Y�7��B�鷜]O�����7qr�y�x`5��D��
,|.kYG��1j'�j�lݾ�9��kJ�}@]z��	\zs��u��\5���aDLF��4��ӏKli"xǸ���yH�>E�&�^|�IQb6)�σ~�!{,�9œ��ZXҘ�f��q�L�7�#����D����U��o�G2#�"�;���JV�"�Ze?� Ga��_�Y�R}?�S�[�	m��.<&<7�73	e�[�'�����1Z�ٶ��X<�O0��֥Ȓ�)E�-� lr����O]��c&$�b�E��	tDt�w��޺4��N�I'������O+���"%�6�㰜 �,?���ҷH�M�G{���ղУ����'��.���Cr"��Z�h雓�o����Z�d!���5�����3�=l ���N�)�U�U����I�O�z q�@@��͒�.��dt�H[pܹRCX_t�-)7\9���x|��t�xT���L4��t7��os+|���_�)�G�w��@�!H�>9h�4~�e�&���`N3�\ƚ��lJ��`���?���� ջ��T;S7Zb�>��.?�p,�d�O'_� ��pH;��@�����E^���F�A:����S�e�1��������E	���U^d6*XNՎ�C�PJ(e2��U3����r���ap��v�?��DdU�j��[;�b�j�{ʡ�DE/'��n���]�4k����z���|�ܦWb��O`�'���i��&��?b�~9C�����ꬰ��p���=Se����0A��^�����lc>&1
株����r�{b��تJ��I����״\ܥ�/Oj`��6�ݟR<�pT��;)�q׿,����1mudx[�;�"����༝�$Ji爿��[��=���&�D\4�G� M�;��7��c��L�r#�BJ���Fv�'��1V4ΆT��^L��9�P:nNgs�p��xeB $� j�` �y�'�j��T��x±ѐ�h��zj��S-��4gjr_CO��Yɰ �SW�#��Zz�}�Ϙ�]N���JN��!,����8H�x�Ye\Xj����ˈ�Qiu�&%�ᒘPo1�-Z��pb��o(�$D��K�p�"ԃǵ�����Y�%6JU(R��������	1Ĩv������A-!�����K1:Zs�%��dhQM��ao�";%Rz����L ����0
h�Ѽ��Yt7��t���9�m��Z��p��<��I���8q+�_�v��}o���k��ظb:����t�*}���PG1�����_G���
�ԟ�<��9ڽU�
�X<1���z�gD�b'ͮ��y��F�>)P����\,I�������2��'E1*�d�CP�!R��-&k1�,���h_BW����P���a����*l����:�]fu���h�9hj6
� "�ղ1]�L����I��������n���X�U�m?Y�Z�Jq����A�`��ܱb+�>� ����m9O?[ޣ���uO�r��B ʫ-2�ߤڮ��w7��-%�H+�'`�a���\�q��ecCMl<��m���10B5P#�{9X�V�`��eF#S�D��������Pq�n���X'U�<A��d�������Qy�
��}ީ�9��z���Kv�w��ž�!u
X�b�2J���J	�F�.�"�V� �U�u�D��Ƽ���Ru��ػ�F��n��@��|T�I%F�k���S�\���+���K+�Z����/Ь�	��ƲY��k�Tv3�
�������ug�Fw\�zw*w�2�S����>�o!����4��? �J���h���w��n�/��)Ȁ�Y�a����6�h�����uT}����!Q1�);�� 0ң��"��1���sˇb�#r��]������d�	��XB��I[A�䝵Ď<�y
a��� �QU�7`��1s��<7	)j��p2ܣh�l5�/X�܅�g�\2	�b��2����!��d�Ȧ��hl{gvA�L7�=x(}+��|�.!����̑��[8��㖪��b�HuR�_VES_�*��y$O�:c�O���$pE�:)*Bk���L��q�}�Ɲf�����ɳ� �p��tW���O���ⓠ���᝔�i��_W-C7��6+p����Z�<�'����������b�	��hA\i�D�uaoM �1p}%I8� N�sl�p;�d�Q�����BN�\`K�Ol��rÍπ��{ψ�:�+O�/C:s����
4^�>�V����V�wJ���r.h�}U���­�щ�H��+��UH�겏�.���)�L�zLͷ?�'b'V��T�8�%����6T9�	<3j�����`�[��f�V���3���Mr�^s��i�j�_'�w	5�y������v芤Xߧ������y�u�8h�p���
um�0�k�kl��$
D\�1$r�O課��Gųኝ��|�#�5w�L61��n��36W�P.�N�yn�%����ې���D���\$���y��=���9z-�m�]��#FV�������Œ�bc<�}
���g�%g��th�V,�
1�J	Y�Z���T���D6Y�e���r`��RU�B�J�Jn�ղR?�Q
�d'���T)�U�i�mڱ���r�"���_("�0U0؟�K���`7"�Hz���~�e0UOZ@�Q������r7A����k�..G�g�K��S��zª��h�����8�G�$w���*c����J뱫�M8��cKP3cy.�O�'�4�)�x���SdXΞ�i-�0x������XV�O?���y!��"�T�� y�fZ|���=�g�c�gC�ڧ��[�4��'�Z�26�W=�Q9������VY�4_��$� >׭�Pn]1-�ğd�j����M��5:��,;<al-I�?�C�P�����c,oV�y��=�V�\]6<���ܟ3X<Q���F�1���^+z�55�v�y���5���b/S��B$��n2o,I�<(ƺ�2_� ��S=X^�"�,80*����vtw�]�����[.E�.-BRH�3A��1�EeX�������WkT~�-%ͫ�iߠ߼�x�Tѩ2<����t���+i:��+^�,	i[�9��_`J�s���.�~�3	�<ta|l�;��ﾬ��.BT�z��!bvw�Z�Y�����$k�?�	�y1�3���u<�i��;{Ml'@�V��fO���d��e����F�U��9B����:���z��Yץl��S�:�)P���Tw�Ǔ@%���h*iӷ���*|���ld��6i����)6yz�P��*j��2�QA����4P�s,�Z�OF��hIxP�R!h/  d�DF�g��=��z��=�����k�6Ķ�Zz�q�?It )�Ow���G������]YR��`��Z��φ�۽��#������V"7���zD�0�x=H���զ�1Y���~ov8�����&�˧�-y5e���8"�I���Zr���)]q��n\�)hb��9�0��T�z�J��/~h�X�b�s ��p���E���(T�Hźϥ/z����֙ia��0ڋCu��7���婖1Ҹo� �r�D*��>��+�ye<�uх��R�A�Bt�{�J�j���!ɟ�USΟ��;,+��VB@l��#1�Ԗ��T� �䀏�2��!�SMx�]�;0�N����pW��j;m��4�˞E�un�6���n�g(��Ж�c�E~	EA0�0|K���^�pq\v������-*��L3�P��1c��E�0@҆�3�%�$4��
�4Γ�#n���ι f�<�FI^F@|�G �h���2�0p����5��M"țh���w�͆���Jz�X�@�vY���۫{dy���deh��c,��1�.V��Xk���.?� ��,�<�����d��Q_6��ٜh��`}L#��:&���p@���`Qb-wҿ����xdu�
z)����oE�JlA]C¸�\l��-�[u�����-V�̌t�"�jztš+�+!<	:�PY�N���E��
zG��@U�@M��t1Д�d Z�Ե�����KUC'\;`$���ݣ�/4N[�bp�#U
/�W��'3�:o��X`�>#�)�ͻ��e�*����M�U���h��p��:'�m
�u��g� p�#�3���P�������ol�Fhނh:I��܌	&�K���F����F�~�+j��C;�y���
��� 3(�8k{ۧ�*�ȴ��X��ӎ>���1�7?����D���+HZ4se�y������}�x��y�BD������]g���-��uL�%���]	��#�ht�� ��p�TL�G?Xj���]���!xF��������j	Ze�As�z{GO�o����R��FnT����6����(��D��)G� i8�Fυ"�<3����[�O��V6��Qv�Vˑ 4�S-�J���s�*
��	
�cG�r�w�~!�)�N�&漢��Ӧ��f�^�OcBiv��8*W7�H�ŰL�H04RY}���b�v1�²�v2�:���u��`,�&��x��	"���*��V�a���Q}��m�/��<2���H�d鯺�N2�a����S�I1�4��d�}7-���qk�/�S1U|�������/�-��?����%"m�?�Md�e�8�bPU��d�SA���~y��������u��C�{~��*C�	�u�8!�6��QB�8�'aד�V��I�����zn����+��Ц>�J1L�b-��UOE�O����Os�> I-)�(��&��8��^a@b7�/u:� &�)ߥ�P��&&�9�\'���x!�s1ANfB�V��,�
��UT�p�`>�)�ͩ5�������'�
%t����܄u!����J'}<�-3����M����,����DqO���L��`�=a���|\���s��[c|�RZ%#�"]��3���W�x�UCU�_�Q��X�y�E����������٨��ӿ��In����w���-�ݻ	�+�!I?⯅qRɜ���Tak��*봝xK$�UԖ`�3B�g�ً=n�fbJmFR�X�Q� �m��'K���b2v�;	�l �������m����X�AR�GO��Yq��I��a��#0�v<}��9hyg0�^ɍ]\Lm�dM>���i��
�p�w"���dU������d���xɀ�TAl�=!���^�Dг9�h����w�I*k��T������G�VS�lN�ƽ����:�ǇX>�������KQt��!=Kݝ�w\��H�q�P�=	 VG�R6�$�/T���_n&��]��eJ���)
M��@F��7�L�T�zO���oCG?|\���%���ǩ�R"�����'Vw��,��J�0�f@��&E�z.�X(�M�xj�� �{��F0)�^�ʵ����1�&��n(��	��ז�~)�ܿ�ej�������KMO*����I�[<6� �z�s�Ϝ\0�lcl�n_ii��kYc�&�1�Gj!�I� >[��9ߏ��*|maO9|�X�M;o��(E��$�|[b4��K��z��yz�FS���9&S�g���{�_�˘1��3'$S�Z`Q����B�2t�m���Ed�%�zm�F�	����ܥ`lxm��t÷]�5�%�y�tf]��n��D��~��� X����^��L�@�L��:̪h������4�<R���_S��̣m1؛��K�A���oׄw�m#d��3�+?���*�@���Z�U6�z�x.z�,jL�k�]�jy���h�9o�ۣ�"b3t����:<������ZՈ�T5)!��B����JO�p��[ZX�2�O�|�s�LR������m�������5�ԯ=(���f�e��%r��8-*��r��� ��y��A�kMM[S��f������q�K<��\Q���$>��q�/V��j/|G��_��au�a��Dy�4K���o3]�Ҭ9���
�Ϫ:f���(:�Q}�\C(��i1����:����.��#�� �tak	�g5&؆�k��qA@�o�AQf\qZ���.[�[���`w�Ug2rѭY�X���ʺ�1�bѮN^-�c[db�n=
ny>�Ъ�O�Ϛ���|ф<�q|�L�d3Њ��&p�|�cG�F=頲qNy\���_��խW��c���ƤJʅ�|wO�������m�����#���4��S�F��^a'��鞡��O�~4eܝ'eLa[��A����dO�0�#�)dơ{eG!�c���g=8S��A>��'�aG��������r�q��B�]7g;�ﻒ��Ƨ0���U������/X��=�ow���O�c�z�#U���p<�_�遲�^�x�@��m,)����YWMfn$S?'�!a�fOQ�w4J��O�nH$h�	N� 8�򿄮�vkC���q�}%���4�� <�V)T_�G���E&s#����0������_��2���<�:� jƒ��U���Qa�[4|��\N�6�n�3�5�N��}bo`(>�W��dl&|�������%�9=�A�զz�c@�7�p$����ut�q�0A��I |��ԵQ���g�{FN���
(1g}1:b4^?tTq/��jyGs+��/:"��KH��N���3��n�~�ŧG��j+�Y��E��AV��b�-�Q��\q<�-y��<�	me�U�F5ۃ!\�y��m��xaSl ��G�]��x���@�gd��5x�G�����zHc���$�G���:^�cQ�^xX�C"������0�p[�	9�H(1!N��ͻ2w����2�r�ˊCb�Y��Ҵܪ!=�%�����zŃ�S^��Z�b�w����ޖ6$d�2���e�Fv���!�ޢL�	�������5?q��;Y���U����1<ؚ�cG���{6��X���eG��ֲ*�c�G�?e-=�`��p�5U��K)�Q�}�)��R�`U��dZ0Ќ$J|�="��Q���t�M�������{"x��Ú�fj���p�2��{|�
�X�)���e���e��˒��t�D`l�W�^M��X��c����Y�gg���E� �,t;�X�i$Mٳ�w�a�z���~��}���5�Qq����b��S�-b%������F�S����/L�����>����g�FTl'��r�z�~;%�zoa{�`���>�g�>���Od�K��-n�@���J�Va�䳸��+���\�4����
��C����V��nC��n�"��^BKy��~}����_.�&=L�\�R�b�o܃#"����T�0~���$�@ѹέ+�3�k����R8 >z};.�1�P�<�N@Z�ja'��2B;@ �.�^�5°�%�t�[����]�~�
��}47��󸋇%�s�`�M������]�b�$���5�� ߔ]%���#L�-�H��I���f ������^�Y$r$�>�k��L�ԍ�5}0!봽b)&���+#�/����Pb�_�T��B�Lй�ō�����IR��{�=U��#);;�Щ!�>Yz&�G�)4������q��K�2^�\S��SMzIh���j��RE+<#K;�e!�-�g���\P���'�/���)���3��?m���:OLn؞�G��~ᙜ��O��Z���._G#�e?{bY�O,�+<]H�~�y���ZɆ]�\64~�E�tN����0�qsU�QCl\�ez�c�KT�,��e��ZW^w���e>t�=��ng~W��թ����d�@g�J�{���#"�^+鼑��D��r�3�{�1�9�x�dS��/�#�{~�"���>���娈�O�ʉ�Xj�C;d-�X3Z�b�#�!��(t� �z�J�6I �#��� ye������d���_h���;�-�-=��pq��b�vi��Wx���
-[w�mX�Kh�SC?A�q��)�U;�����m�|�ݢ�@c���'R���B��boj��ц߈�$N�e��<E	��6Z�XFO�gY�?���2zDL	�aɱ[8}Τ�#_0zu���T�i���;����ayXIX�/�M�&��z���i��0n��B��lh�ʾ$(l��8Y��g[/4|��d��7��ʾ
���k!z�<�5�jM�'˞}�x��A#c�ա����B�*LOI/���5R^l3�}�-koxr��S��<�%g�ɽI�罚�땀R�h��,v��)�nC=�9����\�U�ς�-�w�?.J	�ꨓ��K�/n�Qc@��2�.��D슊�s��̮-м�X#X� qo���+N�R[����%<Do�m�٨�����ha��
I�6n�VC�\�T0����m���_���CA�/V��?0J�"@p�9���Ae@];����^��6y�I����d�AQ�56��i�!HPcv⊬W&��U�&Բ;g=�KWA;��_K��R#������)֢�����!�ݪls2�yR��<-	�� $CI��[�%[�!آ�6&��(Sb*`�	-�n���임�(����մP�m8U2l��� �Z��w�
��:�����T�L/9�����+z7S�]؛���z�V��fߤ�� #��:0���@��z$���A�`�*߰T:k"c���[It��@'�]��:����bt.�����:RUl���d�C�y��=Hٵ��Bd��R�A�ZUH���L���Tm�@�=���h,{�JX	)���1��z	�߼O�%#��f�>�|���;KW�^��f�f�%ҥ���b�YsE����k	��x��y�te��(	G�����b��Eb ֐��������Ֆ�y�݀�8��|�f���m:)Q�y�f����:7~��'EZ%����E���6�Nh���[�n��3"'�?v��u~�0�}�q�F��*�kH,lH�\�p"L�'$�C��uɱ���W�����T$`��M B�S �J���$?�Z�&V.+J&��lS�ƅ͠��mIٽ�����i�%Tk��^z�!�mo�J�59�a1R������;d*�'��iō�!�/�mb3�x����8�z�jl���ߐsFEc�;���\W��7��>�Ձ����j�6v��׉`�� ~�o��D�iWW<�'�j�q=���|��?��tpAxV�/�c|�A(dY�b"�&\����M�@`DJ�?�T`�Hxh����E��E��Lڳ��j��C:���^"6|�rY���Ag+��pF����amt%%;�YM��yk���l��a:��~�+}��Y������/]}���a��XQ9��X�����Tn����R���P�=��4���4�*�5���ecɭ��(�__� m�n6u��R	�Ѝ�pGB@�=x�b�����w�4��q9"S ����x6�|<�>xv�Ѣ�1l��SU������l<��O��nLr�o�yS�d��x8%3�Ĝ�&�
~+y��mX�"OS��`/V�sy��mf�({&~��:��q�Hlgu�����������c���b>*�T��!�1�t�Q���(V�D\Xu���}�H��=5&���[)lgwQ):���q"�7Q�y!��&��K9�//���:zm�_��Vb?(��D�|4������F)Մ�bL��r�L���Mů�w��t� ���M2���1Xސ�7{oܣ�8�6ڞ�� �<�D��5�uJ�ĕ��q�����l�0l�]߹gF��4H�Ƈ��\�f�(�t��Hʣh�I��E��pr�΅;mS���+������H|�#����]vtDKt���dz��iWS
M�/
vIq_��/���w�.߃3hF���[�0�zX������-�v��jw��E2�|s��_��&��Wy���Щ����e�5���ňFI�p�B2�Y�؛>��ZY:��&�����^���k���-�8-�'PޚAuה�	p0��P�����[��X9�%kL1�R�
M �}Kd}a��]wJ�}�z>��1��tn�	a�α(ɳ��n[�3$��!Fq�G�U���ăC������`�Ƭ뇸}rQ��ԩѡi��p��<f|���Y%C�8#���SPp�����&MĖ%�)G��ug��T��I��8��,�46k&���P�MI��qr5��^����}S�1�S|��h�y�G��+Ω7%��w(8:��zj��l`���/D|���3�P�F�����÷��9����2�&9(q�<�k�VY�(�{|��"�Te�@ W�/N��X����T�3]er��5y#�ViUy�ۦ��C6H�9g�O�Z(�]�v�bW������%܎y�!k�NK���oٹ�(�+o�\��w���ƫ�e�P�Mg�!�㣩�[*�M��҃^�岫��SL��n0���B��1m������s���C�|^��&w�2��"�@J�-��Rq�>�j�9"��O�?�kd���f��?�4*s0���]ƾ�E�3>��܉�kn�u
Y=��g���n��x)����So�q�"!�I/b�<(����%o6LMi���W���솇�N}e�o�81>]ej+�Xu849�������{�������-��,Np�;:�+d��%�Д�]T�i��%�oj�^���E��5����������5��)�421���Q#�{Ƌ|�b"�q�m�\	��@)sm�FQ8.<�:4^E�]i�`O�C��L�me:�[CZ���lc�ِ�����Zj�V2<��e�#*cwH:��!aq��GX5��+~����N0
I}���r���5�)u�!��l������s����G���ߊ�����?qźy[����8��c�ܙ�K�T5n���W)9hGy�N�8�Q�2�,4D����ѭ������}�<N�M#����*p%u� �D5p�:{:Q�:&����858��(A?zL�y��<�F�;s���������Y�i��}BYuN��X�v� ��4d�/,�H'��s\��G.D�x�a���a.��<{���he�Si|*h�`q���w�������gV<�i���1���<���7S�����G���$ъ�Ă���)�L吧����[l]�П�N+�ع6�Ab8� w��Y�oh�$O��nSF�/Dւy�����(,2���$ϗ7�Y�����0N��(�ǒ��1�F����c��mf �{(�1��)��U 灟�UJ��3�����;))�a^I.!&������4j��[��ǚ=�l�[%1鄩�宷=ڇ2xq�Q��bY��p,x��^��,f����i�eJj֊wc��0�x�&����b���ŷ��M�"5�=[z9L㩉b�\�y���1�C>	�C$Sl�<X�#�2y���,�~�pty��*�b�~�2��x��Օ��sLBt�dE��S}�#�L�������X^��n�~��������bT�7��ݯ��U�7�H3�V!��g��x���8��&S>C�ﳠ��q,1�������r7?0d��Ք�A�U]=�YZ�#�$�!t�0bㅘ����֎<�*?��],��i���\LK8jY�?k����<�z�9`s*Ͼ]L�JE=�OƇ��b;Y&}� O�I�>���/�N��	�����W۔�ǘ�t�NJ@���E�qJ}�!��[�CH���&Dq-ߐ�I$c��Q���p��n��S���#+V�jʧ�,�����R��s�#�O�	�/��j�oQʛA�����V��C�V�?���ĻT��m>�ܨ���6T42ɔؒP�B-� ��$���,����IXX1�f$�i�ӈQ(ߪ4��
�:�']�����~>d~EQ�v��%��=���A�!ֹ�v��ApH���/�YT��B"8�%�t�y<�!Ԧl,�嘛�\-��)�#�b�{�PM8�N�\��"[4Nl:���j��u<e�pɧQ��,�TY�J4�p�9�������pW ����"1�Sؘ2z��x�i�-6��%P�'�!qhTV���`1�B�3�a.�T6w�F��*�����$�������3�n&�e"�Ѱy���.D�QlE��Do�$�+FSYl�l������{���?�\K�_�ǈ������x}_�a�ܡq���p������hQ]BE'��~m.HCI_р$��s��q
;��z?& �=F�DD:�E*4�@�!�Y����,l��>&�+yTjnD��hP�����˒��F̞���R��M��0��p2�r��c��L��6��zɤ�-e��<���6�XPnY�A�⼣���g _���9)��	�Y��L�X��6����,I��q����&�6�ɉKd�e����l|��U<�ѕ�95��Eu��V~?/�9'��i�3�S�%C6,o�I���OP�X�]�_�8��_��>"��:�z"T����)����j 8�E��F��0�	�k���(�3/j,b����脶B�"�>҈���T����
���mpd���m: l��K&Ԭ(���w��I�Q�����<v�d���^���\�1M��b +	6J��M-��=p�F�-��8�[q�o,�{+)!�"�2
�j6�Ó7�6�Ǩ�J�z�K�n}�*�������:����U�j��Х�z�0 ������X�r��#�X�u����j
0���G��MX;�8]Q��6��f'@B����K��ӣ���� ��>b�uH>�*��M���(VEri���}�f�!?3������;G2W"(<"�#5J�N�����$�W�Y.���҂�2LĦ>}��)	��� aij]�5�lW�'\�RD|�\Ra4u��Vi�"u��2P%]�ҭ��~fzp	}/0�&�N}�+5����k����ƸD�(ϐ{��/Kk[�p�����J�j��ǒ>qJ-O)^�,v���>uR��,�y1��[��T��4C`�v���<��8٠A��r;��"��3�_B�E4M迁4��Bs�e}���=9��Ú�}h2�=��-�Y�'gϣ!�Do"��(�Zu�0�1k��7fI��6����SL��	��޲�^ ��utV�m�?{阩k��avq����}���a���ABb�������YDD�΁Fj'�o� V��XT��n���T.;(:ti���5��|������;#�&����s�|��G`X�~!8�Q��`9Z�����=*m|���Hn�^3�K�� J��[e�8�Lav�L'���FBNMm�2w�J�V��JLi�髽���~�ibH Ff  Y��GZ#Q�K�����:�#��xS�75��JV���)���Z���	|	�d�������?�G��	�Mx)����V����"'Z��>{]���Qy��r�#
u��߾�_�{��t	�����<:Tp.�P���#�(��m��k��{�|�]oza�Tņ_��~��
&V	J��&$E0�;�>�Lx��RH�d�Q���q��	q�5��	>ˬ�ұ�H���;a˯݁���G��'M/0/l�'%��g�%�i��#���P����k��\�w�ף��Y����lQw��>��P��},V�L����^�.���	���
8 ]lI��Ɉ�!���6yy���u:�3�&�K�~~o��T�8���nkF<���������!�_��Z�4":���d�:磉�������ڸ�^���o<�v�ܪ�@�c�G�}r�CL�!�X(Y{����nJAɠ��h68�WL� 8q�t��bX���Ȑt�t:kvf
���G���˄��F>���1��G�^+�K�����G�N`G=`���Wz#^�(^z�H�_Fu�.���S �y�5�|���%��̅�˨��b�Qġ���eH�/�u b��y�c~�����<R���/s?5�m�b||�咣�&s_��O�Y%��Y5Q��6�^�mFq���b����;��!$7fy�q��w�3�X��Ŕ;�^�P'O�r�W�8R�^��9��#�E3��J�!Dc����!y�1��+�;�	�!�wVy�����s�E�UmF���ұ�w?��G���;$g��\�-�� �W�U�#7,֗��oYf���c���`�Ӗ�F;���D��T���Ou��w����j��Nެ� ��9f�ls��X�'x��V�Ⱥ��
������6�(h�v�
�#�"����5|������ߚ�9����F�����i�~�8ha� �}�3�ſ�f�w��7��Cw�!|�I}����_���l��j�����r�HÎb��N$Y�&ܣ��87��VU:J���lV�9�¹�n�a{� 򄴽��9��DWr ;��M9�������(�VC_s��������n۠�-����-��PQ��6	�92�YX=�Cf!_4�K\��|.����gB�K�7����uAI�O������O��L��y�|O�j������mc�޹f�<��XN�b��7މ-��E�\y��Y����3W��<�ù[�(�]/b��I�Y����KM����9@d����8��M3~�=�n��' 	7�B�d� ��X�����=6���M�1��p��A\m�E_F���(v����M(�B�#:����^�.��2����䔳�+^�lN�+㱷Y�3���됋��� k�����a6��۹I���� b��%�[r��z�xh���w�j��؇/�t�}Q�����{܈�pIe�8�MK�Jtïj��m�� ���#� �4 ��gt0�5��4�(�h�8��+�؜���u���J�̢�i����ɧ`~Oa�����5�-4w���3�F�*�u:�^%aÖ�6���)g�`�[5f���$ew8��x~}����rI�Ȥ(,S�%�y�uh�U�)�&��:*1�S��Fr����֮?k+�UE�c�� ut�b:�k)���B 8�$�p�̾;х(R�XA�Mo�$V�m��ʈ\���a/T6�K�T}�b/G����Q���>�{�֗T��IQ�)F���3ág	�o��E(�,D=��k[�P��%�ڙ����6� #O���n ��.���p�~]�����N�ݧ��Th�D �p�����Џ��G��nP|�FR`�I&m|��|
6F[����C˞�JF��[�&g�q��E{>�o-�d�s�	��Cc�"�>ҥ�(����.��+�ă�}湌��� ����#�{vW�W�Y�6 #��
�%�O��9�@,9���m��tr@Mg���U濛O��D���0↠��%DZc�?��2E⳵�c�οv�>Q�]������8R?	sedm��Nf�5���8�=C;Px]�(�(�N'�������Q�|��b�|�\�:�Wq�YqCڲD*Z���:��w�f��T�X]����}%����j��7�2���s�k�K�;���.Bliϯ;�� S}�&^�;Y?1E�Y?���S�7H��8pq�g�i-�ԁ$x4������1�m�'�����e����g����mg��K��F�Fg���/�.@������]���ǹ�uw�a�%*ŏ`�)ݭ,�-E��HXW%c��j<�W�{Ԉ�Į��R�nckpb���������BZ�sd,[�~F�e-�r�#����|)��2RؗG�r��{:~���A��C�"x�8^�������<85ە�S�T��0����+��ө���	�-��%Pz�A$�Jv�n��q�#��<����0��>��s)������j�j�a���8,NH���2����7(�o�*�ff�4�����Ń�Ў�hbN�hGL�u���^'u�]��m���5��]�9ϵz�Է=}�6��__��ǈ���E6i���
nBF�S��Y��d�88���CE1�(�N�H)�^�S�����#�)�~~oϘTv��R-�߲�+���&*��z-�n���bf�*�ޚ���	o��ގbɳ���&�R@�%�u�+���Yv�O��oN�ָ�ۥ$����B{���u�Hn1���\ =^�KD�x*���g�dT��z�ΐz#�Ru�ʗsMA���*�����Vm����#	�0���/8m-��w穲��\U`�2ź�BP���\�y��	�i��q ��KS/G<W,��1VE(v��Uw�ѝHdN��7�����i�H-�
���\������q�%q*m�eV(Ո�KBĈ���ڃ1�˼��Tr��j�W���ZG���9�	��
���L�{����eh�@U�%O Mr�ǟCu�M]�������2'fi�Z��B;0�7�d��' �)|��Y�^Y��Q�FDV����p�e7�:8�|� ��Xh���2��n����;cU�0�Җ%+���l��)`$c��:���<�% Sw/^b��p5e�:"�����v��Cޙn��s9��/م��;4PO�=������F�2�^�>�kib��S
�ƒp\��κ�n�KW�\m0X�B*5'b����0���;�a��6�#��H��2R�)����F�Qq�8��I[�E��QY����;k�����yj	��;�.WCDA��]Z[Tٕ�͢BD\�k�Ug���^Ѫ.řl��hZEH����x�(�(��p��4Ԭ�;8vJ�`lI�0@,�YG�SHO���r�Lq/!6��>%�Yn+o�v�toZ�̕�2;�C�������(I^��J�+pj#�#@�4/U��f9l4��^l"�	"|����2�ܪ�}[��sd#L���_~`4�3���k��cd�S����w��V���o���誗7��bn;I��܇^�^����>�	1���N�e���j5�rvDC�]�s��4B�~i�A԰������[��#a�LpxQH�/w�d8C��i�6�^?İ&I����C��������a�N��[��o	�	ɺ&�&�m��5��?��_4��V8ò^��{���
N��L_�|�M���>@��=,���������c̓�ҳ�{�B�~��<-G�"�Yn0~�y�!
��������E��wX��ڥ�Nor)<ފz�Y��j�nW�#����J�&�e��\��'&���=��x�jT㗴zwQ�z�o;g����[��U2�l��*�{���1�5��^w}��<XJ������z��˸J�J2m��o����Dx�.����d�I_��-?xt�Z0�'�����U�G�\���Qai_V@��A9Y�):U���L�z�]�g�V���z>�'�7L6|�qE��.��5��f��IeǮB�<nKl�Q��^��#gtS����ɁmΙ�ؾ������dk��.��a����U�e˿��G]�_�ЛU՛Cb̆k)�!���C5�,C���D�U#�7������ X;)Z��,�lَ8<aM�!� �(؜��0)g�@��wR��bOܼ�|�W�V�cXd�,e<��(r�6�⛞�( �L�n�@���!�����[Ի��Id���(���t
�L�,�<�+h�. �O[7uY��o^;��3l��V8�q�������3��u�˰U%UO�Y��F�N(]�����#�YB��MI�#��XH!Ya�bg����ec^/SV�5���^e����{���<M	���N͌�I�������P���ޖd q̼��Vh'�/VE栊Y��}L��ع�ā;�P�(�����Ihܑ�zf]d!����>�;�c���ɲ>�㋍̍pN��V�Mm	���r�_�H����LA��^���ᆰt���y-Y3t��b`��"�2S����u0���-�)H+�t��,���0j�I��~�֡]BD/^�\9�8�Oes�2\'�n:��a�K�"��L���9ۇa���n�u���T���6�'�����=���|f�7��AOh-���1��ɂ�na[����K^-���L��bN'�Q����B�`�dz�����e��Ң��������sػ�K�z��g��İ�?w��<�7IOt]�0��1�mIO���$�6˸d6���k�S����0���aFE� h�����g�b�osW��������TR�lt�^%U�8��,�����4 ؏h�G�S	�Q[��|�_t�XڒD|u��ޡ�A<�mw[�� >�/p�U1��J�3	: ��(Id�GYr0�bW�ک��ϥ}WQC9�����LJdt�N]D[�Y�da�`�EH������㗲�B=L�o��=
 k/�V���oj�_G-+]�0X~�F����e�[��p��J˹��Pv�C��.6N����X�#���a]+[ف57h[�S,BP��mS��/�JN�����B�#6a�H��\EC��F���Aڗ�Qu�oIO�����y�����s�/��H�7Ӎ��x�ϙH�#M5Ry\���ʥN��S���
'��U϶�yL����yr='�m�d����w�Ķjpo⎠�D��򏖧��ԫT4L�)���!x��E���PK�m�X�#�0]�Ӷ�����KoS!!�Bˮ���9@5�=H=o5{7�n���˸����*�B,�zy{���en���de�[��_�
�Y���Іڇ.g�����bL(��A�N���!��-�=��w| ��y����8 ��K�Ӂ;����U�5 ��j4�g�����ߞ���ǋ�a#��V[Ui̢�cI�Gl�o��P>��x�UX����'���!�����t���O8�B�����u���oh���A3��s�*���U��":PK,��@/�X����QBz��R����)LD1[Aj#+�ՇxJ�#��΁��[��n}:�蕭3�y�g��foy������w8#��j�DGt�wa�)|�#it��w���ë5 =�wl�.K��`L@Wqo���{oI5��Ğ�I�z9�d�N�0�#&է�Dw�r�JW���S_v��;���M�(����\]H����xZ�{�t���ռ���7)��R���!"�R�����~#n&Sǐ˨g��*�*��b>Ô��\*�^�������9ls;U����@X+��6RO2C��f��'EE�]�w��q'�YԤRQydٙ_��$�7?c�xm���s���oU�C��hp(#��4�?bS�*�-�V4�߆oI_��#�pS�^jAL��iY�^�w,����ڹ�[ʧx_�~��suE�>�0. m�H�e��\F �2��o=$�3�Q���"!-F��o�[���i�G?�Q���L4�E%��4���� �������"�C�ϊ;ol��sfL�n����0���^;��-v���$a�hR�@�9OR�.�˖�Ȓ����-a���NC&oz�6*�V�;���?���r�֙�{��	�t�C��^#���B����`{��:฻�9MU�;bRbP���4����dm�7���Q�����KrR�X��7��wm�y��3�K���qW⪰��
&���q��wj��;\�&d^�F�b���8qavN�M�b��X���y<���U�7��ˠE<��Q����Qj�6�Q������L߄�ө4�0�dŋ8a��5VK�	@VA�L����A��V��a�)�17��N�W5�^�L`�Y4u9�����#+gz���%�T��d"����Y��5.�j��IYB����{��r��J1f�(�/�Z�A
�W"g<G~|9�=R���h�T{�&��Ǽ~�J�	ۤ���a�`I7"g8���P2�i�Y�>6qlqZQ4<vu[tۺ��<a��u@��m���-���������rɎd�w&�z9?�䑽3O�Q��05Ȳ��S��h�g��<D�
n��|ex+QR��Y�f�?�.�ˋ�)�Q��i,���NU�����}��#���vq���|�����8�y�1��p |��G"&ߺx"ĝ� cgh,�ӧ������
C1í,�����;����dh縉.m)���"uF������K�u뜳K�3i�Y��Έ��d ��G��N����u��p�k�ԛ��vXSAհh��[��<5S��^g��� d���|MO�G�}���x2�_�!�f�)�u�:���H������)�,�N���*�?�J��X��M�Uj3�(jW�
H4t����:ɾČ�D{����=l�:*�_����k���ɵte$u,����HW��i�Q��5-�D�<�����sʨ�'�=+Z�]}R�t�(�x��n �e��Z��*Mh�Y#�
v9%�#�w���M9r�e=�,�T�WXR�I�yݦ�vmk������i�^�`I6b��[��Vj0*�c��I��d1�n���;��y���q�p���_�g�Ո�����{�7���B��S/����;�R!�f>u�����F��6v��Wq6��Q�٢�Mi��I��y�����ql`����~E���C:��_Z��b���|>��Sڄx��|_�2��y�T?"��)M�����F"��G~�ii�������-m���	9�,Z��afrPƾY2�ʢ��ぽnǢ�ӳMP�ݴk��\��p�}������-���
��FX�QA�:U��)K�&���~�����+��H�9�}p"������_9���<g+����<>�`���η��~�@C�v*�U����{�<�Ǥ3r�u�Ii���!Ά��5cD�pŸ��{Be*�T��.�`tk���q����+�!�"��Һ:c�dI��wd�AD�ŸIʛ��̒�����$A���#aJf`��y�7Ո�����r8Ω���yC�BA�ZƲ�%�IZ�ʣd�k˝�p�Q�x(���4�h͑(,n>J�s���Ѳ����$r��r�����EK/������ӄ��AMF����⭇s�t�(�E�yc�G��^`<D������\qw��2�:��OCF���Vv�ށ����_����OϘ�#�wh%8~���K%��#�կb�i��GL<᚞�)�4����_g���D�D��'� ����	��q�0�s�5�5Q����0�q>���=T|���.��{���T�~��6%���q��O*�a�bR�4?lVfq�u���k��Idϸ�9��
EWKR���r
H`�ds��NM�#zwOSdP;K�D6����\�F.�Z�8Y��Ĳ�����²��RlN�<�,�*�%o��3�B��� �p������n�N;�������h rM-�n����).,�hRعf��8Rc��;� #��&Y��c
��?f�Р�i��(n�J�:��Az'�]��6������$����0ttt�l#�E�����USj��Ǿ�,ΐ
�4���:Y�b*���6�a�)h��l�p�vnT��;̚�����J1�յ�r.#؟�A�y���Qx�Ho�N�G��� d�����-~���	U7�mD(�sh+�2�Io���wJ��e��`��?l���Wj,����'�%DzR3���?��5Ӿ�؉p"üs�If[�hǨ6������3I���%�� HZ9ݸ���Ci%� �s��x��wPn��XQ��B0�� Q`(XQYǜvT)�/�O��:;�q�4���j�9ħ��n�e��u�w�t�m34�C�ghv��E������	s�<�ɓ��'��`v���ׄjk�/�-��Mƻ�X����e��3Ü1�o���e	�\��Aݍ�ʪ��pi�W[U9	��]�U�5
���{��.;9y.���K$au����j��׾��ڒ�Y�>���ϻU2��#z5U�$}v�I�S��J>0�D
[���ߓ�Z&� ��� �-/�Q�(�ƻ��Rv�\��gt2zS~�X����kD��\�p޵�@lZT�N�H�v��e����.dJ�����O[-����9<#�@����M�-�Է}U�T�� �/ָU8i�4��h?�`��4�(2�R���`��UǦ��ru��Kܛt=}sf&ֵL��# ��g�oģ/�ۧ��Hy����(��x����_fg*��JIt-y�s/n������g���e�@�h� ��$MW\�iY¤�4U�-�������Fw��$�K\g�Twfd�_�xE��-;`�O<�̈xp�pt%mC�??���+f���mc��Q�ϵFt��v'����ӿ�c�n�|�ȞFPY&>�?2��Q�.�ͷ��3p�{98J��U�4i����Д~�{В��U�݆���y�Q(�j�t�)p��:Nw�� 1m[��2p� Ae�����eWo0�K`��v����k�+�EXw�����V�?VQ�{̓�֎u�(Ϩ�7��w*�)���7d�A{��zW�̾s��"����2��,�WYk^��`�8� ��h�k�{�͜�z�1t���n��<�a,%�Ѭ���2�]:(�^�4��β�#�6���bMU�y���1I ���#a����|���{],���VC�0���$h۵��9��]��B9�#�"��b�7�[�jDy�]�s]��l��)��&�RmmX��OD���ۄ/&di�v���C5ҁ,+f��������yS�6)}
׺����7ۇ%jY�L��?��/� j�j�l	<���W9�-�ʞ������[�O�u�xb����ݞ�Zj�ǲ����=��GKq�i[��TI�����4�p{eW�������3�c4v(��a���ڋ�$�}K/�j"�����zq��@�X��z��J+H�����(x�鑶K.���s��P��8@&����ϼ�l��!�_ь�����i:�p�@�����7�~I�l��r�-�}_Bw��eˆIi�Dm��J�Ut诈	�Y��t�:�����2����!
%����\���l����+��O�{;Tgpp�����1�LR�;Z�J[�+�W�i��+�}�t����:H�����C#yzA��oK�����L�����~I�5�Q	�#��9W̘�{��#H��l�� �88hX��_����j�>Wr�V��{3��ے�-0Ǆ�z�u���� ���O�#G��g��oY�Ï޴[���9��T�З��6����S�A�9�z5T���7�?Q2(�����]��4����p�p_z�٪>D�fz1#�S��P�S��Ő��Mr��J�Z
&�Z��?Е��bg�@֭zYm�ŏ���k��]Bc�@2K{wd����֙�I�b�荸��ĊI֯�͎�ۑz�S	�Ŧ��`>f����P�r�gTw��L�R.Y������]�V����9Blz2C��:���">�Q�4�׺A�+����9�j��q��Y0^�/�
l���>tAh�&W��)4h-��]|e�Z�[,,W�\��,Rl�Ģr�ZBw#�f� �]N���!̼�|	"�0�KD:RZ�0����V��Y&=����b��D_klbI��~��U��S��ي��q?Q��q"V�In��j�X�4[1�Տ���ܑ��j�'���ͭ/D����2]$�G��������Y}���(����zI�v���Mľ�X��:wU~`Yӗ���L�]�{,<��|H�-y��?� �FӇ��ũb�Ƅ�|,B�>�*@������iW�&>5���ǒ` �d�����,��X�)F1�쟯扐5Fl���Rt�r����^�i֐�\"*���:�M��K�B<�uvi�����9V���N�r�d�Fƴ�j̳Ny����<Ă���Kk�������W����D�� ��(לЖtB��Fa�?�@��C�@��3Brc(뜍y����O�lY��K�M)[x�D ��>@�i�}���Z��@s�M)k%s#���l3��I����lm=W������l�=oP���߼'q�mN��jD��t�J߹���S�����J�`:����x�����Z�Ÿ?�h�4�l�`��1��n)#v��(�CxY'G�BLx74�FW� w��\c��.[��6�q������Oa���Peq�7נ�"�Ղl�:���6�d�竀���4�� �)�av��Fq��,���U�=�=���ɴ�$�􊦛�uܝ�([4��7�ޟ�h��.h��V� ��Ԇ�B��wy���d:��xf���c�a'��݆p�Eݴ�9IGO- ��]��W���Wn6u?vEU�Ք�����,wNn�*4�8��'Z�5��$�˭b�4�A������:4�*6�N΋'��ė����>Ϣ�wުx�A;�W�VI=�o��Od������a*p%�?v�/��f!����@pi \��S���fiD4���������P�%�Ε6b}#��Y��#�t����wAg�e�Ny���@WB�[{]�K2n���	������]g�87��
�H���W��4!�'CM��Ch��Wp��Vm���Y*��	���e��S���o�3��:0Ԙk�0�i��K7��8;����.S5�O(�b]�QJ( c�u����	��&��*���ɺ���X��[��\�e>G�i��+z1�t�Q�,6&����0��H��I>>:)�C�օC�p-A 4����	���S�%x�=������A��'xk�샓R��j^�����j����3I{�Og�q�X`�9��ҽ�j�ܖ'(G���?����K�B6�A��d8x�7���[��F��m�nfM��}R��P6�����p� ?�!��*��%#d��A���� �+2�wS��Eӂ�m4�:��J>M���8� ���-v��:�v�L8k�����{�qve��k��ʕM@���0��s�b%=��i#��H,
HE6����h(��Zr䛦��x�R�DL0��- }^/~�]��Js�bjY��4X����^: x�4��}O)kR5!Ns	��W��FG�	����Q�i�b�W���}S��꛽�^�>:V�'wiX!��*ӆ�*hv��{e_G+�5���L0���ܩz-jJ������q�[s�W�6ڿ��6��Nm�[�D���$x���	��'�Y��]r�{@ U	��!U���!�T��GՆ㌄̲y�mǄc�a[:����������i��2�6p������7E�g��}a��a�G.��C}�2	�É���;z�1�H�涍l��Ɛ�X-\�*��;����qT���2����IX�_h�6ŲN�y׌�}i4�>��}nieD���ok!
<��)ő���J�����R^\���t�,��ce򿱡ك�%ǁ��2.�i����-��0_i�­| fA9f�0�x�EB�3*6n���f1������Z�6m�:7l��N��_ɬ�m*,��'��1Ƌ���+�U��o%'?�S�e�Ω"]�.s�D�v�Y��a\����ӑ*nϩ��K+)?�� {��8h�'S�	�=��ۖg�v��9{�r�r�����є���r�x��~z�eDUi��a�)�9�nh��� �����������<{�O��N9���	�i�d"�2r7�]£�bi�}��Q���2ʜ�;�a��GŢ��ǁF-������]�> '厓�|[���t F�k9_���xe��5{����U��S7Nb�R@f�>V��9���:��;���x�X�duY�@��&����
D��!\�n�$W9"��ׅ'�D�G�]U�y��(��6��c-�/�T��?m�yۥ�h� }[6��&�df<%$�8��~vp0�)�:]
��Z28W�����-t�!���|�XB]��6�n-�4�|e��|�h�A���8N-[,�!E'��G|�ʚ��	3f���?�����_���P3���ZZA)��dw�����p̄͜��m��:+��G���JQ�z���H�����	� ��cqk��{$$2��@�͟�! bL�{ݐ;�اr�X:`�8]ϖ��M�lS�� n����{\Qس�\~�����v�L
HE����$�d��:*��+b{�P�����6����U�K(�)[�� lN�8��{V8l�=��X!�V"�=��7r�Ύņ*�Z��},sSmqt�	w£Ȩ���iR���r�D�s���~����c��nK�V���sx��WR�L���(B|5S�[k�\�$�Ԑy|e��]mE�=�v�G�ۺ�%Cj�&@H4^��y2k���2������>j\�/a��g�hR�pڛ��먮�8��m��r�]*ϡ�NK��H �Z@f�i �3�Y6܌���ٽ��٦:��}�^�� 򴳸l?/��[ed-�I���8�G��P�˩FO��i��Z,�[�U��W ��nG�dXl{�����-p7�B��
x"e_����>��o� �i���8�Iɟ�����'<1{ԭ��	�1��@i
��B�]�_����<o�;��b�mR�>��_�ͫ�)6�Qpr��^��+�A�����y-A����4Ps����Q�J�\K��pZ��~�2����&h�4�����.�C��x������w��2� �2��ڹv�����&�
��o.�F�G���+|=S������u�))��{|R�;��$^6:d9�4���KIp2��[�����Q
�2�F}�`p_�e�ms�����c��[�����M�ҟ国��Pmf �u둸��,U�'H2R�t�,��	���AFPx�m�i�$�{�)��{�5!j�ӎ��?-"�9��{�x�ԙrUX6k� װ���˫h��$ac���kK>�GԨP���S�1�0�����~V��q;H��;���<�������,���h�Х\�pN�����G���@xۄm->n=�%�2�UPh�+�r�IT��܉8�ˇ<���{�iG�:  AI���)�.9�v�=�GX�aY�*f�eY_E�q�}pz�������>.Θ�́���FI�����Gm��=��<�%�Tõ*��8'��<m��m�D��ܸ��w���$E��)���`!� ��>`٠_���f�k�bqs�S�Y������M���P-z�첼���!�?�v.� r��7 䙷B&�kGO�S��J����ݚAE���l�v�c���ҟ�7�G�]��V8�[�su�Q�
����A4ii"��J-`;!����ԩИ *�n|&�9.6	���|�g�9CRws���&��*�'kHCb�mr4Ir'1_�ʦ�m2U�/�7x�K����� �r�ٝT-��5X��oҟ��9���-&�j��� ��Ð��ɮ4BN�g����Ϭ���'������-({�ik짝�s�����\
@�&�t0��6�6�^�=4�7J��i��1�?a��tF���l�ǣ�F��3ʦ?�"
����D|��|�BwM�C���K�s�U���Y#':
(�%N�@��c��* �3�M��j�&���HI,T��F��l�S��4R�j)F�Yة�(�!t0-�SR>$���S�Nz��a�Y���>H	)��9�5=�_j��F&"�/�l���~���4�[�uL /�֌����!j"�8\�8�[�����Flf�?�x�F�oa(q.#�,h_���~2���j�f�Z��I���U�S�;w<�&�Нs*sO&����*�x� ���p�`@j[r*�˻c�������Z��*��������I����;�=�r��r]�p�eq���Ţ�	���%Où���8΅�;��(�d��l���
�t�������~5���k���A
?��K�S�Μ�㟏���h#uF��O�.�;Z�A�;��H7즊S�����;K�^do~	W蓣�j��	~JNX=n�jgZ������1��G�?	�*�u�l�uU�Ƿa�Ԅb�\�q[
�UU�t���Q�"Bzr��>�M����"��P1
�E:��t�wsbT�n5zVu�Y�ހ�,�n��� F�Юn5@ٻ��Ii�N6|���vlڧ�����[5�J`�s�V��*	p�ų]z��^އ��/���V�ӎacM2�>;�h���~x�DZ��;$KP���x 
P����0G��0�����ۣ0�>Gl�(��u�,+��hB�>r*6��2�5w�EO��[�{"G��8���J �q;VW�(�r!��0ޒ�E$��nLH+�[q��߭E��%1�*'�+��y���1��w�E�K��+�x�s���ſv�>Y8�)��R�f�,=g)��R��@7�o���#-	���99M��#[���J��a���d�����A�w���E7B��61D �����1A�����N0��Y�j��h��F�>��0���K�х69��N��Bu[u�T�8���r��`I]�<_���9'�h��ǜ,���@��g�j���Z���`[�Ҽ�]h�g�W�0*�}b'�\�a!���{�(#XD�m��`͝���&�m8���f@ǀ�H����.�mOi��I ���rJ��w��~o�LԲ\�v��z����Rw.�����ZR�p�����jl&�t+\�'�1�I>���^~>�
-v���֗b5j)!z;� Җ��\�]�m���g��T�>�����o����<�_�&�v��x����L4٦.�G7�(�^wD}�#a`��C���Iʕ~Q6_�A��33��&H�Q\�0er<��1x:��x>�����s�$��3ev��1�iLys�Jvs1dS�Ӝ��KPmy`C���AH~�α��T�w�����E��-���(%�.��P�J�Rp�����%��,h��1��}#hяL6��O�>E���<�H2k^h~ۓ]��ԳF��>�S<7`��A����n>]�GoE�r(��]�\ �?�ݬ���=�`0�]T�B<}�����8���ּ}2�4�{�Dw�A��y��n��A52��9	�:U9Xn�,ܮ.�CW�(��.��jO��Ґ��,�(ى��lF��5�Rʷ�n]/#����v总83����8����G����"�������S? �6��&�@4겫�T�-��n���8� �:��|k�tB��p˹�]6�yA���V0�� e�}D8.�ud�_����ck:�t����ch;�ӯo�����a�t�=akx��j�m=~�������-����	P)�~�$�r'�mG��?���(���O1蠞�A�F�>��]�"~v�bb'�\�5k��L2�q~�j�.��{�v�5{ML؎����o��As��Q0l��P��n���es��
��Ρz�j��-�v��䳙��T������eNrLo��,�q���1��IP�كR�+�s�9F���Q9R��Y	���i9���buM�'�5��c�22`�u|f��	�)�O��KM����X���R	F�0YsBa����7�Ĕc�(G�.cZ�X���fm6`e��0\�Q���)G����>l����|���)�r��P��?�`ru�����K˜����W��j�n�ݞ_"���l����)���M�<�.��B�Ͻ%^��0�H��Ü��� �T�3�x{�I�.n�P��	 ��j0i�AŔ�	��G������^Vn@�q�)��G�0��k
��٨ɴ���'I�˳T����v	�P��M�C+s���	����!� "Z9��qh������w\�mwa{���c7�4$T��O���i�%� 7}��".�W!�����O]�����Z����aK�)m[�5�̘u> .�<�j�%m���Ǌ~��w5F���?6�i���F���'�{��ꎿ.*5OK1�j�2�T�y7�g�N?L�MÁ:V³����
'�D杶~����P&SY�[@��&���!ث"�F�T��C��qm�����z���R����e�aW�H�7�<�����v�.'�����{c���gj��`m�<��`%4��2�"a�,�^O&�Wt#g�㐔�#�Fh��Ι~�\m
t<
gl��F�2����J�3�pYN������ԕϸh$pĝP��A���@�/��YB�w���1��D-�v�*�b�=pb@�8Z��bҢ�>*}���l�MIn��@�P0 )����C�A&�C����-�����?�.X>� ��]s�m�6Ir~�[�S��rF������}��~�Qx�d��A��������B2�k���0_�ةQ�B�,	�����6��z1�A��$�.��L����I-Y~���8
́�,`1K8.�0c�̥��57@�021�yU�Z
_jA�=5����%]i݃�A��+�r�;?�S�:����4K��
K�=�i�L���=�5ak�l�+R�Օ�;�TE�(i�_����5���yN�Ɖ���Ap�n8J)P�aE}^4�]g����j����hZc��Ę������<��Œ2�W��D;.5S��y�N\ݞ�vr0 � ��7:�`���ccF�����C��d��s����^�'}��;~�oT�q�o#?W���h�EO�N�J��
}����(�a_EG*8ӦM����w��0�vȼ�z<��~"�2k
��q�� ���(���gC���:j4ǡ	�/1��������Z&S"18턿��(�}�����q�Wy�������J �ଋ��N8p��%ؾ�G��n-4b��F#!�*����*7b��Sq���W�p�׼�(>����|�s�c�)�_�����O��CA�X��z��#�rf�M�R�nw�^-�l"v�N
%����7m!xa�y.NA����黹��C ~2���o0SG����(wd���S	�]dK�����E5�r�2aU=4��0�MRź)}��l	�M��]<Ѵ�C�R�xN�#L6"�MAH��T������[�^�0��X4�d�������)PK�̴қ5��m����-+p4]�g:.��[=�ʆ5Wм,v�Փ��#@y�dh�g�0%؅3���Оά��y	�뵈�[*�9I��:_�l�̦���֧,o�=m`蔮�=�ս3.��5�H�겟hBu��5�u�8X��|���IC�)�EU�'��|�Us�1��P��5/S�!�,~s��K��B=�!Kg���j�Z�aOM3�Ύ����'���y�S�I��k��"��&���Ѱ�Ŗ�����|�?#���Ƨ���S�ֱ�0��yÖs��e��n���mw��ۦ�7�fp�:]|�|�vTY�o�Y ��z�_ݑ�9�G��^�	uO�j�
`\:=�X���\n���.����wy#��YZz�,�b���)O���|�ۚp>�҂&vp���" n|ߡƿ�$� d�׮�'�#䃧%ʴ]����Q�L�Υ?��׮�lh��b�h!�C����ۅ�a�x��[�� ���b|vWM�Ğ��:�8QhH���y0�ѐ��t;��$���۬�b���������h�mv�܄�S�nmD���
'�|�^:qQ�������^g�$��Ie:�p%'��+�d�THe�F��i��hpR�;����"e����Q���l��+2-Ă�rGp�s�^i�ۤ26/]N�d�n!i�mkH�B�}��k�#&�5Q ��%�:ғ�12m�.~��N	\9G��Mǆ�mB΢�['��g���P�E1��	�'
��_[@�H���䯟FJ���B�ˋ��s>5H��)[Es���H���{F�8(Ȋh�(�8��c�RH{Y���� �ek.UE�QR�\��<��?${�y0FE|���w����q�؆X���!w�|�b�=u;��e� jp����ZP�qSOË�y�C�x���V���b�t���pٍ�Fڌݝ����6�(4*�Sof��oG6d���P$︰o��ܾ�EoH.	�jG�p�^�ݗ�d�Cz��ДĮ�2�%�,��g�]z��1.�p}�Ա��Ϳ��U��d-�$����>�P$��P�V!�X��×O��Ga��2^��Sk�I�"G�� ����|��SIS^R����6W��f��_��YC���1�@OK�Jm�_�lH��&[O���%�J�>+���V��8ӳIY`y���R�66�� ��ǘ����zY�<����<�Uj��W	�`.����8� 
�)�F�!W�y��f3������Ί��%.'f�������(�D=`�]��l��Tu���O�Л��.����r�۔ �n>R^I�A�o�D_��ᆔD���S\��x70�*�
��W��ȕGY*�d��[e�f�s����K	g�e�U�X�4TƊb�n�5� д��$�����K�D���Nj�_j(�ӘB�TϾ��<�WﶄE.Bmz0����"�_�9<�~CH�}Hmvk�8��A�(�z2�Nuy��Ne3YwBD���p`kTrRO������U9�wE������Q�aAf+ϊ���#�6����|�����u�X�OC:��'����>���f�o�.-��)����׍ ���A͑��6<c:ƢuZ�1�ˍy-��z�r��q!T��^�2�I�iKg���j�@����\V���Es�O=�7hFn�j.�$О��v�Nf���n�Z��a]�PU����H�"��$-�⅒��퇴��ĺu�,�|��V5d�Y��I���q(U���?�B�E����ٚ����b4n	,�_���9�3Ƽ�y�zz3{3T�z��o�oe3���r�Qδ�����?&�����E�u4�.�I��b�%5#t=ڑ�ED����$�������c��P7qij)t��m��(R�D�AQ�h�N�]@v��zQ��.)��D��6�mG��[&��3ם"uX.�ZA(O����M�_�p�m���[{Ld���̜hfФ�S��������w��)h�-�����,Ê���x���Fq/��l�c��#��@�gc_Z�"�[\u���4�����l����K�8�+1?�/��.M�1F\���˖F0�}o�����;��g`58���9_+�"I���]�L%�db�?�i-ޕn�m$R�f�HV`�ߘ��2�y�,g��l1�Er����k^����OG$���.��(����<��hv�]�*B�K��1b��a�
�t����z73��"�Q��eӡ���T��l�:�Ў�a����6wz7�t�/��s@�޷Þ��%_�+�6�y��\sy�ɗ�}�0H?�Dm�l��'S��Ϣ�֭y�e���o�9�$7xe;�<�MJ|��M�Z��
6E6]⋍���ɮ��� �;y]�-ZV9!!3h.t��\'�3M��J��e����K�����_0��[�=�<h�çFK�a`�H�E���5_���H叺����Q��2��-�pL̤Ë-%�����ܹ/@��{�x�x#7-�R���O�Ao�{�7�H�5Z.�x��CR�����a$*�?pf*�vۏ��@vKJge?:���k�tvRt�QA���s��n�H?�;<�"Ld?�t}��E��8��ۻ>�wB����<|����=��j��.8�i��
p��bV���!���n,`fhM�'��p���bs�����.c�<��`C�Ӽ������ocP��lI�*��&@2�ѝ���.[����Db뵲�Q��9�cq��埡���s[�p�ð�� ./��g,Jl�8��~��n	][U�G��E���А�}���h�����וU�Nc�C�����e� Vp���$��61Nw�O���O'�x�o� ���V�ɗ�z������_k��P����������E�c�=�s
-ċ׼&(F�o�@���d���wl�����)�Lz�\��c��kOA%O�gソ�����Ӊ�3��~"���Wt�P�"��5��,΀(�\jW,�M�Y��R��2��O䤦H��y��φ���x{��m�7���_�u�?/O8=2&�ۛ���ߚ�
9-����e{�����i`*�6��H^Tv��5�(#�[��U �6"F��u�F�4�Ⱦ����$�
��:D�.�q�!ǽ$�&l�[񞸧�ӓ"�0,�"��k���� ���;�/r���u�˔����{��zTzi)����~ED\k�佐{y�:���c�.������M����89���h-5��edZЏ�2�ߦ*���^�O�,�а�p8r܋T�L��5A�N�3_��S�� �W���|�}���J�	��K����>ߙ�P��$+Y	�״M��!ښ����'�9��t	��k��PM�99�Y��Bw	�	b4����������G�$/�b��K���7�k� L=��0>��+ kc��s��Y
�k�n.cd�+�ԧ����%�$lU`q���e��P������\ί,�(�����`JF��R�h5��C�e�uȪ'sN4"@J���5�eJ|�u��-O��|�L��Y��=W�N��ʳCC�ݎ@�G����*��T���h�cKuۃL-��	�A�La��8$�f-�;���.z�coH'/��5E����j�f�./5��2��;`�'�U�?�ۭ.k|ވ�r9�-���������^G��E|�j�\
�<��Z�E��'�P�>�5��+��f�p�v�����^;���h�oʷ�Z ;z��z]��5��e��\�J�*g��稏�hzU��/�4`��˘l�H
����f� �f��%��K�h�%d�hW�#J�4��m�'q0���}�o��oS��L|q�d��VK�o�TjE����c�W��N�/��ǐ ĕ��jos��/]�����nR�fȲ�A%9a"D������oԃ�^hD ��ӭ2�{6�9j	���V��i��!����K�R�ʉ?�ݨ�4���������Ȣ�(&����,G3N�=�j�|�
���5|�x�%�˄����PO�_��`OV�h�=7�����_�>���R�I2��:�����9� �畓��}�SPH��w&�.�4wɚk��fVE�h}���a+�X��^��7�Al��t����Ra��Q?����
s�ͅ�� Wg0�8�E��b�Yt{lT��n�}ʱO-�}���m�
��#��������O2lŌ��u#� P3���5��ǒ~B\<�_aǧ�x'�L�儷�+t������ן�M��r�c��N����y!�q1�x�>��ꤰ>�R
V�{�@ɓ構�)R�Xʠ�)�hy3�4�C����2�{�\�u��QY��G�vHZ�c�ߍa����,L����g��*����>0x�v>�;�B˘#~G�ML�Ǧ�J��B~I�>���<��t��Sz�jh��u[�������#�:�"�%���Z�e/X�2"�)�T!Fg#��C�Q���sns��Y��;�L�����v�c�ת��
R���&��������/�D+�c��ѹ�柎W;���0޻Xa��<�@�qҿ�9�龇%ܾ*��P޽9�Z�_����qϋ��̠G���'%'�%?;�۳:�y�rQK�0�[��
I���%�Tl;7��x
����{��H��a�"�i����٦���9�~G����JE����>�6/��W?��qX;��6/l4rx�
��wA3vf���xh�:��ӥ�ҽ�N1X�v�f�9.z�I2ű��>ީ���I��z�߿۳ E,���9���"jE���ȵ
ym\3�)4���S�g���!Ëp��թ5�kLG�IO/`�6�抐�/uI)�)R�Gk�k���ƿ���qAx�ھ������|ݐW0�>{! �J�/7ZY��y'�Dm�Y!���CH!)����A��_���M��͒&�B���{�X1Zy���id���;^/`��{/���[�U�x���Ї%<�2� �xq?W�����ݜ]	�ˌ*��;��ϻw8�&�9��4F���;�gC�x�*f`�g'!	��?Ђ #�y9׉���!荂��t��(%����l�8��k/������/TQk�R�77���R�V[}3v�S<�?��9^s/ �R�3{U��[[Q��z���"���?��m3;[�+1ݼ�T��BW,X�[�@i����/���*|�������Z/����^+�KY���=�z��"��Isr8��D��%�b�c\�`T��=�6im�uG��q8�y�C��7[6Q��v��$-g�8��)۲�Z�l��*5�G���I��V��r5��-w��-S@"�y%F|�g4Q|Ǉ��`��Yu�d@n��J$R�1�X�4��
�kQ�hI��H�������)��o�2���[�Z����Jl�&���l!:e�n���&�3�����Q7,ح��_N��H�xTN�R�}&��Vs=Qx��Cr	6��d4Z�|�$�9��Q$A�y�MJz�ȶ5����{��x�
K::��:���2@��$�W�>>aC��H� ̾�TOFy��?���F�a�g3�jv�*qf�l��t7�ӄ�jR�z��N�X�7|��X��	���U�#���+�1Uѫ-D���ā3��N,Sv�ݑ�R��s�L儡�fa�oܙ�w�ě؇�fZ�0$k#�K��eJb�I��S������5�.��<��#���C
�������`_��d�����:4J��0*���ؖm	3��������Վ�*�^��J9��~���8��[����b���.(���X�O�G߼9<{��[�3B��=�% @oӫCE�3�y�����O�Y>9���Uїrwj�aQS���\�����a&�tm�j�b��duQ! ��A8x���9��x ��q�~�S�������CG��?�\
K��Ѩ�gt����^���3Bmv��I�`���Z<�[�8P�i����rE�U�]���&
���R'cd;�4���_���f]��:+ؤ9��X�9��I�^o����"�8j���Q1�OW��������/|>��V�������:r)�]�x�.��_�ɥ�z�9���lҭ�"�]��y�S��}u��j�i]vM%��:K.�ae�ɐ���8~�n�o�1N��/�@q	�VBv�>f�<�
t�/i%����R�<�A��A���>���d�0�@vuj5�X�X����ߩ]�ұD]�yw>��Q�G&*ڰ�żvU�K~�NF�'�5� �]�&|��O��::�)t�k�6;.�e�qU��M��~G�K�|��dy f1�)m&T�v|>	5!��7����A��"hO�u)c�����=���$Q~��?��s�,�\�20�\z_h��
4���-�[Δ�t��~נ������xP.fթ�k�~��8��|2�W��	�>7�B/n�<w�to'{y<��R�6�+�,<ٟ�����}��#Ӟvz�!�o,(r��	���T��!�߿�%+��������vz����'ѻ���T����
��*�+�1HN(�:Ո��?��8Jg�gX�Gб(�F�X~��z�:\���S� ��=g�j��Xq�Mс�=5.�	�����4��jA�E�J��H@7�gICC-�7\��O芳>}���N�+f �«\��s-S\�0R�/?)�~:,�G2�R�z���>&�;�i���>��󫉚�vk:ǩG�'���>n<� ���TKi
V�_�a��K�/˞n<��z٬�_�|�9�����N�t�V��`�0��.�v9�J�z\:܎�Z��i(x��×�U8��}�&���޳)?�砶���;���
=k�?��^E�W���:+�"p ���g��")���۴�ߏ9ܙ;_�7��y����6}7�W�v���k���d9���	�D��8����)%0�x4����ҩp���L�>N��a6l` Q��6�/�l=�Ձ6��oe�~-�t�=!J`X����>����0a85�;���,,��~�CN)��^mn��^P�����0����pɧf���U��P�v3Dg\%�n�ۖb&�T���r|j���7:�M�3&� 9�Q����f ��˓v��^YG9^�d��O&m�4�U�+h6.��w�\�`���L�'�����yb����Ԟ�*��,U���̡:0�L��T��H�;�B��d���K !%��h
�.w���h�T��Cnd����1�}F�Vj5m���t��ѹ����i�kW^������M���?����ɽ3}��4���G9ێ +vD*��QQ�= �b����*���txY�H76�E\�EM6��m�ݏ|D#Gz$h����v����U�;T�Q��̸�L�����9^��>�$�1bɥy�t(��IYcmv���U��+'�,���ȃZ�:\ba���p�Ikb�{XYc�Ӵ9ޯ��-�^���nJy����l(��@|�X����b�����R��K�f�D��L�N}��"RA�� �� 7T��J�X��O�u�jmK��q�olU�(���}����D�C:�^b���1Y�FT�zZ����me�N���sG�����5
f�@y��ۖ��̸�E��r\k�vFz��1��#Y����I
�᯼b�� !� ���H?29mqsv����v3p�T���kr/�ק�'�kت���:/��a>S��<-n��F�����(�N2�)��n��n��2q��Z� t�K#���AL2�Ru�7'����I_��~I+b	���������5�+D �\z\�E�|pc]w5�a�Q^z���i1	��\i�.��ۇ�ݙ�+��;��JIYk� SR�B�i�*yɷ���Υ-����a-J�yd�Х��U���9�ڙ����u����/6<Yf�֥XR��x� ^��ү��0�6�Lﲶ�6c.���{*W��amhU5)6/���OoIRte�����xʱd�r}DgDa��.�̩�Kr��1��CF�@Z�|��jZ�]���R�N�᠎U���e��q����DB�;��yJc^T]&rdI�ػ݁�S�C,eS�5|�WJ[���њ��0-�Ԋ�[�!t����H��	�z�#�O5�P1ɿ�b��@u3�
�"�я�! �Th
<u��^�*ӞA	O�?���˔�($��Uv�A��1��'^#�9�ٝ��]�b������l�9�N|������O��	=��{���,�D��1�7n'�T�c�8w�Q,�ݻ�2�_o��ѭP,����E�V��S6"Qu�!��(��!0��b�������[�)�'!dShX��B�
S�������L�%��&�������a~�rx6.n�C����*W�\XX XsH��}}P�+!�	��,���.�^ٌ�	aU�=*Ǒ����֐���X��l$���}S��������湔����mK	�S6b��o���S�HLZ�����cĞ�r.�+S���֋���뵪$��O�z՜���y@3V�hʭyAm�{�˯v��`�pչ^k�D�i~P;��u�i�0�۽+�n�����Gq߷��C�׊)0�3U�?�gj��T�kR���V��t
,!�#\f[�L�ƣ�¸�̙A{����p�r��٭���L��4	��"��e*��������y�'ǭL���1�Q��\!��-����"qp$��-���a���:�pqw�
C�p;@?�NJ��]0�-I�M0q䴩�ьe�;������O��n:��Y�d��K�$��1��"�:L�I��+��ٱl�N)��:��ئ�a�a�>un�Ԙ��yް����Z ����9���Xo_����i�	Y�Y&��ka�	&�`�^/Я���E|v��<���l�a��F��<�R%@ +'xm���jM����g^����y�����R[&M�t���&j[�o��w����3�>+]OQ&�b�T��T��!R33[���ө�,M(J�b12�8��Тy3irO����ۼ�|�|˫-�w �3�����!G�"-0U�ae��f$��S��6��B��m������m86ٿ��@.���MRi��|BL*y�Ȼȑ�����ҝ^�<�:��:�ps4�ۋ��en첎� �Q�����X�A�S�=U�z�3r�F��pN����JPW��a
T��Cq���yۤ�C�p��+��m���igl�Y��H�*HQ1��|:t�b`�#����'��`�?�@Ɠ���������DԻ��*���X�]�A/C�	ٶ��jQ YQ|�HX��{�m�{�R��,dq�m�K�Bj����4^�e�!s�R��������\�w�(�|��@���H�9�����s����O�0�d�d�,/��IN@xt�����o�#�qV�i���=�iC���7�*�י����%	���K��B ܴ�hX0],��Ga��V<
������m��W�
���/��[3��G&e��upb�$�ƥ19�X=X������e|����xݺ�-5�#PK�5)�Y�	5���]-l�j�p����}z="u�[M��[��4M^�!L	�&e��h�&wK,؏~	I&�06���Р�P�(-a楂eP@�?���n�` ��])���i���ǰ�;Ьl�+���k�k`D~
H<�.�p�$�\�m��~s<�D��Nf�;G(?�Nry��E�o��-�����A����T$��x�>{ԕR�Z�!\9c�|�Şu�w�/�t ��W(��9����M��$-�V#�>�3?�ci7��#�C�|ܵ��DM;P�!4�&��\RP�m(r�J&�Jm��慀�{��+e �O��B(x�M�q5��D�E-Q0���,�1H	�hi�$P�O�-���_���K����q&�Ne+)m�$N���M=:�whɛ���5���3�
v��p�vZ4N$8��A�R�W^ر��K���a�Af6`���fKR��$�2�
��k�����d���a�݀�7��-�ހ  k#�~��lT�	�������$����
�8�<?���U�+VY_�Ƙ��RE���0n�DA���m�!���N\�޸KR�p%������	�Y*)����6z#��8���=Sk����/5�%N?�x~+.t'`�=�~��$�״����2�$���M<�yC�b`kU���GwﻥT�	+���Xt��g��;��V�Ѹ\�ė�<r�a��a�+��ҏ��Lj��L���;���$`���y#�"p4��|7����U�,K'�j�_a� I�����a�u�'&^6)c���W��id;���t4��p�f����"`Ф����Q`JB��d�?��:Ȗ	A(�To��7v|�郠����eq�ts�ۛ�{�kh�I;!vu�/</v���F�m���e�Q+��.=w�d9�lF���3�G�Yn�\Dʂâ�AS�sT�x}1�8.�����b9���B��j��\/e����!��;2�3�N��@<��+_���#:���=l0[Y� R}��>��/��LGg���
΀�6��꒨���]+	��"���#��#�X��2/]�S6;c�$j��#�֑&�mƼ�&�f��CoZv�O]mu�_T
�����ڭ<p�/��8q���=�����(�����U�=�C����8�tu/w~��`>�����-��A)nZb�?��]�.��K��#�a�Apo��Q!���W��'���p�u�2� ���ա��r �����������I}� �/II�a����/d��72��`��$e�#����{��/�
�}E�����e/b�i=v�����a��N#��!�H%Ho�������k�3[NGi�@7���Rr�ݶ�d��Jɾ�~K�V�-��n���Ѡ����ʻ����k�(�?�ẳ:&��z��#�m&�_��la�Έmpt+���͠me�{<��^�Ʃ��34��.�h�u�WG�i#s�/��:Z�׾�Z�	�)]U!K�y��L]���Ӿ���T�� ���-;�'Ξ6.P�8�t%&Z��Q�����|c��ĆW�:j9x>I0%�97��Sw�$'l��%�um�HUWŁ��$�,wYr��'n�<3Y�ۦ[T���_+X�i�`Af����1t�]�xIfпnT�.�º~^Rg]�z��뵎WA���k#{h�;h}g����7����on��'l+#�H����LB�e<h��_�ߌ����Dފ.M�Z��TNy�Y��V3:'jR��Xyd���,#a���P�ߘ�1��\��_���8�1�q7�A�*���MYe�� ٥C���w�BmŃτ],x�T�W��BA>�ެ�w�[q���'�:sS�L��:��iNh���	�g��Q5�������s4�ߥW���-k�O�sq~�B�nSs8��f�`�5uk���P����"���ֳ��\�����A(���V۠#@<�	х�$��1��+���V��]�$�.�-����������ƣ֐��<�w�Ge��rX���4��,Ld�U��������
��?�kB�f]�MS7� �C=��	��:8�����!�z��s7�l�"���xJ�0�_$���X����'��h�N���)&V_5�D2����;T�ڼ��{y� )�2�^ִ� >�6�"��*�^+��F*ׯ3F�;�Za�Q"\l��q9�!�f�
�F�{�4��#��@��j�=Z�t�֨��!sD�A���a��Xo���͝xfN���Rp����3�
^��i��\R겷��ZB�-:{���{ί,�+� T�Hn/�ᧇ&�������:��,��jf�=�{�쒰�"S��[H���Kwe����x��ػ�؁+BW�����0t��O��U�Tw����=�<��?;�K�*�2kΫ38�tX�!Cަ�|��[��*�J�,HD؃�k;c^7���,�ln#	�wBg�.ވ=�,.�=��6lQ��Z�K�<���9K1,БG_`��ۅ�Jr�x&
{z��:���vT�xӘ��b�i��P�!�����rUP��`4y �ܡ����JSw�P�A��=�BssJLC�f�Yy�S��YVB���O�
���4{O���v�9yl��fp��	���Y$	�+ ��H�3ud�tt3��z͵-G/ۘi�L 9v��[����UQv�{�ۚ}��n����VPz�$�}���Mh�Ԣ�
�e҃z��{�@e���v?���ŊH��I� �/2I���+�s���L<j=�����\�Z ,$VT+��A��H��v+!������F}m9��u�HBQ�Gyě_;lM�P�^���W�O;��Q��a���LT��`׃�����W��`�Cb�[kY�9��
�]�~�h�[�1��ϣeF�_S�$��W��5��#��I�a��YԨ�$�~��SZI��!<��0[�yq��Q���f��DǬ�69��Ue����M�TD��U���8{�gR�73^�ˆЌLjD�\}]Q,Hg�J;¼OUyB�i�w䖹�D�오+8�r"�:�Ӄ�����)�_!�`�65A���p�lҰ˛_�Mxg8�3K�)`�>�����c�ZV_�sŚ"�Q(~V�n���#�A��ҁ-k3��ř=���͘�k;pA�͚ϐ���DC���wZ,�2���m��Y�.�K��X��Y��rM�j�}�T��G ��8jMqX�?�1K�_�z��~�+��B��^@��Z���B�u�6U�ۚ�Ak��uNPoMw����e�?P:9��ey�a�(�?j�m}hvg��:��
�l7�����25���]h��Ga>霻C�0xf����zd����v�ϫ��=ܞV����y�W��ⱪ5}�����ʆPM�Z�����O��q��_�\������?$�	'���B.�7 �2%3b����WRs��l*�p��b��b��4(?ts&='�}�L[���q��䵟�Dmf��g�}1(�����X���_H�X�ݔ�M��m3ߖE��b	O�ɛ��-����<7C�w܋���!k�5�eH�?A@s��l�5��y�Pbp+����܆a�d������@�⾟�=/ �,�1�b�N�d�����$�QN���a���t�r�~���`e�8e-\[���0+<*�6mM(��b_
\}������Z0���YJ|o�M����z�L�6�G^�"�����Թ\���=3F~p�<iu⛩V���d<��7��Y����9��ilf�+(��R�L���r��^釼�#Xq��$�Y6y(�]%X��� �������������}z�
��3������p(�R�8*��y)���Q���E�~ �z¿	��V��I�:[�T#	��:���t���T	��4��&��n��H���}��	0AK[����	���dA1���k�>�����0�M5{��|���Xkm-*y�юC$*��!`)�!���4�Z�fP�����G%��������i�����Ƨ�\�����~c&��;{�#��&����zWh;���Wґ�]C���Ͳ�^N_�7?g~���l��55��@�Τdܪ@�|��t�@��:5���Jn��~������B0r��*/�%B�H��+����%��e��>�w�&�2Hv˪����G��*�m�=�#gΈ�@!/�(e��SRT��r�:Om�������UMG=Td�"?�s��]�e�=�	��i�T.��
����L�>fBfT����[9R����笡��tM���!�g�����J�D�A�0�\��L���5K�Va!�Y! �I'��M�8���k=�n �]�p���ʬ�2m�O"���r��6b���e��ezE��k5�e�D��m:�kO4�Ҷ"�փ����d�Y��HHFҍ��H�!����%�b�waQ*��]�L��x�,�)��J���@\	6�k��<M�S��.X��������/#�iO.+q�� p�btD��A�!���_�P����P�-7�l}-�28�j�X��6#Pai,���,�co��"@Z�n'��B��|"��Coo]r�$��n�^Ͷ�@�t�w�G��B�(8޽��7�>���7�h���"�p�w��]��F	)$@�\?bO���.���j�KM���N����� ���!�����|����S�$̂��ެ�r �ɲd.!�v��9�R�eAĺv�\���'�'7=G)��q*��6.��/�m�sM�'˞�D)�.��=���25F�9�5�'��
���M����k���K[.�� �t�����e�m�#2f���juNL	�S����u�h��)�x�**0�l�򀍪�|��"�Pp�0Hqo8*^+E���Jf�Q9~�Ɂu����r�����ZE�ߤ�'�;>�=8Z�f#���7�Se�(>��ZB��&�Ond��������kLeU�� ��L����#P�7�!���`�1ߦ��Y�I�:����@Y	��J]659R����q¤�0�1H~~�m/v+�+p�Oq�o�	9���{�4��6Ȩ�D/_�DX��.��|���bގ)X���H�X��7d��M�ME�S��nuy��y\s\	kh�;��ڑK�ؿy-a\m�ؕ�rD8�P���s["�yg܌�4[J��
g���V��������'��О�������X���[�P�?9����P����@����kY��v�v[�bq�I�m�X�gŷ�h���۾|��CI��I]1�`;�"[�5�zdVr��g�Æ�i�i/��2K6�#��a�aohZʠ�$�p �8(l���-�ͦ<xQ�}���qy�PL�:;~Ưb��:2�I���a��R���S��$�V:ĥ`(Ԑ����]nń<��(�֏i8�w���R����޲��4��ov�y����[���)�0=��|�4�モ;�L�Ȥ�!�6w�I�o'@�3����6k�����όW�Y��=�cq�׎PM��q����@ �Ϟ�0�+��C|����	DDPbXG2oXW�����6�bX30
�M#,P��Kc�����u�z8��,:���$*�`!E8`�j,���˖�Ǚ��l�9�K?W�1�7[��6$?����n�I�y̱��Fٷ�>���QJ�K��X���P/{)���`j�xN�ˍn�5_�#��U��y���Dbu�S��y�В��(�s]ߍ�P(��PBAk�Jc5K����^�%��
$4�㪿��B�;�TT.�g�t����U�J�7ݔҬ�=|ȳsՄ1X1����f�Yх펀RT*��3ţ�bj������˵5��C��f�[�ӂ���M� ��?TmKK�h���y#6�Es\��i-0O��4�jM/������F��5	}��&�&�/�Y�t�d�8Rx者���S�|���V#*3�HY�t�$#��.>}Ŝ�X����8bx��pT@Q� 8�P'�9T�3O�:}�`9�(�&9��H�0	�A�0����V3����8l&�_�r��Yh��"��y�K*�gN!
P���x��7L�S�" $�5��e�׫�ź�w��!:�mX0Ez��f_߇��RS	����=�]ehA�?�0`hBQ<�Z�����!�����-�8!��L��J��ސ�#Dt�w%�]r�_��c���W�ZM~EA���\�����aą�-�=����R:!x�2�~�. ���iz���kЇ�����E��=7[MI{G8��qL(v �+_:ZּFG�<��LW��+�P�1�lr���.&��f<[<�c�m�(���OiS����c�T��>���B`ew��y��%��g�A7n�����JM4���2N��<�	��j��HKc�d0w�Jǽ�� ���	P�dۈSKT�3 ���E��<ID!�E�+SD�2O܏る+6N�p�� �E��H��=�Hs|�$a}�ff���)���{����l���x���/�zC����c��n�3��YR��03چc�����x(Z����4��x����y?A��O2������<�/�v~���Wঘ�;%읯�'�$��B�j:���5ա��rr�&r��Z3ih8T&�b֢�1%��d�w�y���D-�5�� ��T+Hb=�-�c�YL�X���oN<)-���-r=p@�qc���>U��ε0��g�N�ą�y_�NU2��GA��g�&�B�4�C�`o��ltbzH�Jt�e5(�,����])!3Db-�L'A�8E�� C���]T�V���	�B]���,y����D$�xd�/�R��r�1�l�廘���s,/��M��&��w
�<����=3@��6k��z.0�م!݉�.�M�<F"���""��ٳ�'����o��>������� ���Qm�&=������ٵ�!��g�b��� ���B��ي��D@�J>G�䚄�d:W�O��}W�Eq�;��
�UT/��.��{Q��%�T�{�hj�oXa{d�(�xc<ɫ�p1ᴅ�x��94h/T���Ϫ
��|	�_9��/Ч�;ݻ=���pc����Az�������v8?��/T��;� [V[����\��j��2�~��h�A��ޑB��A��L��^xkcE.��XФ�}�>Me�߅�M���P�:�wn�F����s��=��[d�6�q�P&q�Ѷ\���oR�����\-�z�?�V�]�7�*����4^�e��:��so$.B����{��Jp�i�j�7HƲ�a3�T^̜>TJ�aͅ{�����<�Ylu9�!=l�ۃ44�o�Vy[�}[e�!9�aE5¤=U�V�a���6�y�]��^�$��ɳ���yO��o�{���"���$[���7Hn7::�d�`���P:�[3L�E��_
�PH�Ke�)���U/'��$JӨ'�UY�=ľH��t�!���q*�J^��f@�ڗ�/,����}ڬ����o@݇@U��Ul����q��m(؄(� �kJHӜ�TAS����]��/!_�_�I5c�����01�v�W��	ʐ��'��qbh���̓S�h��t����h�,u�-C�iAM �aŝdi9�;)1�2;�M^�9�`C�qy�8�c�Z"&�ô�\�5Ғ��M���i��}8b��kɒe�=�~}�1�{���ZC����H�"�ި��M�s�f�[��������ya/Hw��O���*Y-?F�فG���5p�'��l�^�Ov^p�ߵk''�j��q+ܢ�d�NlNx��z�BqTto�S�o&M��5�)}(��vb����%�77�.��v�D�H5q�L�k�$)T�ֿP��m��s��E� Cox��`�p�w�B�����˕Q$C$��}_��Dw�sj�hIJ��uW��1�|��;��jj���ѽ��)5�I��CȿƳk�=#�#������5��BK'9��%6�u� �*>%��H�L�! ��q�s!u;�PQ��$���ا�b�9��y�1�K7Iě��v�����ksvA���
4�1mE%�GN9T���߀��2�����~g^���jq"�N]0���W�f=�3�L=i��w~{۬�o`�Ut�-L��n~
s�a@!߰X �o�����u��p�A^9�Ƕx�U��
������W��M��;��6�\��A{�6|��!'F�h�5Ӭʫ�Ui1*Hj�������֐���"�ҍW���T���s�<O�R����4����\B���<Y
}�k$��f�� w���#W>�bTy���6�(�t�xn'Co���ui�\Y`����c�������⧥��0襑f��F��'<S��b}�O���ū� <��^Ѡ3g�Nz)��bAL����#�Vj+�Ϗ)��)���~�� ��q�+����`���`���Fc�Qk,�q�S��#���6�Ud��	����� �5Ywu�b��ç ,���׭��7|�VzVD����.x����#nJл�S��ke0zT���W0c��7��Ժuu)�:�e흊��
�<��A��wQ`���> q��"X�6ɱ�6�r���I��'��9�\2l�n8a���q�"��Ź�z#4P;�^iI�6�ϴ-
0d��P�AY���\&$�Cڼi��p>��#��F�us�:�d]Y��)��I}��I|bQ�&j._4u����S���˹����Z���0����}�α�wա��������2�;/ uj�3W�j�����L�#_�9Gн�E��H}P�pU��4pyx[l=�7���mD�Ũg>D�X���gC�;w��%�A�X����wƾ9~�Z��
���&X(�©�~�0�5��ݏ,� �/7m��WN��?=��sxz���>Є�z�	j�v�9+9n)��81<!)�|��Ct�W��ͦ3L��4��r��e���bl�$�פ�����W�����Jն{u<��k�^t��lzᔆo�0�a\���`#
���i"��vR�a$�V�+6B2�B��d��F��Ɛ�p�Ӗ�Z���K$�q�i�!�e�/�	2H�Z�⨥|p.���N���S4
?:���˚%����&C�&,Fk\|�T���ط yS� �N�_,I5�Qv#b��@�u�f�C�B�xp�1,k>J�G^�c�m�))e]�����%{7�����.����#�i���"i<�Fݍ�:����(��oI�b"��D�S�o��L���*sv��X����e�;�}�Fw�9S����� p���\�d:�%�@H��~�������?���卥��7�I.gyUʈ�Z@��
b�W�M���<Ժ�n���8ڰ2�L�j
���}���l�6�>U�:��*�����[!�����Ȍ�j.Lj6�/����mW "�֏�bƢ�N�[��ٟ�Z�۩s��=_��Sq�𬓪���	W�f���[�l �vQu�A	،�+�3~��X-��n��.T`�ԋ�p��N�2(�a}�g�N�c�6M���5���1-�C�.��F�+�E�2�������T�x!v���$��&r�Km|��1��5��Ju���4�X�����G��#���@my]��[�"�4�$ֵV؏����XJ�w�����]D�4~��C��S⾊�N3Ś�x�t�hD��{I�0/�`moy�X�%N�#_ص-�'����4��X�]�%T�%Pʢܸzl�Բ�AڔUG9�΋�/B�������~�b����9g�s�}16��b䩽�_�1��*%�ݘ��Ԥʣ��y��x�1�z3���|�/,��N�gws�)��#�6AK'3E�t�Y�K�����̦���h.��)yۿ�����I���W�UH1�8?x��E����� ��Il��\Dg���*�A~U/�:(��7�G�#�����u�dr�[�cz��x3��NmF.|fO�	ynO%VJFcC?\o����n�T�x1X�Т���bI��Kz�"dLF�P�_�O|)0[`�����[��5��#���? �$��U_�tl�����3祤0LiP+�)��v�]Zڋ��D$�������jOIW�I�@���ӴŎ>��"���d�+,�V��ɱZ0й�9
��1ku>��c�z�EA\+�RX�d �SJ�TP��&Ŕ�6�K�R�j�tNx
��@��Q�rI�K3�f��Wl"�����g|W>쌰�L\��R�7�jmjŒ-	��A���p5C�Ѓ�gjY�5��5��:(|�gQ��s�ۇ��Q��3N ����ݿ����������C�!כ��#5��}�����[�K���� ������_g����/b�.?X�\���eE��!�ݕ�܁a �B��[у��(�6�{��e���Ű�_L�_��[."�s�_���~2ˏ�Թ�6�8�62)�����Dh[@���n�6HN�k
����Cm������N����@�q3m�'S��vn����Q4�s����;i��b}�C��2����'քׅ��xI��e�y�KV�l
���(w���� V��~�u�����L;��?E��n�z�� �������F@�`�~m���d����4��Dx[r�~��3��8�΅�)j�r����oj�h2��r�j^���H_�o��(r�X��#L�� R`����`�U�9��N�F�KOf�j�4�)��fm�(��i��!�	+��'_��>�>���ʍ�^����SX���`hC�.r�tcZ�����Lc�Y�B��{�D#��2��]gC����d6ќ�cab߹��:��17��8a+�%�/�%��
]�*Z��B֕�`����T�ˤ�SZ�_��0QF�����ohG96�w�.k��B���y�$��T�������!�-�����a�(��H�ӗd��^T��W\�.��EL��=q���Ǭ5�ajV�XB1��s��OaJ%��i���k��X�,<rMƬ��<�0�f���$($>��:&"�+6w�#��АMV�EbL��bFL������cJ取:���t.�Q��3�4?�{�n�A����K+ᢘ�F�Y����U�{w��6p<e��u�8�6'N_�u������W2ȵ�+S�v h!H��2ޚ18A_�U�̗<�y�]����z����>���h\QD"o�(o����y[�J���T���jl�O���݇i��7����)/�zQ/�^���}��e%�&���ֿv��q`ՉЩ���CDC^�h���ζ��KQ�ӏx%0��3	�*��j�����5�1]f��1�2��a�wR}�C%/`�܀��/��(Y�������fu��gؔ���f<�8�%���?É�ϕsEh���\�p�Q4�f���8X�H���rJf,�T��P��D��[ڃ������zsl�+R���P�cy�
[�f(�ӻ���Ս|y/������kQ�{x����/(���L(륷m�F��\4� �I�с׍���tG���FY��C��d}�y�0��0r�TLG!k�Z]� ��JA/����	�����_p!� cm�Bc��$�E��J�-�+������� ?$�ߐɝ���&�5/f[��CK�t���/������*7�	#;�X�CG��(�=D9�i�5����9�qb�B�{��㓭���Ψ�u�� *��[�$+��w�[���2�����*n�o��՚6�亓�TE����1���.xVW+���G�5���y��9��H�h̒��`K�d�'�H���S,9�{���:��G�3����ٴ��Ăi�|�cU:���~�E<h��9�]��6����Pc��2e�X����R�u4����>G�W��|���Rƒ����>��cr��	u��L8 ��=Б.Bn�S�X0���B�:t�����?J ���&�TsH��1�=G��R�a{��9�B�E�e^*ue�[���ID-n�����A����Hg)�h�;߈�*����V�郯��yg<����)?T��
+v��y�n?w�����)���=4@�