��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|��I�ɖ�a|*A���SzV%�"��[`���T!c"V���t�^h/΀�y��L� ]�m�jk05"F�a��B�a�l�\��!���U���%�1�Pj����RG*�Ԑ7h������<��G�����$�7��9%����w4����8^��Ж\(�eK�K��B���ln���U�Izr�-���J��e.��5������_"@~	�n���E�����\�|F��[8�wr!Ub"�A���Q��F��B�c�pv{On'E*e�ήpI*�?*wV2V҆��M� f�I�M�'����djԤM8w��e�
l�����J��z�����a{QP�A��BK�u��$��/MγV�.C��L�����K e�9r��~���I��3^~��	�xMuO�uy#���z�����{j������%��E��ʅa� Ԕ�Z�R?���k�/��&{`B�V�N�"T�.�a�d{!Y�Ah���`�����S���N��<uJ#�,ǉ��-��_�-�� GLG7i��f����1VV�����S���Oѕ])�c<懕��0�2�ri*xO�r�J!�\�[>4��L�c���Qb����l���m���4��2;���Ms]�����N�tI�܂1$[#� �&ձ�kT��	!a7��L�7��iz�S�4��ua���ܻ��%��V��m��e�<٠9#��������:)��f,�R���/>X������p�����j�D�v�H�?��/8Xج!�ɏܹ'��Y�Y����$E,��5J� $�����y���ɽ�]���g��g4҄��l�O�|��ä��Ɔ$9�����ѓ���0���&�[��[��K��)�
(��w�<0[Ǐ�\���{l��ojX�W��n8�$�@S�Q��x;�<g~͡ɀ��2�Ht���,����wĚc֫/�cXr2� �w�
n�.Xs�~Vu '_�Ê�ܑ9�����O��Q6B;b낄N�Hmz�Ea���i�
~Ж�� L�xΰ�I�.� ]K 彛�"U�u�]9���^#ݲ
�8���n�f�PL�͎6P��VK}g%��=�#z^��Ҥg���\^?�7N�R���FJT�����]���p�)v�_����>��qb����~�D]�di�μUF�����^�}Bg�c���ܲl^�ZA.V4��(����r8]�!{�@�~�Y��v����Nd�՗�o
e|��V #��ƣj�<���װ_�^ͅ�Z�KZ�Pd�*��&���}��Z䞤��Y'��E�%n�����N7h��[��u���59���t�7��Z׻�Y���E]\��3x˯;X�t���V�^�N&直��c\�2�m}�9�#��i)�t�[�]�jy��h;�vׯ�M�L=�-gE�]��@t��0�I�÷4�^�c0$�-_-j��$��n=��@��ϝn:��;T�8?ZA�t�S�^��]��]-��<�Ǿ��ZPK+#�q������P~��-~F�B_�x ͓FB�~Q@�]���i���i��$ux��'�;�K�;��(����'��ۓ��ܵ�j5I��篏��8y�����T� LHZlt��}���D�V�O���r�a'�ͼ��^���r�g>`y'��L_|4�֮�m�2�$Q�?[Y"xU�9�~L����PTH��/F#���+Q���m��܉�2�,:�dȈ6�.Z bҞ��������e�L�J�����I�p�tx�9��x�VPhjw}*�*m�T
x|l��P��� �X)�[� I���`-G�j��;��v0J?s��cؔ���4l�XQ��gmG|����K:(�X������ �֥��w A��W�0�-eiF�B��E'!�bΈ��� ����z~!O�>)��+e�k[v�&� �4a`�O#ŞM�&�zY�R)��h���hzx#`���H�&���=2�3���@U�>���7s�ry���F)�DS
��l<v@v��~�u*�����
��T�9{�a=�KɄ�)�/�3����dg�_��B^���D�|�#�L�+�!�I��~�����#�B�6���f����NkU��������\]�0�Vi>+�i�h?�����f�z$�pSd���"H�����$���b��%�y����������v��u�<�2ك�Ƒ����V��H�c^�;��WL�a�!��)�
*���'�s����IA<�l�7[��f�ܜ'�wK���H���Wg�[��FFt��cc������(�S]��n�D�<0��=m}.^!+8�����ҋ��I�=���j	SÙ.���:�V��N�%�yY���U�T�+��4rƎ��.���y���0�������c�=>R�R�5��|!�Iد�5��dɼ��O����;_`�8�G�����:c[�{L,��}�nd'MC�]���S��0�5Cف͞�����	�3���m�܈�9��ZH!ð2�ң�1�vv��<��:�W�}&�
��=�I��E��K4�q<%��]�¨6;R� �#m��Mu��_�[5�p)��W��V�	J ��_5�)W��S�X��U�!�8fx<
l��}��ZEW7o��tq�솇�$+T=P�"b�h�1�� ].d�a(�p9�`=�f��t�����`A���2�{T|�r�@4x7ǿ�������6Ԡ��T���U�����|�l_R}�$ �(��J2�9j���9������GŶ�q!5�r�'F��/�{��:Z����bʳ"�`y��P��* ����0v#��*Y\n���+�(�N��xS�$��.��6��k(����gy�<:1�3yW<1usA�W��5�*��;�ҫ�ݚ*���-݋�#F��mz����ܧ�J�!_�T��᪄�Т��a�߇�(oH��)Hf4��v��_�3�y�AUhi9��X���Q6����t4��6�"a7/$�F�FpYg�v�+=�����?��.A����od��`�Tئ�!B����u�F�%v�e���������^TL�
��N�����H40����nyĬ�9$�e�������9�'��"�/+fa{k�\Nn��������J{^��R������D���-�S��"�g����>Ra6i�C��r6eA�9R(/�½�X�\���w�c��BYH'AE��"��H���7��1r}��G����\Ȧ��H=��A��� ��Xp�q��W�'dJ9�O��M�V�0�Q����t��ĭ
����+|kf� Q���DN����U��M�)W��h%&���$l>��EC���N_���9aŝ���W�\�5�/��+u������" n����OL��(s���Qk�	���(^�7*��oS�<�]���{l���7��!���|�
F4j �t٨������Tu3�]��L��_n��BWS�9�,�Б�8c،2 ��r�8/���s��%��/���x7��m�M���xB]� �����@R�a9J�ֲ�q��*�aj����ySwE���i��酅H�HK'6n˹�d{���ƹM]��������2�W�+_Lw����G�\�iI����)��z�o�&�$���볖[y��4�nY�� ���KHP�-��ی�n�	0��đt5���-MA��ׇ��H��y�����k�锹l
�TwLW|�R?,�L���ܲ�0���U����Y��&���D$'���z�u|��\=��y����}a2iYT�