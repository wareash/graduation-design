��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�k�۸�m�i(b[�{�㇌�]�i�5'�`;Etg
<������H�W޵α���N-�`��6����ݾ�FF��eF4��_}<�ےA�[,�|{�?r+-��5K�z��!��[��S}Σ{$Gx^����c��Ʊ�U�I����8�v�#��������)�3 ��4�Å�Yğ��p{�O�B�vAl��|@&-,�����@ѪqEN!��Ҏ��o����T��'���D�앦)J���$���wY��k|S@e�2`�ul�]�B��,�1u*�� ��^�
�VH �p�� ���/��I��:���v���V<Kb�i-�EV���P���Į̽C�Ӗ>��K��१QWy-�P��t���D�������j#��q�q��靅��l�� /K�_w)�)�Oq7ѡ�ݿLv��/�+��-mMr���+F���xp+
�.(�RU	�i�!��ɼ}ϕ��F�~�;:ٸ_[�t�c�K�¶y$�5�dҍ��@aM��6G�ƚ�(��c�>���F��td�|��������ALB��iq g�!����SUަ!ώ��wa4P��@�9�`I�0 %��G�E��yA��chdZ��W<[L�fQ�A���n@�.e��D�Z���uL
��4e�����u�W� ��h��ϣQK �����p�84?0����Ɲ�I��A����ig���ApOZݽf�B���!��/�W&%�NW9��V�6�똼��jh��`@y8��+�[�Ku�5���C^X�ܢ�@f֬�S�v���>�&�����m�ͨ�N��j�j�_�h��;�j�ެ*V�"�,�A1��a�+�κ��U7�%���S�0�M����� ��iWr�ۍC��
�4�h���v�·ϓ���@IId�~l��~eP��u��4^�t=TK���E�zp)�M��jk�m�s�+BF*�p�Æ�N�?�{�����s�H�'%d�� 0��c]sV���vE�Qo5����p���e�FA$Bԙ��#q�~��{���sk�N>��蛝sG��I��Q���t�c:�D�[ :!����}a�u�p_d�(?�����ӡ;���dLd�%d��}�Zt�A��✥0 zǢSa��^@�[&n���h�d�������pλ�`|SZ���I�t�
��¯84Ӭ��.v;���ˀq��ۦ�(��_/���PT;D_wu'����,Tn%(mH�'���7p7e\��`�h�#qʜrbB�|�sq��y&t��=[�$`��=���B�^��8�2$��بq�A�4�������ўWH��#qQ�xS���s^�T��8���=����b8_Ѫ�wc{�4�|��E�g-hץT��
y aYZ�nv���c4��S+A�9����y�$��������4mK��O�6$T�'*��������3J�g��]<F�^� ?�p�Ѧ~V}U.��F����Cav~N ���w���'h=)�����p�[��?�N������B7l&�P<�t��b�P�G�h�<g��}yJ��*��8'���@Z}���csT2��\E��YU�T;;x�x�C��7��v