��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jåا{�\�u�?߷�dn@6�zf��r������;,��o+�[��C�����a��a,��$%	/�1�pi1@"��5�~�4�K�7���9b2�1�3(v��r�Fz��Y��\sG,��-��Ǩo�V|%SLV)�д�mv҇^����gM�[-M������;{�e�Q���A{&:��XB�s���p/(��[;&BUM,�ѫq]����F�h=ʟ{L��cxy�D�`�.(,��1}۷ vKB����$�A���R���r�3ī-�*v�|x(Uz�!%�+0��@Z�Cƨ%x���UV�<+��s��x��Ǜf^�%�2ܲM
.Bm�I����bJ+���1�@�iDrr�E� O��LY�C`8��-���@?�;BQp��9����fE���mr����v��#SU�Sݣ�PN�Y�L�3���z�m��������и�K@+Q�q�/q�i��ln���m��cB߄��' ,��t����� �tn����{j���+#�b^U�X������K�=�Sy�cs�V�;�-�N�b���f�|0���~���:J  5!H��o_
N���w�⺀+�z�b)b���2����n�M���q*Ĩ��|�CŮ0�1��\�(��!�����F��[��mHZl�BzN�&y��E��+x7�-0�!����<.=�[�5��e� 6��e��d���(�a����P(��//�~՜�����bc%� ��zt�QE!S�y���hqqF1>�ܒ���3�4>ZϤ0�r󱘩p�NVY�}%$�\�&��`n�%�`v�&7�=\Hўa��Ǹ+�SL���Ǳ����	@mާ	��<"AJd-��xh��0�9o�h���;��c_���i�F�JX�H���ǁ��^τ�g�VU�ݓ�~ �~�N�!m\!����ʪg3��V������Y�	��+���]gU����z��i:���a��&q�����gIX��HK�N�����M�z"�D�$4��@K�;�NfΈR�2_88�;��p�{a-��vR溱���,�Nʡ���������ܶ�&I��	���$s������t�q����B-':Y���	m�,˦	dM%5A���+뀅v�U�H\������ ��?�z�r"�R/��u7L���dA���'p6UΆ�M�q�'���?Q��8_��k[��/�C@�\+���h�J���~��$�����+���fD�UF�d6(��G���v��w�����l��=�F�[?��֎�3uv�i����d���ڵ�ex�8bt}&�*ū(���πp	��۟Dqp�	��]Q�K�{p����(����e�t�`�w������vZr��|	KW��'RF^�!�������j�W���2����b�vY}x��N�r�Q��PXaZ�O�Q孌�h��5�m��y�Ucz�ׁ�w�7%}f��3n(<�A��B\����C`��n�[�*
����2��-��^����0��5+�D��������.5��9��f�N�x?�����d1G ħ�n2�ŋc�(p$A��,;}�x�������l�B/�$e%�e���U��bގ8�ĈE�n���%dG�������#N_$�$9����$�Y@S�M�^b�P��Y�<a߫�Pu�g"��h0_ڳ�J2��0œ��v�	(eگ�BSh(R>����[x��W��3�.:E�V�H���r��-�� �!���|W���1���u��wnC�Ϸ�`��G�p���ĥ��ε��	��#y��"���h��Cá���>͉���rQ���˓5#}q�Zk�����|��+�-�<"tſq��{�*�]]L6�A����@|'k����^�UH&���z��eM������$���+�?ݨ�ʘ}��჊���3��_bI�R�x�ku�.(}���Z�V{�w�Q��xy��L�C�����YK�^��φ�N�%�Ƞ��T�`}�GT0��ۅO��.��xy<}�sx��m��0R�^�\�m�򻘑�cg���j��XS�'V_D����#4�>��NJl3ܬ��+��u�5�H�����F��zKq�d����'{"ha�v�$3S�����hZ���J��)�!��G�����P���@���"6�^Z�^�������B�-��MZh쵅�ȭ|��Z��q!�m�a,�W7�ߦ�<��E@֟i�>����?;[���{���|7ʚ�����@F�y�|u긯�a%��N�9�_wn�����q��3*�=XJ�^����JY�M;��;��8>��]����)A��b9�~`��$V˞0�=�����ɟ��nK�D6�&`C��l�����ѧ~nGr|Uqd�,�8 K��+��<'�����u�8R� )� �@����l���%�
�e���8>䅨�O(�|�P��خi�� �a7�NWO1�oh&�{�f5E�ۆ�C�Z�so���&�Y���Nncwy�*K��k|}��]�~�����I��U~Lyw��ֆ�Eʬ� '��-������G�}&~���n���<�9��x�}۬d�jպU
��`�%\�T��b�pH���R��=�M���~z �d��i���"<-�7;�͖#<�)RO+t�/����ʩqυ��]#lWa\�a�eٗ{�1�:��x@l9h聂�9�y~��������ځ��E��R=��g79x��6�ƄSU2L��h��)�(Ǽ�0ź�l3�Ȇ���Z䃿0a`c��Kex`�R����AA��Y�(���T`7/��/�����/FK�*�V��A�֦pv�Ar.l�59P4�صǣTy���r���4qW#q"|�@��蕦:�/�K�B
�ǥ�0��V�w΅���³n)��rb�"U4��W�S�a�U�Fiy�n.�tT������ m�M��8 l��Z�ތU�'�e��������UG�Y�bg�j@%G"1�V�2� ����t#��
�臏���s$x�`y�4����Zs7$�5�g"mc�ߴJ��$Z�����s�ܥ'q��6�;ͺK�	�uv8\:Yo�88��3�hPF	�`�K�B�rv��Xvw#C^�@i��Ӏ,:�� [�RC�W�A��L"t�i;4G���Y� ,ѩ��j.�3���zRlQU'PJM����s�Ɨ~���RA���a�3^9��@~����JF�!�D����w8�H�v���)�)���ǔ����#����T�H4��0��G�<��+o/�1~S�ıA�Z=��v�����\�>�9J�|Z�C��FХ֎�:��v� {�T�喪O�3[&�sβu"�S1���؈���Z���ܠ��Q܊��r#���#�K�=����� ��j�J�����U$"�&,�P�YL�uF��ݓ[R$-&&��I�ft�_�H�K��B ��՗�������]Q�Z�0�Pڿ��c��7�5S��HX"�B����P�'��쮥��ɑo�X]wt'��*K�^������@CE9���P��Q����p���,(g�p�	�$h�;,����~�i�SaO�b��t��jF?��@=>S��$����"�X�x�Y��>w	��)$��9���l�������@�~ū�C�f���9��=xQ�JR>��+L�a��� �����_���y�5+��ɏ?����pZ\܏��{�,x5����4�����F$����[p�'�u�_`��S�X�ퟍ0�;/T�0�Q���U��#μ� ����o�jY�-m�{�:�}��l�����@-Q��/5#u�b��(��Gta,6=B���}+m4��l�&��1����]���·�,����m�^�3���ϣ����-M	�<,ԩ��͋�����׮���)o�q����5��Flo�.Lu���h1�El}��M �
�z������ ER����Ȣ��x��u�la��y^#�k45:�rJe��]m���̞�eb�.���`e`҉CǦR2vθ�~��YQ���/�L����WP�� +�)˱����!��a5]?�=mu�ER���/Չ�e��PD>}�[}0"I$t��E�/�C��d���F�LW;�3��6�(kQ/�H�e�!�uI��c���nk R�Wj��Fm�]gc#*bwٞƧ��9��bn�޲/֚~v�Q�/���nj]*P*��c�I�n�F�rn�I�:� W�ͥN�+ ��b�:d�k#*5���Fҏ��?<�s=M��Z� 㪅���Yp�Y����{�=�|j<�{�LE���.�gށe�5ҽ������G�{M�\��q�"�ޓ�8�� ���쑪�/!����rq�#�S��i�£�E5�D�$�k�[�7�ûfb��h�孛�]DW�$��|+n�Ϋu�g��#)�e�4���E�aH�����hqI�LF���=��x=�X��hO�?I,���v�D��e�M\M%-���WL^U��>"���5�.$5]�Q6�4�M�*�-ɑ�~���Ƨ�����܈�a�,ڍٙ��7U׺;���uD�b�����ftU'3��$6	|���N^ve����=�G�����?o�I ^8D��K}�to���N�oV��yb�E�<�03㛰%�^(�j��o!� �i�4�<�T���4�}KN�҄��)�.E-��+>�U���#�0(�I^.sn�ա��c��G�f��A�A��)}4�E�jt��f�iFN� �!sd����`�^���&?\��l�?������'h �q�\(�u)�m�o����^��}]7���Ӵgy[�b!�z�����S�Q���>$
{����ckc=���+�u	�CF־��~B�t%�d������?f-��nU�W��
�r�j��>�\�a-��Ժ�S�`��2Cb�z>�9ö�#/�bO�E�a���������u������vw@�qm��q�ՠ����6M/�U8/����q�^�4Z��9]���ө'N��}h~~���R5t���x�����Q�!߹1��#��#�	w�x�[գ�(���
���܋l�B}���OP�g%$�)�G��K�P�
�i2�"�m�X_�����9�rf"5MY2��#/d�P��Jm�>V,M��ɍ�q��`��e���QH��*P��P!*�Dyq��\~�?C�Cu�"�54���%��; m�p�5��_T`U��N���,6\����eC��}&:�*����@���4zЗ��ջ��C�F��"D�=LO.g�5�?�c���T:0����@r�T��XN���K+�У��V.�r݋� ����m�#}��MZ��Sbr6�R��6u*���9v2���qa���[���h�����4�(�t���쾖�O����k+�u���c�7�0ǅj�vbgO�h��O`����!%�Qя	]��B���5��{h��,ݳE�-��v�S�56cJR���1lmV��n0�[�D�'��hB����Q}�8�Z�_{�ذ�1B2U�b���7!�QN�&'�W PFa��	��R��ʤ�Z&�pA&i������s�T{��*������M��(	����%���h>����C����ޒ�q�dn���Afj�9�;'cK1L�����awy3i�4gJ+�Z�a�^��o�ފ2%��jNI�"�0i��b��M*��6y��9�Q��5�
�gŎqnS����x�M!0*p:r���s��������|v� �oUt��k:����Tj��pʵ0p�t���|?�����ɽ$|:��6ήL*��XU~N�������k5�-�ÌA�Z7���ѯȸh������Q�U�M=�*$o]��*���ը���K��b.�� �ȔȈE���7b-o�wCs��P�z��v��XG��;IL ��@aOb\,0��+�Ly9z�tjZ�v?���۸"����!3��̆���Y�lk���I��tB�M�/W,�}bJ�4=��#2.Z8Db�ar��,���P� ����A@W������3��]���W4��|:2!�Q�/Q�Ӳ��Cޣ����z�0�)��T)9���;��D�q�&h�읎"��t�ɻ���xf�܅>�}<�A��ʋc;я�b���=z�+�8���*���6	�
��0#U$����J�՘�j���a�1�V��4e�#f(�>�����o�a�j�JzD�>yqvA�{?�b���-0��4y�R��N���I�_=�Թ�U����u�tN��/��#��Ǝ��u�E� '�С|��;ω�g�R�WNE��v"i��։ѯt1V.���J�wK�/��m�؝�ꢴO��O�'țX�'-R�D�Ӽ�f>����]�Ʀ��A�V{5������Xp�*�g��lO��1�	���ܚP}�z���B[��x���K�j� �`m�� ~�wB���f1L�����nPq���d�I�jZO�d��4����3��J/T���媨2'�3�����(�ӊ~�J�u�C贋Hmqr�����:L$��W}ͱ�ვ���Uȁ<�c���VR˨�n3��4[�N?J#�!��l�P��"���a���{�W�ͫ��/�{���Q�Y�(�|&�k�h1�S����q��)�� ep5��P�w��83緒��Ѕ	qoT�C�]/v9w�K�=z�7��q�E�E�"9(�;%F���-_�@4��mR/4!�6��cD���aW��Z�p�� ��{#)�� �r�q���_~wS(��yu��ώ~�z{��_�y�@Yd+܃�rj�7�=gCZ�_g��y$qH��N����u���6��Ƣo�r-��A��X����cM�t2���:}�
I�%)����؋9���cz������h��^ݥ ���`h��{I#;e��G���������r,n���5[�_��m�W�dA�7��r��> |z�4���Z��w�:�b�%6��?I��N��p<��O��:x{��P)�"/��S�?���K�>~�3O�P�"�kmX�b ��$V� �wy�w�$S;;}��3�������R	�­9 ���-���?�=L0��ѓ�|��*�Д��3������]EqSY��|2�ar�*y�L�Yץ�S~VM������\���'�~����j����|��e[�#}�C@w@ЅzW2��,��ou��Zl쎂�A�ܧ"�����?D�����O���c�(�����.��P�N�R�{^���E�m~4D����������Z�\9T��y�_�� C ]D���Ff{�Mq���t�Ic�m˲!]G����_����X��q�
���^+�����D_C�ܲܝ��^:�������-#x��#1�x�����o��݃͞�{.���S̩�������Kü�|�G���D�G�&}��K��� �뮺��������C[	�qyY�w�
�ϝ�Vy��(Չ���=����ظ]���֜�����E/ *�9ڬ���>���m w����5Na3(5c�(�qA�OTS	�Ʀ�n
�Ī����hn*��2J�<��*A���4�w4|��R���UjfP���C��{:fA�N?CJ������,X�;������>��n���j�P����	G �&���L^G�	�~��(?�h��L�p@b�L��x�P�f���R�����MD��E��R�JH�h��~�*�TA�qϳa��ϳ�H�bWf�QATL�U7+Oah��L������:��������S���TQ�ж��7��P�T��h.C��r�&p9y�� v.���-�Q۲w��X6��G
�V�g�2�9�+�(E���c�*��F���C��B�{f�vQqv�� IR��,�!�Mg����?.m�Q��n�b�ي�.�";g�³�S�vz���bFp�'��A	=7@�G�V/6��f�ˌͽiגt����Js[�E.�k�X�`�KP�۷^��xߋ�d��1�5��'%�P~R	�o����-u�e(UP�}s�B�*�E9����;#.l�����N����]���8��RSQ��)��K6�z�����<���N���u�>L�6��6�#M�
`i,W
;/��U/PC�qW���/|v��'�����k�����d��s8;pb�1�y�K,�l�ƣ
�$���^��� )��{&=��F�_۪@t	�:mG$���s�`Fj��g湞U�T�>�<F:y�GVS�-�����.w�c�ĵ�rL+3Y�`�:n�6?���+ÿ����)%A:Y�ͣv�p<��:��mγA�KG3D=��T�P�^�H��v�2��q��M�+s����
�:7��M�w@S���u�U�R�ہ�qn�i��Z]�0��`P���~\p{����C�T1l��,���M}�F���t{�O�����uP���*p�>���tб):>�ߍUR_2�����7�(���C�~��{���VX6�"��_���������`B'�$��,e������Ұ����G9���f����"Qx?q(u! �Y�E��K&/�R��TB$~�8-8܀Fh?�E(5��|�� �yda�-4��\�ד{�aq��4"n��00�0�N�����h%�;��d5�#]e�	�\}���r�0_����H�����J�r59� 1>�X2������PjM���Y�_��_�n��Ӄ8]�G�* �0�.���N�K�# bj��Lt�ʣ%��� �
i}���p�4�}��U)\�M�(�R|��scȞ1�kZ��_?Wi׺���.V�2�յ2(���:����|f���Qo��g�l���R���G��bI ��b�0�5q��]y�V��`-P�n�>�	Β3���mA�'��U�<�)��D��������#�P$��1��H���'�a	�)�I|����cm�B��~���G_�D7W�=cU�?4�*[>!T�����%U�׳�&�|2��%�?�c����U	$�OI��{�X� �U9<j�XВ��	�27���+�,��ܛ���-DE�^����� 77\�Qr��o^c�T�fn`�M�o�mQ9H��̖J�b�(7[>HZe@w�+i�8��9��w�Lz̈y���!���lB<��%�M��&�����>�n-Hx�pIq�J��� ��#��dZ�r[oF���T��g�?�ӽ�y�K��ޠ��)XLv}$5"2�[�2R�W�m��3�K`g:܊{+ ������=�:wi!ԗ����1:�3(�Z�誃���Fa8�en��6�|� ���&&}��$��ͭ�V�?��oJv���7B�(�3�j�fm�B���B�XX��_�: :�J���G�Sw ��>��LjO���^h͞~o�i�<0>�f��(��4���y�}�,��}KA�������oe�;W[��iL�u+͛��-Z$�yc!�G~ފ�bA��&���0~�0�My�mrJlw=��q�εG@��^/�<na&�AD����4��{��x��U���B�|2_���ZT��[���S��K0=����:�y�\���B\���o	��dT^vFFeu��_e�/��2/��Akb}��;�/�LR�eG�nc��9� 8���@�J�J�#�ba�%�F��W����2���D7�W�ޚ�:����+�n]���蒹�{IЩ�ihA�a����RBT��e(^:��A�U�+�$�l���pN�&qy��dP�Է=%�٭�]@6lhҲ���6�|���>�w#�0�İd�j��z]gxS��1�KB�CJ��L���_�ff��B��xup�q_�D�-�J�M~�X�+�H@�A�n�C�"�� t&	������%����eT5�=6�Ĵ��
Ȝq0<A����wI�P2���� �a��y�)��2����"
��B�S4+Yj��L�o��N4��2ծM̤J�	��\��0��	U;M�q��8��Yo!�W��~�J4�d�>�Zs�z�ha|epL�A��|�Ǭ�Y��:��(u��	̴�2\ Zy�G�(��w�:c�f7�"o!^Ei<G<c�;�4�{��;�t�G�왕�R4��z�$���y�j�^����:t�۲Ǫ6sʆ��UH[��`<Ѣ(��#5�!�7���Y1/�H#�Z�3�/����P��d�s5���Y��E^�O|Q]���\+�������u�>!y������j��a�`7-T!h/��s���(��1t�I�5Y�[��럆-j�*Ɖ~�R�F��K+�b/�i����:6��,�J����W ��W	eQt��uC���E�k�®�^�5Զ�dn�S��l�<S���+��a!�C�;F8���� �*�EXq�0&F���`�'Y,H��.	�0iw����V���>���յ��H	�_O��V�e��B=4f�3����M��=�&�ě�� ��6��e��cfB\U��W�z�d�6�=\�6��`�b�|4~W%�W��H�'���-�E=$P����*��Ys�6k妗�p��h�Ffytew��]�A�^}L��
�t��[�.oX��l>���O�j��JF�綠����3r��֭A�o3�k�ع��#�y�D�V�Dx?�U�b0��$yP��D-���T�e��;��à�g��C��f��w��0��,~�=��N��m��Z��3#�^��`(��y�*�<Fu(�����:��z�*2�S!���y�+u[���V�vI������=���:����mN�;]v'M%�Y�9�ʠ-D�Gv�$2��;���>B�]s�@�\Һ��V/��2	"�=����W��3K��Cl�_�c��9��aLw{9��ѕ�ͷ3k?���1��N"T}*�h]y�Oɶ���r��U#K��3�x�)����Z}�9�a5�r���Nr��P�6������J�"z�PN��Z��ʇ�{!�*�Au��X��N\�t^�Y��O�ޓ��18H����������@�Yl(]�w�i���#�G�iJ�j6�0�
���#c�| Ǒ���y�U�r�)[�X����o������78�a4O����Z젇��[4�N�6�y�n�:{G�H�pf����1*^� S��5���9#���p)I��p�@$�ek
V�eXN+�`�䳄b ]2�$�g҅nEp�Ә�	�R�f��	?AЅu֞`�x�~S�3��t���]�,>����r&cm$��.X2	/H�_�*�X|i��g�4,iT�$H>����a���<�&�=�IXA���Fd��CяzžVt'����6�1�����ʜ��Fi�����'�������ڠ�����L+xIl���i���_�̲��τO���Re���B�'����]K�����ҙ�w��Qq=���fm�y��ԛŎ0!sΡzC�����7�G�"�(�^�FI����6������>w:�r�1"�u�G���rF{f���1�����2i�e�KB�R�2���n�G�)N�E�z!'����BoD����?�1��i�	�/�>~��o���T�5���u���m݉L�8��hJ��}���VUҔ�
ORz���V4�n��$�>xт����� Fy��v��:��/����z�4�b��K���C��$�� k�)��_C~�We�P|_	�z1̱C�"�ppGE`�"SJ���P��>G�0}��8����]������7���<�b�:)3�G����`�J��d!��g
eY��Y���Uk�)� �?v|���Y�J�LH?O
o��eN�ʞ$�8��dE�(!�w��K��a=��3�|m�9=�i9[��f��,���\ǚ�'W� ��H��J���6���j��+��%��nr�	bwT#13T4���%W\�'��=
��"�H��9���
�	�I����%��ѵ�H����e�q�EW��,�_���O��C��uU��>�ж��3��C��vr���q%��X��ŧk
"D�Ǎ*xi3���;��]�v$Ҡ����:.�����e�
Sp��5{��Y��g܂���S]���|W)Ԇ������S�YX��REei*��vK�;��i� �Cb��u�"�)�e������ˌZ�Iq���ҋFY��m��L�q�7�۱��7���U#�S��aH�E0���Hmp��)��n��K"`w	H���*�lK��}�����$p�*���5eLl-�����Oׅ�I�b�Z��˜.�Ⱦ:m/pI}��)����iMc+��)�Z�tϑ�)/ʿ�)�r���6�Ĩ���@�ڿ�>�]&x=���:���֊���y�&r�.P��:.�<����;��9���[�ʊ�'���`n�^�K�oP n���O���B���H� ��ɏ=}4iI�vԝӯ��r�("+��,�ֵ6J�0U���J�I��ټK�\Ѩ	?]sdSߒ�w���NK�t1+瘴o�R�ϊ����:��]hl��ˏc�zf2r-��I��1nX ����Ӗ��z�9�\˛����^!��tJ@��K�v�b��<{�Oc��s���Ce�z��)��;Ҳo��U4���rW#3��f���G��1�)����";35쯥iό5R½���'�B�V���ߗ'�i�PP��|vgE)b�w4@P#�� �����³ ��0*,Vq�ꉗ?�y��/K�������ojiM�3v��	rh����T�5�q�cs�ף���T�#=�&rp�ʎ��T��wcآҌ���$���9�b"#�+���V>�._�v��^ �ȚP "���֖�(oU��4ˤ' f�a�'�@ObP��y0?
u'Y#��R('�Y�EV�!�[p����5�P�O���УW��I�}!�AiGT��Z��3��.S���x:�ipb1k�ua;p NC$���r�:V� -���|&�i���8|��ϫ*
&x�?C�Ђ�2=@Q2S�i��K+�&&%q�z�Gw�d}t�������,P杀�(��@���
-ZX�ց�1�c���s�,���}�0!�l��R+)�����B���mNÐ.~�g�Ft>=��k��\5����Qi.VBLf����ܳ��F�NCzZx���k�����d6ʅO'�v�⩗�<�I�� ō��Κ19L�$2����,���k�6���y��I��(���#Ҫ���Mx2��Y������MOYɻ������N�<�꽧�dW�a����i�B}�k��fܱ�|	�`�Ob�	�pC��0{�cRr�P�v��/�^�SG�)���y�v��hL�TŗF��:!#څK'�TX�r�u|P�ha��Ƌ�h��d�W4+��`��&�iK�I�/= O���}Zcr�F�L>��K1�wd���'S�M\�e�K��'DR����&4��q��a5h/����{���A���f��-��s�:`QF�ƈ��62�r�P9���o�:���Jy�=� �$R�����ew��<�R�����)�Z���J=<�1��|k�����j�B<�1����5-��)��:�6�Е����~��s�3
����<!%r�a�y5�e�
�$,xc�x�������3-��*$���"��q�d���T:�ë+)(s�9���|{�<�Pc�U�ظ7񸬋��)�x��g-h����௫>\Rᦊ�ĢNwW��M���]�k�zQ6�1g�Y[���ui��t�	�^�h2����=u[��z�􉕞G.��j������� ��>t�tB.yL9/�,�ĭ��A�C�Z���ѣ�#����r)hkj�=�>��[S$�`.���Y�dI'�!���q $s1N�9�A����	�m[��H8����X��л6��p�,o�����cI����%�|��>j0��mC�����b�Tlv2s>����a	1l ��9gs����o������l�޺vr�	�|]��K�/тkMr�Ea[�m3 _���C�8)o"m�P�8����\	V����e;l�R��h�AtV7ƆE��aA�j�1����@�]���s�A�K�S�1�^�`�m�^>��.�M+��Ar2$`���1iͲ� ���M����5��G9�Q���ōC��DN5Z�#g���	�w���-E���8 Jg���4��k8�=5��=%�fK~����q_2|4(L��D�˖BʊJ���Q��,��r�Jm�ѥ�X}O��H\ۘ_hzLvT�5��֛ �]��P�<{lO��c%�B�:e�|MCf%)P�S���ڑԡ��^���_��?Z�W�����'6F�[�q݁Шd��7 ONz6�p��Y�;8Gb�����|�ՑN�ҊND?���d��֜�Op3���M�3t���aت²��!��7��4hjCC8 ��~���
&�E�it���b{��+���?ɗ(�C����,�n$.D�������^��@m'XV��#c�#4[�S���J�b�d>-N���(>$J�p���S5c�#�o`���e+��7'+i%��M���I�<��'���X��PL6����~�ޣȝ��c(.�]IzLu[��+v3-����J��$���i�.'� O'ْ%o��2�T*h�$�U�{�s��Jy+?缓{��I5A��I��0�c�R�]DK�P�"�ٔ�I��0�Y2�[�u��:��I.0�.�rU�Y1��)�~�f��!&\ҖZ�����G�g���g�9[��a׭����Ԡ����Zv9I͏��a��F����A|~�rd$� ��^vب�g���Kٹ��J�a���F�W]�t�R:��sc9,gvb� vd��s�����I�)ET���I}h��d���*����X�w�V'ls�2��w#ۋFGs	0��r����ﰞ��V(���r���h�V���!/ɐ�vcz�ɘ�*�b��������T�F��DΟs/?��p\��[yr9Q�*������KE8�ceM�;>��'D-��a�C����jW%aq��j�K*]l����X^s'����*���<B;E�̤�;�֙�C35Y�S��JaB&�+�e��I�:�9�r.lo�����3�ԎQi������҇�L^����D��"~:�H4u���)��Z�1}��'��Ks\$��M�<�5\��T3x�i��G*Q�F�[�y�NJ�F���+��mf�hTr�Lb]����4K��U��!�gK�3eT[��}1c��cS꾊Ғ���S���"�*�-�opE���>�fj�/l��4�����*�,�<v�ϚKّ��i��H�Q�Y�ϗ�]1�d�r�b�'�0����bH�=��_�C*����J���?́XW�l#0c�rC���T3�gr��:j>�ӥ[���������M��x�Ωbg��+ ��]�%�@	�/1����W\&��⮃V�S^���>&<v��V#��P`
o�ڱ	j��}��$m�^��i9?מ�����!�c�/>�mp|ڠA��g������3�DG��rN�`ɋ���c3��+-�7(�	�U+g>� ƟrR�(��3��Lb�^o��
\ј~2wIqK��Jib#�uu����Uċ�凜�
��8�0��c2�Z&x������zLT���]�ֵ�
���4w���=�� rڗG�q����s�{���n��L���b��=o�=�]�L���hc��Ɖ[k����Ub�D5�����筧�)�W��9��@a��J���o
EB.����'�u���>��������%}U�O9�𶊃�:�H�0-S��S;��c�aِ�<A����X߅RG�[�֠���1�6��Ȗ�6H
�j��Ӽ�L?|����f��iDd� �a��E�$��+P�>���XFMuM��2��f
Q��:[��-���~i�jc�;�t�R�ONZ��m��H�\X
�2���7:i{�77�l{�_�S%�\�3�Ȱۥ,3zJ�!c���7�8���=�yoA��ZM����"］��.��H���-�����^�R���|q�/QSi�x'+4�S��<������ܓZݑ�]�T�����\e���j	��y5���(��f<1�FmK��͕t<�YqY��v���ߧ
�YˠZn���]&��XOZBi�d�I2�����p����C�j>οX|�)�i���u*�_�����h��XJIXUb��r�M�T��FA}�8�
Xs����1�Ijt4���� �񁄽�MY�T��>爖l[���x�9`��,��idi�G��4L���;�Y�9���oH��	"C�~`���*����j�D��y���et�a�U�J�~�8G�R�k�q�}���� �Y-5J?]��ߪ"��;ѫn���L���l�o���r�5��ߔx������=��h{׏l�ڴ�����{Ս�!/���'�Xq��V��۫�M��wv����1������TdO�$y~��b����}��X�}��� �x�.���A�_H"��\��'����5A�'3(�����Ow\�g���WMu�N~����fv:�ѢJ���]qm36|S^�ol��]sS�\m�峽�J�c:Ɲl`Č*5t�X=�Z�X2�X�m�͌��8��'s+g,U|��q�.��B�/��㲿��P��������|��(./O�H[�w�BMX����]�*-��^�����;��|<�uB!�H?�����j�p@�}��"}�*���4��N��T5�
:s		�Dȳ��I�IS�T�#�Iy�I�1O�5����Ro�gCF�
��g�Nb�� ���&s��G���ץi�F������PN��	����)�b�������WS�����ScO�n�@dw8-�Fwe=M�tp���|�5jFN~��AA������Had\�k���C�����U�F��h	[z5���N����պ�Y֒7E�eW��f�0��@�tk!�ة��"1�����xm�2�H���f�Β��O8�\��(�Ő@=a
�!����X�
�͸�����~�V��,$�wR@���z��� �1���T�*>��J|d�4Z�����a;R��Q�n��BA+V�]Ҳ5Q+���:���AG�?���s���]�S���U��=ļr����ޣ�|�ǾF��$;�T��k��G��.���/�=C\�9P������Z�W�@ �7���x��#"�C�C��q_Xg��觬����ܦ2z�})w�����-[��eC180`IM轔kXF���L�4�c��ȝpg<�$���I>��;u�����o�m._��q�Ķ�������v�= �}�v��Ku�tX�1&��j66&U ��c���<5�=p����Ύ�Q��qt�\�o���в$v�1�41pd�2ݝ��T��:��"r��Ͳ�װ\U,��dQ�P*?Utl��xu��
��/*����+r�,���UOaȠ2�*_^;�@'���� o硘��^��d{J=��b��#W��Hd:��k5���,���vE�
�°��1�����	�TY�|g��sC�9CJΠB��u�j�q5S�Y�*|���j����hY��L�����}d]����� "�L�� 5DT�2��.NǏ]�y��Ou�q�J���LP
^�zr��&p6��Mk���v�j������j�lO~{f̢��x�11�up�]ȻD�'����"��k�47K`��	؊��I��%;�3 ���iY�~X�m4"�iCY�O��O7nao^��ޤ��E<��Yǵ�^��{Ӊ<�Z�	
l�RU���Ry3�f]
�6��,��>-�RƆ��5��Bs�u�/G}��z�&ǗyYT��Zr���#�/J��a�d�����2���j�'�4�J@
�j=��L���VM�\4�!-�[_���f�	)���@|D\�H!(�m�����0����Ũ�����~T���4y<>�f�O/�.}@)<('�(�mQM6ܾ|G���{�����<���]�_�mK [m-�}��:����^�]#��j����Oq�'�Kd,��I�,�!��}kf�)�d�@�zl"�w���{�ͭ��*���V4M�g %J�o���\�W�a��Xqn��`l"��5�$j#K/���n�e���\A{c�����ӱ�}��1C	�6���bB����2U��
���G�F)�� ��Z�xUY�k"��R�Ɵ�`nU�7�5��S�����z�hC/�����i�����I��R�ba$�o	?��q��C�GX�ږHB%�؀�+
���@�����;�2�ہ�m��HA9&��2�&�M�ρR�ڄ��NaE9�K�0�����p��XU�:�Wi�*1[
D�k��&ߨ��R�{�R_�xj]F�F��c�((&�L��F�������Aw����1����L�����k�[�(��q&8�K��~�O5��U���?p^�:[�Ŀ��S�&k4���(�M�׮���0n� ������e�g�1�i�ᐬ���n�`1�;(�S<tH@Ҵ=e~r���on��$�ilw�P!����u@�Ĥ��#gE�N=F����|�:_c� e���J�܁�Ub�ڀ����sg�=i��� �f�d^ ���9���b�|R��9{�RL��f�w�A,�Ђ��	~���X�D1� �3���o��"9Y:>S6��5ڸ���! 5��%���]8��tp��
+~��_f��)�o�>��7���읱!G"#�z(�p�U`֪o�\8a���Su!�Xiخ��4#[S�5���>��|��	�.H���.l?}i����]�ds�6/��jmoq�P�����e�K�	7ys�>V��zs������~��.�gvHm�n�:fw63n�㡷X�v=���&R�Iz%�b/*�OI��g���J|�z��Z�Ds!��$	������3�L��rn�_P+������&ܠ��c}�y80�ߣ�iӠ���������S�0�B��?��hW�Š��%�ś�%�~�5��|���Z!�B=�Y �� ��_��1������iq�_s$N?����w��3�S��-R��v6`^ֹ�2�͉��<�j)	v��m��	gW3K�m����3��ےP�IAJU��R3�	�sO�F�}0+"f!��c�.�;���EP@
�(H�sO#�	�A	d�[�����u��$��`�O��4��>-+����w���>��m�҃j3���j(euiE�D�ɯ�������dzlB;�^/*�.���:24��"İi�b�x��z�2�QG�4���9t�|���x�ba�o�=��Ҋ�Ӹη;�S�z��F��(e�|��^�x�R����,����<�� �..$�
/�L����4Z�6��sȩu�� X���?�zD�X��.9�r�h�������L(�D&?�4*t� �1uWv��t1���0Bf����E��1��~,���)�]J�)�<j�N>,��(�hU�ds�ܝ�eP@D�s8α�tzc)s�y'S�Ho�mSltw��Tm���<~F�gƿT�w*��gXۭZ�������l��\���'ȝ-ǀ}׹�����)�q��7���<��!m�d�k�(��,�dp�*4�t,<�]M�͛f}�ua��P�K�!�@�[�[�'����}*H�z���w'�f��M�at�YH���+�fNY�чdBϜ��*�
�<'�n{ȉ����l0z��!q��^)�����bW��4\��򴮗��$;z�Jk�l*���8wܣ�.���
����s+��E�U|����U/���^z�r'��y�� U��\gq�z���1k���\����	���ت*�������+2I����j=�~�6	&	-\���1\��(m��(��0��
1pA�ˋJ�W 5��JW����uQ�D�|Ud�+�ax�0��Z�"f��A3�c�W+�#��yү':�Z-V����>�����a��l�A�aV�����mX��U����|��J���p��y Ht��EA_Wa�L����9>��;��a�7#�4/`p9'�]��uOÑ0�j�4��;��e {���j0�>y`�0��8�Nm� �b�o�؋�@v��@h�s���1�캁"�����{B���BR��.��JY���&���$=s���n����k��GK-���&|��<ux��ڽ,&��,�.���Cdg/<���t�;xq�h�P#פ����Tv ���%��.��wQx(�¬�c����";㸞�v�"�a�|m����跉U7��K(�g�h���5V6�y�Lg+�1R}�|�Zq5/�#r��W�F/fO�L����v,����s�ð�Xʗ��9�Jݟ�[�^��.�Hsq��9� x���M���0%�IX����ի���{\�s��h"�EE�܁�Z���|F��f|��K9ݟ�M��!(;�lW���Xt���2R�A����tz�Zvycr�tC	R�T� a%�r���{΀ x����s�K!r[V�b�0�Å���ӷ��IQh�ڽ��l�+�"�v����0���#s�,#��9�@�{,4V���^գU�&5�Ȉx�8���[Ve���K7��i9��p.�qg�h)�����c�Ñ/j��]�3��?�K)8�0z�͘�݊��7�a��K��wt-� �w��,X�FaNu�|�����mR��M ���A�1r������%J&j���g��g5N�M�ynT}ηm^�	FeW��~-B���y3}[�d�P�I'�S(ɴ� ��� *����N^L?��[���wa*-��t9�\p����@������𑸜i'e��x*��%P���u��'�v�7�#��1?V�&?0�/��E���DL�pv�h��I��#���5�.K1D^�By�iz���o���@T�K
5�3.t$v��=��ön�w�h�����[�8��i$����jlh�;]�o�5b��$p`/8�df@��n��4�վt�\�� �S'4δ�M^<k��C�`u��__|�|�b�wݖ�2��6=�n��͠I�3�����͖=��nɗ����Cʹ�U�a�f�����<2��p0b�H�3��Ebvoc�^�&�u\)��J]��u	�����S�R�O�g���-���tq�����,u�0Z���,2����z�\%;�A��lX�K&��mdC(@ۋ��m�P��4��3`�w3;J����ML��Y����Hp? 1Āz�����cgQ<
.�zM��&�	s�����/G���S�]���͈����צ�G��RǠ��YN7�C�콹 tV��2Y;2L��^7��*�o/�ggE����֔ÃU�Ì�p<�JW��)�i���f:~v8I_�hR���җtC�ac�	w��7%�je����zr֖|����ٻZ8�p��u�����nwv;+t�f�^ؚz!
����}�.ʌh��竚����O��B�W����Ao
�쌇셂ݚ,c/��=5�pN(��Ů��{hb!��aFz�� ���x�'��6�p���_Q��X�������OA��WC�0�j]��bW2��HP�3�1 0g�~"o�|Y�V�$п��ژP��cc�`)��ZKS;�lq���:���*B��b��
��j|� _��X�@ủ��Z~q�6�3��2#y����˸`�b�r.u�� �m�U����M��_@�h�mgς��QM^�(5���U��(̂j�`W�@A��tI��P^Ȳ��q�j$H$?�2���׭V�G��〭!U��"���&9=Q<�ۨv��V�>ֱ�f��!q>T����� �)jDSq��}�_1�gU8ѕK�)(����!��w��ôUA�p��4�2�jya�lQO�/�"|f���8��S�4�ub{�b�5���4f�C���in������(NՏ���Zw�.�G���lÃ��Ԣ6�&��!!������y}�Ӡ}��c�Q�ri�(�I��E�.o�����ٖ�?xedk8_�3����OXe�l�s2����� ��֘8����V�`�A��ŏVs\��X�A�`��ް��0�}���@*�e}�c$2V7J�u6���ç���W��6�~�6�ż'�ph����zqgo��c��>�o=�>9�U��lk""���a�&�\J��N�#�@�Ӕ����u΀��32�i^GI:ܩ������đ�����\�9U8g�n�+N��Z���/c g�CE@�C-�yH�T�yI7 Q����Tc!N�åpm���w<�&5D`B��C�tU��*WQ���hF�1ۿ�zPLs�w9x��8PIx��)g5��D��q��J����KŲ��>�%�n���;��E����b	1x7�tw9O<��|�t��]pY��q���[�� ;�XTiH���"�r^Ӽ�����Wt��;��A���	(�2A��bo��X��|(�(�H�A;�$���$gwe�����8	5e��L���q�GBV(	
��h�����.�k<�T���eZ�v�햴�#����H �/)lUY��б�~5-N�G���@^��=E�?=��4�g}R�����|�����eJ�8[�������s��1�ϕ��ZZ����>{�-*�ѯ[����8c��w�G�E}p�S�8��_[珴?�m� �.�T�B ^+1�A��/��Hn7��)��[	K����G?�r��n�:8�6>�2�m|N:vhȢ�^�J�(���4C����I%l��,��pF:.�q�;X���]��v(K�g�����xW��	����9�5ƅ�*��=�*��ʻ��O];� (Nk�j�4�?�&�,���I=~�7F�Ŋ�|��T���YG;���6�ޱ�)�wH���fp���!�
Kn ��ܪk-V�m��e֞٥�	<R�P�ss���̠���-\�h��%{<�n�ך�D�,�vwŗ8�c?� r�v��S��$>�����\C��đ�W��� &��ɤ'h�*��ˠ����+f�a�~
F��!gC��	0���spn�8���wV����p��%�:�F�g�Q�vy���J94��f�fX����ؑ��ae�N��2PHUb1�D}���e�<zM;z�$u=8��E7��ru]�����S�3E>��We�e����g�H�i�C����+�Y�uࢊQ�,�e�>���T�)���>�Ķ�=��GlP����2=;�*LK�C�^��|�r<>��N��B:J$�j�:�"RTd���x�('�JuLv#bs�ءk�H,�ı���U[휾����!��l$N�E��q(iP�^b�U���l]
]����4>�O2�=֦�gUFo� [%��r�5�J�֯T�~�������(p?��jZ�傠.߭)N���T���i ��J�A�֛f%��P�e�m�ـ�7�U��s�I��Y]:���^]X�}����N�9h�rm7�e2��Ji��ؙ��*�::�oH��<�+��yb��V|,�MXJZ�n����nFܱ���_�bt��vU�t>2 �TI���˽�ߞ�O~�ɓ�@U�F+ټ�RR9`VC1l�CS8��ڰ�����n<`���G�eҦ���%T��hx�oGsI��^5N��?��G��=���n>��FȎVFG�ifZr��S	���c�T�O�����|a��L2�7n�1�g)҇��=���<����z�F|/0��cO�BI��~>�=V��ΰ_�I��V/���5(����U�_萢����	�b�L|�zʨ&����?g��:�C�|6�b\ c�q:9uߚ��++g�o���ܣ�}��g��� t��Q�C�������JtR����3�0-U�+��C=��Q��u,%-k��Q�Y��|a�~��y
䋳CtV �t�!G%BJ������W��4^t�\H���M�;��?�#Xđ����.�@���PӋ�;�F�o�R�����6�S�������$ZZ�<^6R�b�y��:�ɕ�@4[��k=��%�o4.�v������y����e�&����u����A��1"[g^��=����I�{��ʹ8��!Y�����7y���0����A2d�v��a"l�����$w���Q��yv{�oԕ���aG�-����a pOm�4�����&�cZ���Ԡ�D0.x,�9��1YB�t۟�z�����cj��BX�7�K/���=�߃��ܽ=~���Zq�
@k�Wu@�L=��0�o�Q9b��OQ�1��	\)��n���v�`��-k��e�i�B����Lk��f-`t���Rf"�����V�DWK�G&8al1ݵ	>�q�U��(8=P��x`s�3{�?h}����?�*+�R��6�+8�?�֔Oiik���h
̷�{$@�6�f�C�!W�>�Ar�1�;���ͥ	F!1(�sQٰ�2�1�/�
a�����gWO������/hW�{Qж+�-	�B��>�9@��Yr��n-�E���Ơ�ɼ�&,U'rv��ӏ)D"X�z�F���+V�I\������e������Q��:ȩL������?�}��6Ӭ6��� ���Y��<9�5%W�eu�M����[�+4rYN�Gx��lsԅI9�'���1�_}N�3���7��a�3��3��m��Ld|���L����)��Mwӽ���U�c�M��M�>L�	ĸO;��DX����~����6�Z_�J�w�)=�{a�9}���&��%���p�`�S�)�b�x��:C���P����-t���W�UŸ�dn����?�u��0�+��:�qk˷ΐ�(�2Y�,�y$�R0q� ��vG^�w��2�m�I��2��-}�ŝ�����Mӗ��a��^�B��k��1�����\��X��?ogST��H�m*���
L��T0���S�[e=6��ɲRMp�sP�ҟ羯���)��?��#�23�NB��fj�T��y��^mT�?�[�e���� ��
���!o��{T��_���y��b��ct��8�����J��uk�y��!ꦚ��H_V���x3�uj��u��VW�>!���~���M�	5v���$�l!���@�)�`����OF����A�m8Kr9$	G���j�ڨ��l�~���{
T�U����3��]X���G��SH�`�p����Q��%1i_�Kb̻��]��W�Ŕ���:�f�Pg���o-<S?���}K3��r`�x&�w��?��'��4re��[�f1����	*x��<��?����	�"���#�aHe�q���aL��S�ك��$l�g������I���~�FiP"�dw�
���C�Pr�a�&&�������S�7��w��4� �a;r�p"����N�j{�����Өᰚ���A���1����bR��i��_��~N��+�Sb>ZT7�O���#%�ߓ+��dM��T�VeR�qN�IŢ�TdYC���0H-2�����rr>1u��,�:\?����0~pG�Z��	h����Y�b﷣ra��1 ]��P�ޝ�j�6g�����D0(}._r�u�O�W�b�i��&.���!ǡ���Ҵ�+��I
Al���6?C�W���"�-�3�����˷iT�+1J�a-�մ�i�Y\)��͌.�);�N��~� ;� �����������P6��'B����Qsr���g�L�L��R�ݿ�MɄ���^/�9sm��d�f�&������\[�Nӓ�D�L���5F�;�mV���k(g��ɇ������*���r����A���a;�<�gE��U!`�$yTk���3ꍏY�y*/���ѡ�=C��2��o�U�B�3�ǖ��$W�l܂S�b���L.|����"#��4_�w��ѕ�Ү�b.�R�T-̖g���,�Gӧ��@�r")|��1)TJBJ<K�iH�MJB���W�ʛ�����&(�4ȃ�(�=�Y��)�{�ہ�fr��J���P}u�N�CT�sE�O'\5����a���������Y�s�铹��Cy7 ��/"���`ำ�6_Q�*�vl���3T���HjEL��n���K�]T�~���m�m���]������W�f��=��P��<���y+S�ҁ�{_q�UQP��}8�
����,�/7���?r2����1 M��ɎNgkߠ& ��0x%�rF�w4:Ϝ%���z4j� ��nI�Za3q=A��1`O'��I�inG-��T����9�5�'�7s|o˗�⚗d�"��ox�;|���{�6O!޶D/Ǘ#�"3`;���V���cQ���yz��bh���b/�JJ���>�X�f������qM��[��`��3j@g�jVp�mBQ�ڧ�`>��R%WWy�`̪��ig����}a�Z슑�A8L��*Y�����*&�p8�;uu���2�~Dw+݋bjI������p�%bz����P"�v�\�9B��҉��N$�{Sؠ�dYOu�����Z�/(��(���Z���w�&�J�wr�|b���,ǝ l/�$5u�h�NNHO����A�V!�3�a�������?L�غ�E <������9�-�Xq�ڰ˳ �pΛ��^�-6��m�.˜�)�=�ڬp�A^
J�u�ӫw���/B���XjmO����ï�@p���w���7G�R6E��0%$�n�nJ7dFmچ��ĨʀkwyA>5�!0�W/	�'�ճU=Zg��?ؐ"�ؖ�H��4ʦg!�:ڰ��E7l�J-R�=�I��?5
xZ���}sE�"��	 ���-$���/��o'�!��B���xew�}��p�B��r/�	(S�h���9Ž�.K?������s�!��7!қ�����7ySCy֔���q^%����/ԃ�ny7!�Ktfla�R���߰ĻT��3PN��r�Q30!����"�$��*U���'`�M�Z�o�������c����ȉ��0��m�F&�N��32�^x[���3b�e�G�۟=1�+LN�����5C�@�-�P~�z���y0�󨘵���Ê�@F�����+5F�&#�*!�S���B$-��x$���Rv����U���YK%��B��0�S��HA�mg�C$cT:N����\��/3CirF魛X�#�d)�47�I}o�4�O�U��,�	���=�[^�k_�1�5c�]�/ժ��p�C�!-`�$!u�1Z�@~��t� ��Ý
o��1[9J���n\���<��`ʠ�k�E�/��&-�?�J�Ǡ�`1=R�|�ڵk���zn���ɀn�&Rx�o���o<0���b���=��i%�Ǖ�kˊ�lo2%_���ǦWc�p[_�����IbN�0	|F"D("�Q�1�g�v`$ٖ��T�9�q޽8?�ETH����
D������`$,��`}��2&1RL��3ỉx��$�Dעb�)D>*)��p,�v�ӎ̎)�\poZ�O�$U(�F��j�5V�hv¸����C��ޮ��O��C��$k�Q�K4�!;�qN�/�y�5��#�v�q� �$��m��������C��%T1��/5��0զCB��ZU��"!hr�7�s�B(����K�`&G^0u�]��<cw*����n;�"�x��9���_��N��
dCg�,B4�����.�m�����X��F�#�-F��e�Z���'���쯳��~�p��}N���y�M#��!�"�v�P�ZS+�RH݆V(���#����C�E��q����w{�,l�:<�Jc� ������0=�~?Hͭ���z���n.� iB�e��1�k�����9��.	��a=��C2��]հ%r_��Q��+d �ib=1�=�n�`��ԭE�(��Q���ߵ�'�7Y*.���咱-Wx��l5?�5�R�r|TZv`]�0GV9m.<��s��
eI*n,�LI̚s�%�+Dij��8�.;v�
O�FZ
�:��ip��)��bm���<����ж��W��c��f`�UG�+�(9�r�"��n$׵{j��T�W!Į-.KL�Э��!C<^B=v��?<G��z��a�9��.�C^[}J%O`��JI�� ��J�)4
�4[�1˩�1J���L��֌RXos��nF�g˨���}�/̗�)g����H���SML?�N�ePpks��mW~hƻd���L8�`��ig�G%L��K��*��7����`���㷯��ۦ�5X�-��7���o5��r�Z��u�K�m��!�R���6�B���o{G$�Â��e�eB��W������hh����5^<q�E}�^�뛟�L̪���rZ�+:JrV5O1bx����m��DT>]e������3�a�M|B &�yNm_Y@�z�LP����s�^'��NԤs/x��Ge�jY9qXڌ��w��4�%Զ�������.�K��[T�g��Ek�{�	���u�Ѐ�X��:'�$C:����Ys*r+e#�� ? ePoj[k��;\�a�4�0�#��ˣhp�^l�`9C�C�Qz[�������S�h>��%�"�E��q���y��רJ4������H�O�(�𬑪vl[?Y��pR6�$���a��cR�)S�?�Ҝ��n��E����dPEA54���(5�t���ia�2�K�t�0��K%��k��Ӻ�s��x/^����B҇��Ғw���Y񕩏m�ROᄡE
��k��k�:7�۱ʛ�0�|�,̀�+�&�;��A��P��n�9Qn�� M؀��@u���Ĝ�q�?_@Z��L��NA�� �t7b�3�%@a��S�>�e�I�:qk�i��,��˄�v"������pA�x�S����޸u�L�A�M�3] �sZ���VFU�>ҨXD��/d}u�)����_�$�K`j��:���Gz�uk5����"�R��$"�|_h~�M3�+�?T��>�C�|���\d�2ؽzĴUq��}<?0��F�n7-qc*�����+��	�7xba��1a��~�w��2�(PH������O*��SLe{��^f�.�+�R�K��MƇ�3
����hK �����θ�����8c�9-�XeX���Яϯ�:)��4��+.e�{\L����v�	]:�?�K��UB�w���y�M3��s�>L&eH�i��@|X��p��<mƦ`��x9a�0��l�����yL��l��h��P���#����i1����6�9{:����T�8��0� ���;���$d�&�o��F��X�ŒN����oM��dX(�jΓ�%��Th
,���B�4�Z��ը��L�B�z��-����}b~)A {�_��mB��c��^M�c؟#!˅d����A�hX$�2�"պv=�G	���1Ń?*�ɖ�(��D�f� ��fZ�⧪.�P������mg�a�l,����S��}�)3�?k��<6,0�l4�l�G#�g�(��D�Xx�F�����:�fp����(�ENNk������PSQ��op�������5�h�t��f�,����}:�]�J�D��L�j�8;��nm�dc�ʞ�<\n���6K�jŁ��z]��_�E��tmW�0�\�������v��Q�ƒ�	@�uѮ\�7k��Ú�
�mW��E�	0Z#���x�ĸ�ʰ�8��-��&�{�,���٘�7Ɇ���p���#�R2k[�4��jߒ�	e�x$��O6X����w�E�xF!
A_��'��ڣ��|)pl���ѼGӷ=0aB$�D@ˆ����W>~�3l�9僧�߈�Z���Y�#���55��q�c���Y����@ݮ��3�Pw���@�9H�x�a���ik�C�mNP�ʻ�sgsQ)��'s�v�U濂�h��#��?TWi���	������?ל�r	��Vj$�U߈���ɹ�?�rD�3�#����Lpj��R�\q["n@k��4�3\�B��6�I��->1a�k��BN�ts�q�̸��T�]�W��؜��@*XE��&�S^J#���.`.��(|�P���$Mf���o�����H3�w�B/zdh	��bB/�mm�.A	QE�G���'��T��=���r�'�Z]dq�e2����7���g*����a��6PƤ�8M��,U�D�V�j.���8sLV�*�g�/^L�JN�x���vo���a��t�{�����+!�W(���	,�Q
�A7l�sdR�s�x�J��0�����W���H��L�,oV]g��~fu�{,�7�6D<�/u���L≷H\�����ٓ!�	�=&m�g5g��>��&;����\<ɾí|�ľ@E���� �q��t��1z���2ل7B> T�%���'r�Ɔw��ؚ�vh�9�x��������K�܌o8�)�U�&�5�ew�LT���L|��+5��~}���C۹���.�\��H�'�=~<��U�q�%�mmh7����S�Rr���BKn�(~*�>9&�6uK2����-�f�0����T�;���|3?g�"=�r|r"+[y�7S�]l�F���т�"o�e�#&���"�ʍD֎eE�Wz�x}���O耢���i�~sx��>)��,X?$Y�ѝ����4���(g%l"B�����@���-�D�⁤�x'�i�1��?H]"K�`���
��_C[-0auQ\�ڭ�J�U[M&�I� �˗�}���\&ĕ��O�k5|���ћ��/�[�Y��|-u$DLv���?�a�9O��.p2� I��s^cF�a����C �C�L�*:�8�2;l�);z�����P�Me5G�{~:A�{�n�K�Pﰔ�?�q
hHmPz�wX��1:|@|0���}���&��1d²[!Td�L �̝/@�<�S���~ļN�����XQ�>�0K�����/UU���"#�5h�I,֘Ew'PY��j�"I�H�t�)��,l��.�,ѻ����=�������[c�F�MV%�¦髊�b�=&��E�	��{o��{���)֔�!�x6+���B��b�����5�AMLr��~��W��i�4+L&wV��Ĉ8���1������ޣ|?���ǔ��b29��	Ʊ�0@ajT
7��$�nރz3�[<W���rU�/e��ww�]����|�G@��o�h�O�Ѩw�sk�%���J��	�3"l�9��M�2҆}����G��bO���<��p�&�KDs�{S���܋�ȫ%w6{kY�P���S�d��C���6���]�0֬�V#� ������ub�0�&���a۠���ag���W�?ɷ�T����qh�b����୛�V���4s����-n��栤�cO}���Wz�h���D�lzS�v�'�r&�7:
oƑ�36����B��m�:�2�4?�D���lxf6B�>M%�
���,�Ӽ��^����9��*�u�Xl۸Nm��$�S�_�K��V�Q:�UZ;S-���"���qX=�������'��8�\o�U�๭�na+C�a��a�;# �]�yRg=��&�B|�kmU��X¤e��x�fyL�@�"�$�//;�;���c[�������A�5#3B��W6�ΉY������P�ׇA��Z���}:����\�H+��yH
�s���D�9y�
-�$���J�[�_Mm����-52)��������J�±i���&!Cؠ��0��������E1u�K����ef���NQ�����L?�Z���>��*�1^1������٣3C�Ѩ�l�c8�[����+���p��O�<�hwA5����T�]�#��5ѯ�լ���r��Gnt���C�o��.יִehk0�n��Z�z���]y��&L�O��=.�}���u]����V�<�6s'����0�G��`���I�NN������ �u�����_S�W��M��f�i��kE-�L�4W�s/���o4ׯ���꫎��s�bގ����ݡ��I٩𛝔�����-c*#���U}�BQ�v��Vx��"����@v�i�&��oA�*϶>D�C�NN����[)=�m߃s�ڞ��R-�c���ZЦ�M�+�ن�u�*�f���2\\»�'y�¡i�3�A�m�H춝��j��F	j�K����˪�n����^�Q��̲ÈfKb��ߟ�7Y�L@��e��pG�}�����@�Y�S�f�YՒ�"P�˯"!�ыU��$��TVp=�;�Z��%Fg�-%�ށ�+����,����x-���dF4��I��E;���5:�M��o��bp��8Vw����D���3����6��T���_��%e�R)O����K^�J��M��2M9N��p�.�:� �m>O�ٮݒ*��})�6�S�GD�p��h�����%
B���5.�S�}�~�5�6{N逃d��C<��
�N<����)`�"�c;��ŵ~�e]�����n,o�ﵞ�NO����q����3�q�m�-{n�y2�V���Ok��!|P2W�@�l� �8��@(��QWi[L�~�u���]�bٖ��@�[�v㠧K;�