��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jåا{�\�u�?߷�dn@6�zf��r������;$���K_��+�i��(���ذ|6b���F��eP��cт_�z%�f��/'�yU;�+��R����}���s�y��V����Ka��/9��(�!�VKKZ"���H<��Xk�Q�Ipi&��ܚ�_m7�����Y�1ST+�UMm���-ٶ�@D��Hn�w��UeN�V��%�d ���������}��eY�?!]�\;tPtÎ�����+keu�6\�ZiK�!�];|S��&��X���ͼ�V�R�K�gڇ�7K����x��c�Ň� Ŀ�"�4<�j*.z�E���~����������t�&~`�6�T�
��,,ȡA�$�Bf x�� �$[p�8�X���U폧�oA��?��DK�<��q6sĶ�s�t��DU��0FK��ee���Ȕcm�7�D�3����������H�A%�¼�ժ�Y�������%ω&^o���D�!ض�j繜?��T��� @����)V��C¾R&9�ȋ�6Y.�Q)�k.���ʹ�/���4��	��V(�ŭ����3��!��3}t7��G�!5�}�;��Gsc�{���_٘j��L~���K�Jsg�6�LG�%���a����qFe�,]�c֖5J�t��-���Db$� ��fb�V|X(B�x�h�T�����lVE���$�l�wNag�z�_�B&gh'D�P�:=h;�'TQk�S]PC�U������<����HO�h�ٹZ��,x��qQ螖'��M��&G������<!b\��b:I��b�M��{�K�|�k�P|�0<���D^]F��`� ��JD�l����)h�~Fˁ-ǘF��k�C a6^,�w-��L�Z)���Eo#m���A�,Ҳ�y��O܈k�&��˳�H�qĸ��H!*({y�G�5�s�d��B��7�pE��B6s�9"T�1�[�d7z�FX�~Ŋ�e���y�GG��H�
��F�=A9Ȩu�DJ�o�Y#�#��C�j�p�@�4��ɋ�m´�d��@~��`0��<�SM7%����I�UEM�����%�0k���C8A_.Hw�l���kd�&Y�u��J�%t�[�D0
�:���'��k��k��a�J8dPv�p��\���+e{s��cx��2�bB�1���v�EՏ���<i�����V�{�� !WL��G8<:�9/+�N���L-0GH��v���3���,e�U<'
�B�o� W������2�蠹3Y(�R���`/�!<Q��0IQعb[߂ �20�u��f���(z97,/��>�^n�{ ���O.G�4���אҀƈ=�2@�&;�L|X�������I�IXy�݅y� ����Y��R��bJ�&v�`}������R!�ZR��G�U��Ў�c����ٙ��&JciYRM���U��h����bL�-30��Z���\W��k.���*���*�y�%C���+]蜌r�Β(��2����b�|$㾊<ڦXA��|�H�;t�)L_��W�2�/��D	yuҪ���H��u��M5K���w���s&:�t����	"#��L+$�[q��-J\<����I�� $Xņ�:'6��+a�.7�]��C('آg�7���#��?����Y|1]����Q]��w9�/�e��o^�}�IMP�n��e�$�Wλ=,~̼���KWN��e�*�~K��  �0��M��dU�u�s
^��Ǫ����A#�`��iʎD���d���5o2+����A�*)a��/��m�P��K.+!��~������N5#t {-�i.��*����e���Vz��H��W�)Kv�Ub�A��0Ee.~E�	k!(ug���R˫�m�<�:.
~f�O�v���*�aD��l�`|vP��|Z}G���."y>w˅W	�?��	�=9���.�yӄy��ܗ0l�6w��Gta�{P�|w��(8�\���X�@��$�T4=��(Ot�!�p����6Πp��BS���h�U�o�(����U `�x2D�o~�^��F
#{";������,� ���G��jBd�ģ���O��%ԡ.M��5au�q�t��%d�n�� 1�P��#�~�@�m[F*��`ګ~�Ȝ<qd����|���7;�p����G�b*s7����I��e4���"N�c/�?3�c����M�+��6�黠�g��t|�7@4������]x��"�n�ў����X�_P0?���C����Die�AΚa{����(Ij�_A�R�9�;����P�՛�n񐪑��K�o��b�iGCc�)�v�&�=о�m1(�^v�2rz'zG~,�$i�R�L�E�x����Q��ke�Ž�PJ�.�X-E��^�r��s`�a�tZ{$�-��)��ۘt���k5��D�*h�J2���i!�	 [��3���Q��|b5@�A\N�����u��kmz�%9�����4�M e�S�A�[�n��
@=��'R�)u&9AО�~�	�J����א|�0e�Fr��vr���Zꇔ���X��uo�8`��Ƥ�(0�]��r�y�V�B�4��:�"5ڿk��xO������@4��`%�k�Xxx�R�� ˱�����V	pCIݴ�'�Va���6OkKyt�n$�g��W��a~��ާ�.֛��͈~2)�:lM3�U{cg �
L���A\�g�\�>�D䤭��b:��Ji�� ��??�#T�:F>���W�]��:�����L�����
��A��ቹ@cB�s�����`M���Q_n�v��B�a�f�1~�t��R�"�uM16�h�ft>Ć��8j{����~^`����.�d?C[�^7�(�'����LЙ߯Ͽ��3:�	�
�2,�A�gw2(���8��r\��!|p�m!�%.x�hU�m'�����s߷�%���!Y{v?*�.9�S8����6_�iYD�����0�C�X��R�9��_�����J%C�Oq�|cK�c�����Dف����20=��n.�Q�8~Y� 6��l�~��\w��0 l~;�FPwt��z2[����W�*VBh�Pa��x�\�f��I��Җ�V_���m�1T8�D�m^b�dt�%^b�"[�D
zO#|Z�~V��2I#�����e�"0 :�z2�e��-�������:B��"5Iܘet)�&i%YYZM7'Se#�w�����VpD;��"c~��4ƵTR��r����J��ҖUe~G���6��G�C�R/W3�teZ��J`��(��^C��Y��V�Y�&�c�P˃�ܨΏ� �J.�|A7?��u�9X��xU ~�4a�c1��	���$�FR�Xd�O�a����s�_���L�/��m����a��[� ?���X����a��gm��:������,�pk�:��G�M���x�Fq���	;����E��)N�Yq��P�C�"/��-���DJ����G Ҫ�d� wa5&�t�]J�`�� (�/���ޘ��d���S�p-�6��`݁��f�TSd�g͐F|H�t7tಟ5�ʉ�gU�ǥ�ɔ+��_|aa����bM�\e�gW
-F0,BF�A|�m�1#�Ci�1�+`N�8�-�03���w�\ьN�o�R�>"V�jw���Ru��1L����j|�V�����r�{bb�/M=]�!qʙ`��C���l�9��̙s,8��2X%�������k��.��o4;Ћ�lx�v{��4��r��z{ZEVNi�B����)ױe*�ya�B��P����_Hy�UZ;[jN (Hb0�WW�sN?T����X�rP��Ȧ��ri�B�;9���|5P���oP�98zuymA��*�59MH:<7���ӛ�#�+Sj�"�S�K&B�՛�@�``\��#\��M���[���oE�	���L���I����9����)���{�؇�i��բ�Fo�e2b�5�G��MkG�^���!� �	��Y�3�$�s����o"�j�	�A���Z#� ��Y_����/��GV�B�v~����.Ŋ�fUag��M�$�?$B� ��t�{!+�&����櫴��{�Y�����ƻ@�����{E��X��t���l)���&���修!h�#4�lsY.G��	����Ԏ���R�\ӧ��{����Kw#��P���C��B�pN��g�r�Z����(-�F���Wyu�ŕ��I�O�M���oI�� �S�!�e��(��	�>YD�c��ݔ�)���8T���������<{f�2h��Fl'�jgXeo�r����4�D��������z�:������^V��J:�x�ZOlԈS���pP�z�6��YFO٩2��V�:��61Ō����h!^�~��-��_�/��'��$V�Z0`�a��?��Q��U��KR��f
lZ>�`�^e���D����-�1B+`�4��̡ꖠj�����ΨT����#���6#��-�w+ùU�'�ߴ��)�u�ū�h�@gs�TK�6��A�3
*��߂b`�Ra�	è����.]t�$��O��P���u�s�M\=ʷ���j ���)�3�F�[m�dDgL2���n�~/��B�Ĝ��8��+!�ˀ�����	ު������F��k�H`絯��z�#��p2�mR��������dt������'�J�066%+)���]I��.�z�
X�*����U;��?����F���꺴�"/�՛�������r᎟}�Y�tvzD�X
�R���UϙhOy��L�O�[ˋ|-����\�
����i�p8:W����g*r�x�;3G��ld�#P��G�ċP��~k�L�wT���:Ŕ]	���l����@�����NxП�?��� &�1�vE���Q���K�c�hG9��$�W+򂼢�v�צ�*vtǚ���("*��|^@�	zXg�^����>����A��$Hɍ��Ax+1���=F>SN9lL�V:��t���Ň۪�z���-XV�䇐M�d^^��4Lʔ�I(F�C��3sj�r�M#���~��"o�^��7[��a�ػ0��>�����|RAm�D����go�v/*�ԗ��)������iߟmz�%�g'G/���v�L����$��}��T�ʩ�İߦL����M�R�J@��{s��}��Z��'j�gIR2^4RBᑦ��D��(fK;�tJ��?�M[�'���(�PERmZ-՛ނG��0��ڰ:�Q�a��M}}���t�`p��|L�r��d	��t�� ���(����
b����<��z�a]�,jڙ�_��[��O�  �+����O��cr���;8
_\��Ws	�\����fg�M!Q������� �m�o�~��K��x����p,����r��,�� ��U&���];��� �%�4��5@;@O��!����z���w#vר�e'��w�]�)�ǿ��,v �K��F�:������"O�<��3����w�E/��Kov���&���;ѽC�4����Ta�ҎT8f�ħ@��c�M�5��o��&���p�XTJod���p\�C���1��¦T���51�����BZ��lßE��������f�G����c���� �G���w� Ig�Z�+�R	c��H��
��_X�f.�n-���x��2z_�,+I��q2B0�u��Ď�!'��K!<v���C�� �ϹӠK�!�ְ�t��{t����-�n����c4�E��kÎ�9<L�4��+-�e� �-	�i_��W�P�p���{X����0�s�_v������� ;$'Od�2ː�����w/N��<���)�Q4��xy��؟
�0��mp���{uP��N��Y��q��H'p�V���"oM:[��4/��fڱ�qh8Iq쵁�]��/�x���x��uL~��i��#�%��4�yx�����wXi�6*
��&�D����/��Rͦ��`ز����U���Szr���V�t�$�D�j�W�ݕ�)�\Ķ X�7\]�E1�Op�d�|�ߊ����F�$�*��b�R�#�nzgA~�]�O%Q�(Q��i
��.qMhW�Ƀ�NG�ti^��T��������>>*��2ֽ�EMT�k^y��eme�]	(�-+����S��n�����|�X�7 AP�8���S9M�����&�;H�?�d{�dt�t��]Фi���>/D(w{+jGw��<E��.f��`Xr����_4�����]�ot���e���y�����g/ƻ����&q�Л*n�^�=�4'�b�@�LH���<wb�E*��H%�#\ն'I�������Y��zyC�>I,��WA�*��\�Ϻ�k���QCJ^��v�4c�j�-WtQ}�ZZ|<Ɨ�����
�LJ	��_�z`���U�J#|*XX5�`}�)���?�mm��A-��$��m~Mɫ@3��H��:g8
?~",w����1z��\�G}���,�r���(�9"P���Z���\�?si�Go`w~�a	������9�
˧9�gNÅ����ð@*}$�`��/HV�Í�Ff<��z�2#f�������1��w��ê�2-/�Xx ڪ��;�t��T�&���(�� �n��_���2�gy*�'N���Q�wL�Z�PDo�+���*�r������&�|����}�]L���o�9eL��gp8���v=*����8��H�	Báٙ��J�1�"�a�?��)̕��H��]�n���0�_�@�m/J�K�w+�ј�K{V�y��j�+a@G� c8O��=V�6	v�%-�1��fQٕ!.ı�~��_㙺���Rkn-���	'��LlF1���*@G��l��['B3� jX}�wh%Y��V3�����,���]�-�u��GOA���\ڍ|[�T�R�5�� �d�;|)�� �5���@��7�u|�C������;�E;�u�yAW,���^�t�
.�;��a���;Ay�_F]���M��q��ROM�f���������@���'�����k��?{,��(���[3�U�]"�M21�l �n�=[V(c��ܓ���\��9Q��v��pR��v?Һ�A�d���Dk��G��>�*>�X����Y�	
ׂH?[�#�yiQ�!JJR��QeƳR������+j��ND�Ԋ�"�Μ"�r��@΅��Ii'�����"Ǘ�H\���x�ȕ\�C�5����6�2�����NΤ��v���[��)���:B�H��P�шP+hE���*RaR	�E�A�����n�kn#g��KC�Ymn�T,jT��ݴ��h���Բ�t��x�G�U��m=#�jdI�>��Q�����N�Y�@�.d ����-iHQ,.���Zt�s�Ϙ��#oXs��0�ܝ�����5�Cڌm�1&'���S�އ��ӣ:���q1��N�[5j�m+ܰ���ċ=���8��}��@[c��iP[�N�=��/�<?nzrf���>�z�3hɋ8È ���ۯO�]�,��=�[�n���9P�N˥�b�I�����"�]$���{�77M^/�WyC�����6���6��.ơ9�we�p�����8�^b��1H��K���I���<�h��k���w}�WyR��sg�ȗ�&��1�����x�Z�)��)9����ET�B
�^��Z�ml)�6>O�UԈw簁�)� ��2� �'��Y�f��_ŝ/7&6<�S,��G`��QYWO��+2ؾp�-	�*|����:v{�����{[�&����C/%$)�D��t�C�y�9 ��xti3#��/i���u�n ;in N��ٯ�|Ċ
X�Q�!�z�u���,YUBf���ɽ]B�\���������b�G��̌\��q���U��T��g�0��/S��tG�g�!d����@�I�& Bߒ��,��uG-4�����<^��:��N�<��+oޚQ�o����S�e0^���\��J����mp�7Yc����>�vv��[s��$מ�d�F LN�Kc�(�?��?�dCT��=9�՘*��%4�3�Mm6.2�o�r�Tz��,Ք����b��7Skh���R ��%n�tz�&��k_�.ď�B���n)Z�Nb���*T�Z�鍥��1BO.�L��XM(�̏��хDE7�܌�u��&���$�xFh:y,�&�C?w��K����Ҹ��+�f���g<���<d�����o����O���h����H�NB}��WbE֓/��k�Z�$l�%)&�DK�:V�B�ɉͫ�9e��.�*�"�JKM�sF�$S&�T3�i�/��r3�6�#IO�\����`9��x�$_��Y �w� ��Nt����Y	��ef�8�~��I}�k�λ0H������^Au���Z���՞�ڠ�j��H����y�a����&�+�K�I��uOt��[ka^��[�Ǥ�������'�`���� ��S��h�W�0�e�Qi�eM9v�ѽ7	{�������by^z�	hY��Q|ތ�����.B"�^�l<����ќf�k�~�RHTr/�o��1�(~�"?�|D\�Qn�[xG5#�U����q�	�H�<�\�	�͐�=������3"���X��=C�<ɒ�"9�	l�|��w�����9j3�~��~�x�wҀ�eqW�
{����~�b�T��D�s]�/��j�Ր_�Q-C���╫I���<4����٣�Gˁ�W.�`Q��>N`-C\��e��X9Y�m�A������{�}3�d���J鼮��	:i��˻p�7l�w��8��p��_�̜ ��1��sL�>n�_���n[{�b�D�H���5Y�\��
�F����r-e�ʠE�BM-�� 6d�)��uM~-<��oi�ZfΡ��F	���\B*Cԭ��ح
�I�6�	jHIB&荛�mXK	]��Va���A�k���D��s�%v� �Ӆ���,��8� &ZUS��r�'wg���;���V����4�K���^�0{�~� �I�tKa++��ڥn(�N��Mu ��e��m�n�2�}e�K�P��M�byk{:6���) ���&��1������d%SG�NLi�6
e���,�(���0��ǝ1�B��7�~� �Z�7�$�~�^�P�!@G
�bx�Q��*}�-��F[� ����WS�S�T&�s�D�bH�sK&���+�e�U[&X���t4n_H�_cI�������L,���b�Jo�� {���I�<�mM9n���`��q�eȵx��<���w�gk?У��p��6�m$��'���p~VR����8�<��8N/�t }�������16 �v��ђ=�"C;�ݭ��*$A3� )k�rU%�jD��2�nN���9�ut�F�%V d�$�E���.Ue�$VVZnF��/4"�CM'!�DTY)>��T���@�r؂ͧ>���	o�W:���s�f;��u�>���	�{���X:��$�iV�2}7"�y-�B� G���zM��I&���R*�"�M�.�Q�Ig]�Hay��`Cu�q����1�����%Ǡ��'��P.�����ߣLk�j��OY&�� #D��Dnq�lJ�i6`����t�M���OV���<ϝX-]1�F^�::؅"E׬l73<tT���2�&~�0ոrĎp� �VY�(Vv�u��zMEH�j�<$#��A��ddn(4)����G�Tϓ��yʎ�]�����.,�5T�~������vϯ�o�0XVR>�IA/�[j/�l9�#E�%�8�B�i99Cﳡ�J9TL��>ٔ�}�Xա-�O������x%��w��/���ϵhJ�Bl�JI䊾V�sv�����k�YZ�NK`���Z�Q����~�{A�[�3��~}/��q�[�џ9�y��dI�ڠ'f�#�Sl��ȹj�\"�e٨��Nc �uya�ܲqA.ی�od���O���I�3zD!_rsz|z�vD�N�R=�ybs���㞉2���A�����е�'��ey��ds�iث#jĩ�?��qߞ���':A5�ߦ&j%��&ٽhz<Ne鍒l�8�Q���\��U�˭��og�#TRY���)�k꼎�$�Dc��5�m��6x�ۖ��ګ�a�N3B��[�r�R�5�#�M���[��rȁ���jǼy~2�!���~��>z�0J���wn6[Uj ��v�~H��������"� {��{���mSv:�yOS�W��0~��׿7[�;����cY���Os�_
J��"sX�мϥ(V�Kؼҁ:�*Kl���ͼ�ճo��TD�J6c��u��<E|<߹�@��まhׅ1B��aVÄnqq&��ӫۭ�ɊZ�?wj��,Ѿ
����"��Ba470�m|&O)���SS-��p��B�I-���S���5QK,��F��m�U�F�f��B�0����l�~P�1wV��o2g�Vl�o���ٕ�,���0�S�*��V�K �1}�y���Z��&�-�Z�Z��G]D�c��RB�zS����}QpR�Ȝ�`�;1��|d��`���p<���8�\6��"_�-*�8q�%�˾���C ��»��q�fY�}�de�� ����\w�W
;�X����b�s�G�X%�U�[ 5�&/���w'�Tn��B����t��3�B�ka��	�܆Ȫ�|�M��DRO(e�29��kF ʜD2U1��F�"B������n��bٺLj�޾	,�\�F�&��?&�ܥ�?LX���Vcc�
�_0dc��D@�ǝ�_��oy��Nܺx�5i:7�bn`:̷��;p~�g�z�U1�BSè�I�D�����-�G��yA��<�k�(\�>�LVʣ�qx�{�M�r����t�e�,1.�� ��o�Гgm/Qx)�!�{ ��o!�#���o�q+���7j���ΐ��mm?��7�,V!�uuq�$zo�;w�VH��!�vTU�	�d�O%���ƸI�1�o6����<�֮��X���q�{ZV�����o���&;>)��K���LR${����^�yt$�l���E;��z�(u�)0{�`f�yU����IcS�	 ��m�Fތ�����t���� �^>h�h�Ol�,ǔ?�[cd���=�؟[H�$4Z�|����	z��
d�?ڑS���L������p��הG2��7��Tff����Az�Y_v��;��x�@
ug�lB)��ⵖ(�����Qh�mgG�FMY�F�����tfq�Ƙƹs�
ђ�`Ot7���1����w}���-~!}����V�0$Ϡ+�~<��Υb�n�-�g�g׽�j<�"\��,(S�l����n;�U``9�N�	��-�c�z�����!�PO�G`�|�Jnp̾Px��|
Ǥe���9�6��!
��j���+>�i�}��+�w+����y�ۜ�-����Wg�%D~�շA���\D0*u�;�,�	�׮���ԯSH�s�zD_|P��5Q�$�9t�J�gy���%X��#p����,˭1����9Wc���~��A�g�ˌ*�R���:J���u��W��ϼ;��hX5�a*���
^h����s���G��Z��rS_�^A�B��~ b�(�r�va�����#"�����(���G�*���5�QA2*�.���ݦ��7�
���wҍ��_�N�/,=��B*���(�(�����U\00A�C�/Aة잒i�d�D�۝��K�v�G���/۶�t�5Ԏ}$th�CX��14���1�+��DTDS�����;S �?8���l����q�VtD��tWg�V-[X-Kv�>zgh��Ṁ��#mS~"Ƣ'�e�K Ե7�F�	�ar��U3K\ik(���gՠ1T���{�l�g:.$���1�&���5��Np6מ�B�ӡ1cy��/P�Z���O�mm��ŶA1���������	�;��WC�����p�i� ԇ{���õ�	裉�O�1R��H�,�H�F���'�F�.`�GE�!���d1�S���᠙V ���gbˌ���E'p!���� �/}��]vc�=ܞ؟ �A���8�ĬX�m��'~��/B��Aʹ�ҏ�J~�8�_Ut��ɉ��$PE��G�á�:c�T�@�V�XW@3c�֠�iY�z�j{ؗ���l�=�^A �8uC � ��Ʉ��~��%�?�n��^��}`��p�H�ϟ�)Z�� Lo�C�.��|]�O�5��ɱ����W W\�-Z�-G!7hy��ϼ��$�4�e-A�ͷ�3N�+W#g�q+�����cH���Gګ	��)?�'�k�5a�;�OU�&�B��>I��
�K6��F0�y����$����-�X<7�q��&ݾ�����V�^�-u�����9v��u*	/���!�6��� �N�p�ה_�S ���U���P�{���5�1n$U@�.�� s���4�a�_LMu����'��l	��6���uO�d��,�0h ����6G���=,���!|��Qǿ������ǉl*�s�ʤ�?	M���֡��h�G˅�p�,X���l�Kn�,���kQ�4n[q�sW�I�J��%r�c������
[��4�*����t����PI�70��\��M�ꊬ�灸���LI�SV�H.��� *̱���7"2r���j
��B`yZ��~����\��D�A�aUy�m��8����MP��uf����6Ρ�R����ŤQ�JO�]��)�K�ݙe,a/i�p�$�*�3��@�V�����������u'I��f�c嚕>|yr��(�V�Dn��-3t~u�����Az�x���ڣ�Ӡ�Ȏ�d� �Km7��r�SP9Nu����8�J���/l-�kM|�r�b�����]��ӫW�r$:j�9U��]������yJ_�F�)-Uvh靱g�֛�(vE�Ś	$)	KG���y�W�9�(�(�ĪX
�_�ǚ�Ƃ����u��o� 1��{J��-f�qΏ��"Es]����;ӭ��Unvv���6�|��7XCH l:�򁆴��H����#����뼠�������O�ѫU�D�9��b#* �uT"��Bo&v�g$������=\h�B���n#�,�12tJ��#!C6p�H�֣y�y��]�X����T�����k���T<�=������ �П������-�R��|�ؐ�;}P��h��̴��4H��1��Q���-J�2 =Og+q�䧨O�rc� ��p�}��D��C^Ȫ�1��K�g�aA�?�+'�`u�j}N��Js-EBғ�D��\s����+�E�������|q�����˜����u�h�����æ5��ہ}�;h���!���3�.>�d��TNY ��o'$�|yK8�}dL��H1p�{��d;C'T��b#�[i�=�EB�Z��8j��ߎw�2��Q�ъ����K��ր��S×���j��JPC�U��/�</P����A���ш�-y�R5=�?�de$$5�99��_�3��A��2|O֙>��aM�z�	�Q�����qݹ��qv�}�p|/uE�:
R�Ȳ��ח6{;��6�S������V`�[����_-`G+��|��o]�����B�nD�}�1�+�X��� �>�Ԙ�EY� ��R�?�5�Ԟ�V�g�3�Q���[�f��[��g�j]D`��!0a��r!���ּQ^���%����K�a��Q3�j��T�	=m֤�.�Y��R�"]�q�О�0+}�!��'�i/��S��LW�*z�<�7P&<&BM�°{ٖ����x��W�S�e�ad��$y�S,�Q�$��|�Aq�:ib�'���<�l�E���2��=����z�;J�*{0���jû�>��|9P	F���󷊘��p��F������t��i����o��ݟpȎb�ݡ���!�{�b ���y��m�%�B��"2���׉��K�ߥ�- ҅>��C���T��9�-.D�/KAD7�$F�<I������A�rؑʶ�F��Hu/�#���Z�l��3ef2�v��6k�\D>
阂٫���j�@L���A�Y}C
�e��$����)u�e��6��5���I:>2��'�)�������a�~9!��I��)
���?qI��j�E�m�$_O��[9ke
?eV�ˁ6�#Y�*��%�ˎ�-\m�a(C1�)r��#,f�__����B?&ƿ1_�I�tAQ�O�e`m�t�6?鯃������\�}6P���~N����(�go6���'ᕞc��-uG�����3
��X��{u;BP�mH��g��T�o�I@� �N��&�������)�aY,Z-BVLSf�'/4J���[� �g"#�l�p��鮇�|]��8�[�CBϯ?Ï�3_X�1�Z��-��9�+�\wa��^�^��%�!�ͳl��%k�cle�(vﯖHs��O3�%E�G0�:�3S�F��ճ�R'����i�m\���.��0���R[�d$+�����9A�?ѳ�?���XVf�	���9J@����2s-�ó�S2^>��&�d�5�����5Rg
X�P�]���_gZ��|�r������]�U��څ!:|LR��j�3ݾ���]2����'��U_��w�������w|��8��j&�,ɑ����װQ���Ta�zqMO�P��-�(�yd��:v2	���C