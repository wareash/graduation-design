��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���2�U�z�[B`�#�� 3�����E��R�=R��1��TH�G��N�����` �۠���<q��c}�޼Y%�(�"�sڙ�AӛXG�{|��AT��x�PL(�]������r�@�h=n�O�^����	�{K�*�q�a�T�FV���:`��Q�օ�H�m�Z<A�=p�/R�ؙ��a8E?	[��C��|_EM!���MP��� �R.Cw�j-1�,?���Mׄ��E��T��� IZ$\��h��I�d���cL�mG }������3���@T�G*C��'���"t�a�3kM�����p�s��7�Q�0�[0�yS-*e��۞�`4�,u H��{�k�p	O-O���I\��vC&�] �oV�T"f��.�=�-ԙ�v��vd��__)��#� !�z~A�]�=�[Ԓ@K�mw*�i� <���A�Si���<[V��6��C~�Sa�R�����?��d�R�^�^Nh�x'���PG)��T��ɨN*P٦W_E��żI�5��̠�����T�bJ���#�]=�3��4���׼a
I�OU�e�H����]�Wqj���+/A��|2~�wY�D�|B�SYG����8�[�+�`?��~�T����e���(l6p��kT[�9���L��G&z���w�T����[�<�K���/A%!䡢ciB:���)}`-9�T�U1^�U_�p��m�#�ba�y+�{(�9������\,n����� h�c�Y�n���:� �PG6Q�> ��a�.�M���eWd$��E�����Cr��� %�OUU��W�)�(���ڴi��Cר�z�WA�I8���QT�.K�\�� Q�<A����Ѣ��� �K�;��b�1k��Gϓ��\� Ӡ���I���3YX@�P����ߎ1�K�+Wk��^�����޲rU�mڔY&�p�|G������N81���r�^��r\�/k�F#)��g�Ȏs��g�E�CQ��]�� �(�ƙ��@�^�U���q*>Df$�m�.����Q�J�v����H��9dٱ'^�h�q*s��D���I�2�CU���|�s��\�������e������M�7� 8{ݜ<��7�z��~�a�V\ϔ ��?jM�c�����eHnW�o͉(�N��Q����Mv�X8����MUx�@U=�/r
v�ZL!�2��;��q�کK�5;��sα�'�B���s�Q��(O��0��?�]���>M�>� J�v�!78v����F��o�Q�'+9��U�P-�"GX�����`�70id�֮�"�蒧���Dm(�{"���l~���B)�@���|.�wKZ�Sm2�éF}q�	G��u=�Љep�A`�OAR߱�F�3��
L���~������y�������A�� *�*��w��2 ��\g��; ����"�T5�põ�����ɋ:4N��r���Z�)Q����ř(�F�G���؎���О� C��X��b�+P ���߭8B��ABA�/�:�5��>�R#�A_x�B�45�=~�^|q���1�@��\��ϳ����r&�����Re*b�=rݜ�����P�I�@9
[G\�&W0Q�@����J�-,��smاW���tZ�ݫā�F����GЖ��܏�(���]#��w�J����y�~��1�CV��y�7��� ��a0��ja���kݺWT���AQs�V^<e�#�<���}1�ׄ+�
г��Ƿ �n��V8hQ�l7^�)c,����7��r��������J2t�-%���mH߷�]A.9�~jD������v�?ڝ:3�^��]���Q�Pu���ܰB2��+I�h0�0!���>d9(nO�x�f 6R[�3��ܭ{;Vj����pW\<,I����w�d�����=x�Cx[tF��|� �Y'�}o�����8(4�j�IH��^� �x��˃��K�Z���g~ۘ�v/�':��k�
	���du���;ʤN�5���#�E1՚��;�(�ӈ�B�C�e���_�M�_��B�
-��Ÿ'~{<��bd����^6����r3<��E�H|H:D�}=C"����u}�������{_�u!��S�`���C�n�*�vj^Qj}X�H%[�\�mTn���އ�^�w.c������s��A\���X����?+{����ʌߢ�d�ŵ,q�s�tk�ꮻ�	�T�
�r�	�K�=!�b���W�����ӥ�k��\�U�Wگ�`����A?���*��;��{�d����� �ҥ���3
z�Z'�zb�/${�����;����ㅡ�S��K�ٟ��h\���˴����M9���.G�Z
�Q��y�\���I�i��Y�YU�Q��7��a�'^��HGO�
��Hd�ӐT-ҬS��
���a�V�gm�3�o��|�P�ͺ&(�9�S�\�'_�ey!S�%�ť�Z0�[����futN��!,P �V3�4L߹o�٤��Bf�/ȁ�iKƔ���O/������sۋ\`T�}���/cz��p�!��股�����!�{!M��ᅉ�rM 4r�wz�򇬘��kuGx@��VTFx�֚.ગG�%�D��,�9
���<�n��m��n�a���U\��YТ!��若nSZ)Y��zRd>���'��8��h'֯�Aj��� �5�@1�	�̕�U\�f:�x�5�bн�L�-�U�&���'dC�G�#SV�����d�7-��:��� ��;'�J��Zkߵ�#֩N��=��J�Ļ�yD�qGV*8[��3����}��!u�Qom��_i���Dr�,P1���IA-��;R�i�A�9uW�(��K��Zϙ���b�Th���Զ݁�QH��]wT�m>�^іT
� p���=�;�er�5���_��¢�RVi�Za�	�'��YK˭�<���w�j��{9���9���&��uOi�Km 4F�l���@��E-=Oo�bN����ϟw�n(����.b^�#��E(����F����<��JQǹ����q�`��e�R�g���ڍ��oP�����t�֟u�5 v_��3���B��WinL����v�H<�ʓB�A�X�ʨx�`27"k�D�_֫�I;����J[�Yr-}���sX.$uN��?E����u��PB�u��k�ţ�F�?��hXޑ�sLleD{���z�㺒qݩ�����_Z6���iA;ښp{8)(�'c�i���fS1v�0��ZT����y��e8jR�K����M�"�M8�cQ~�0�V��x��M���*��HVEXN#%
h��=�V,�nF�Hu;�+�\���j��w?�ψ��׈b[����_j��(���q�n���چg�F2S/M{?�D�U��'�]�:tSpJt���і�E�6�8�M� ��ʇk�+[��)G@ɹ�#'F���7�.��)��.Mi���v�	<=��"�S�k���nu�E747V�ւM���i!��#��Ͳ���}��g�7�9׽����.c՚�2�<Lo[4�IB>�Jq�y��2' �<r΃���"(�x���:�[M|y���_��
��{ZJ��7	�z�;����H�6����������ٴ��#�O0)�ڿ?��--9f����i7Fa����	_�1]c�7�EAe@T��;P|7,��'��x�}?��9y@�i�rwL�?yB?���`>��4����Ad9�Rש1�Ѕ��d��G]���LƐ�F�J�v���hx2O��Di�~�L<�d܄���"	ėE#57��m��D�M�`�V�1ğ��iGT0�!�JDnŎ;�� ��	��`-Ϸ�4:�Ӟ0�xW�WZ�\6q�9W�P|�Z��_u�9e�T���$��.U�"����~�r�j�9Ί�����b�?	`��g߲OVݛ��r�����^��	#�v9���9��5�,mgF�⦛�-�5x_5ʚs�M<�e	�(�,���Ԝ%�\�P�
%,��Scu0�]/�*A!n�7ժƽ�gM>����ݴ�U�#M:�����f��U�B8��D��4 f̱	?�v�;�Q��������9,��е�����,0���xҲ���kc��}�!e�3��j ��Z�b��{#�h��6�g�Ɩ���+��hH�ߞ��Zq�Kʂ�8�R�CX�vvq���\]�ow�Ub�w=Q�<�*q�2U��}�da,���>g��Dr��S`,{]�IzG������2�����}��D�N&V� �M���n����;͡��5�V��fI$����1I��:�YC}�3"���E�����j�R(	�C��,�%�}�@�����q�Z�L.-���1���K@����aq�
�;A/�պb�/��j�t�<M��ݝ�f~����
H��#��Q�#�K��G=��4&a�U�k{*�8�t������_	ХA��v��?�:�W _��r����w���@l{��\ f� Z�r��=�eR(i�n�%��gӏ���@�\ ��*-��p�*䄌�����%U^ĩ�7��(av�������o������'Tc�����&)`c��E�`3#�d��}Unn*q�J�˽h��rٌ�2]K�I�eR C�䴮c ��o9����k^�x��!�}�qM�~6�eZ�@z|���̛6݁6���
�x(��Z5!B9�rӟ�̮i�_��J��O���g���4ͯ`�O�&�J�2�v,N��oT��<�Y�5?��R��).l��g�NK�����Ë�.��A�F�  <.l����8MF������#�?^���D鬹ޓӳ���8�����;�n�#����!$��@�)�H�J|R����91~|�Q2�P��������x�r�ʕ�ƪ�Y�����g���v��
?L�h�[��8�*
�IW�_'�yU�_�l�n^�����if��o�8j� �Y��U2Dg�n��LXŭ���j�����7	} IO!��0 ��z�
�񨚦�$Xii�o��̣gB��޲�,r�%�����\}�0�Fs­��J���D�UL�W�i+2a(��IΔJ
��c|�D6�Fí)P���b�������Q��&��o�<G�9�	���:��F��~L�W�6K���}=e�p_貎q����AP��1�r�Ȅ������,Rz�}�3�w�T�����X���f�t|PՎ�H#�1;k�ӥ�!]�Lm��ǫ���ԍ����4p�͕j,b�ΘSP��%氊/�gl5i�R���F�+��g}B$;J����~��8���C�}�0�9�❰��e�|i���y��B�z�҄U1�'Q˓�� +���ڋõ����o&�"�q��Β��Km)�g�o��IOx��:�]9�k���"�(���ǵ��v�K�l16s=����^@QS|��Ɣ�E���6��4QS���M��'Dƥ��u#d��龵���~#��4�3��iT���q����I2Z��K��9&�jn��ZI)<5���pK�;�����w�#J��/��s<�镁 ^��!a��(}����߇�G�n��l��E�McFN�tKh��68�Cbx�>��)I��x���mXuzZ�>�%Yd�('�����`�f�8�+������$J��f�l>\h0�~CWL~�}�t�G��*b�f�덽uTOh��F"��5.�NXS��vk��Ω.2��Wn��ZZ0)���v���u�bU=��q���r���u��F���C�<��?^�V���
�{ �V3�W��ln���E��F>�d����!���{XP!%҆ӹ-��?�2	��
�c�� �.�/:we�@`���G�� ���Z�=�t�<~k���P�'}'s.qƞ�&�D��=���s�ɚ5$��1���d�D~9�ۓ=}��vq(���q�'�_�4cu���$�����S�Y#�	a��t
-,��k�vR��������:�Mx��� �%���V�)�v�:�a�>�:ժ��dg﬑ؤ�#�.Ƌ�+��w#;H�(�(��y��]"䇺"�t ����b$�k �!:�C�u8�z�B����E)[^7��{I��\/�Q_1ڗgIr�1��`�N�/�2F��%彁�r�.
ǣ�M��v�T�)��=�B�t|^�܀4m翵����g�z�������kݗ���5U(e�˒��:���-.����� ���I?����?LJ0O�q� ��O��d"o��1�E^U-QD�uq��c5������z��Y�e�͐�Y�¬����w,�sj����3=�zV�ew�?�D�2I��36s��#����5rG����L�o"����0��B�Qg�&���ʉz�:|8����Ĩ�j����}h���OqdϣVͳi$��2Z8�=�?����U[}k�RS��8�f���o��!�9ȩ��?���4�#���dQ��
�d�hsb��8�p���;��cN��\�fZ�����(岿M
R39���P��57 f��}��
S�m�.�(�Wܕ�9��Z�3<5�.⻔�(�lʻV?+��)6�;���ݫ܇k�X)z|�F,&ed���&�5�hqqH�}�	� p$Mձy��e�z�%�gZ�	nx��[��r�YqxO��ϒ$���3�����/C����
:h���>Ggn���I	����#�R�V����|���3�dm��X�b�hx��
����uL�r9�+���.�gg�JP1�pݞ`I� ��9��w;0Գq�*��á,d�T���^���D: ƈ��Rv��a�~��';I�����=ྤ�.\Ď[���K\�#z�����y-~��4 &�ƪ��΋�\�-yR��!��}�%ۏ(Pd�2��'�$Hp�5?�/�l:~uOrg��й|�!�� ���=F�e��槥��ba����+TØԿ�غ�d�~�P��ϒp�\8c��ߏ��%2��n�$�i�0�ί=�K�J M�R�x8�bj�2�]1[VW��l�Յ�&�T���Zz��|M)^�]������$�O�r�r5��_%]�+�a4�%q��_�"�p	ʹ�����ZH��x�$�!0�B��zm>BVD�V�����^�"��Ӱ��쪻Si@dD7"�a���0������y�9��|������o���z�a�Զ�^�ݏy%p��y���ˈ��!�06��bKw���	4e,'\Q�*�W��ta���HLC����8;T��B`ʚH)k����ͥ�!:���=c�)'����� .A?j�>����o��F��Յꔼ��������n���+�����T�nEw�{���@{T{H�Y�����Y�u��Rqd��u[R,iq�m'�x�e���'��)�����ϸ��D[��n��D��z����/���"�˂��:_"�_�q<a&W��	W=h��������}���OUb�#���#�WRA�]�-W�?^J\�3V��>�5W�yr�i��� ]�lw��4�,�{B�.Zd�Ό�c�����m@���qD(	<KC�`���d~�C��ܺ]��)���z��ꂌ��0�֪h�(�
�ʱ�<v�_|�!%��H�2���2��J�	�	��Z�>����"��L}�ew�S4��1j_���0dۓ�j�O��[��
{O� ���s��(^q���EuP#�Vc�_�N)�(%�u{G�S��3�RU�Q�����7��{8��o�$�uz�9�2�5�Pu���i�c.���	��2��	e_3I�6�C(�ߑ�VU���|��w\,v#��C�/T���K�L}8<��R ��G;��s�Uv&P6�a|(}�]Q�,�ɶ�-�����s?�o�,׾��m��zAh��8}�g�FB���"]Qr���m��$�B������ ^H�����Q(�eB���?'0[����%�QG4%�Fy�� ��pI%��#t��%��ߪ�5���\�D%&��`��v��OBlS��N��&�19�2����.o�6lϐ��,u���ғH�ٵ�w��?���@<s�� �݋�KP�) 7����U�k�ñ�l*�{�Acr�qBF����z�ك-�B��Bj�U��*����S:Z��yC�����H�����ym�,,��p�|��nM�Z�M*]��,Ǳ�aI�48{SQ��T�J@i���]6�6Y����4�E��V����0����h���O�z�n���n��j�(�)�Y���t4��d�'�@'��,��O�����HyWN'����	dI9�]�tL��W}~P�9���?Bn�W�m"4��;����.�_6��A��i�/�2e������:����Z�J�cn���/X׫��i.��
�ܩ+��𾃶{Mu�
N���V��U�x���)M����"�ba�7��v��D�[׭4�#&�&�������S)�e��q~gV(B{����T�)$�|� <�4ᾚV^���$�v�,�߱"�򖻆J	I_O���~&�RU��7͖>�y��aF�m?ns�L8�<5�K8�Ƨ�X��SW���0�o�����ٯ��kz�LMnE�ҕ� [��\�Ȧ�~[o|�jK4j��F�L�=�,����@�~x��M�up1�c~s��YL��󔓧�'��Mz��g. 0��[NU����a4y��&����33��(�0o<"�z�c�������/S�b��pU���i!�y���d6!��`C�؍[u̕�K�ï\a�7jAg�[��F$��e��&_�n����\�i����!�=V}Y
��޴9T�Y�w�b�PP��� ߵ�D��)W0�,٫	#߿��5BK�``T�XwΎw�Iz"�����"���g[߄���3��2K�s;X�xA�[elJ��$�Xs�ڶ��tU��5��r�b�J*:��A�L��.�h���T��b#��JhA��JqVԅF ����O8��/�T)C��G�.a����O��/ζ�U��� �g�52�����UE�������@����Q-ƙ�oL�^-2-y\l�KBO�V�W��)�X��������:7������:\�<�bP���"��	|�s?�~�=�c%Ohیpd$�S��4G�O�µ������,ѡ����J�5 ۣ�X���'Sa�J�>0̃���s���ɵ���18Ϙ�y�ͽ�&{�p+�1	X<����.-\e�Vr���j�v��pZ/oއB�+�����B��Ƀ�~:D%�ā���62� ��=˒������6��0K@�0te^�������O�=�/Q :-Kg�^<��������%r����2!褳f�T���V񗞢 �]�]*s"i���)�HM�<��>�E��p���sXl�i�N�4Y(W���y"�ta�$�n�)'�bL�?�bQ�
C���V{b��h$�UŵӠ�pp���K��iɻw�X�y��31�.Nv������8�M�Ŏ�%�`����0����E�lB��p���֞B�9Ű�ܕ�Ty��TX<�� ��,@�o1�q��hI��৶�W2]ٗG���m'D�gXY�p�Fb�MD���76D伻�F���^{�
�j���{H��+1���ȴnw��G}��O���8Y7L��q&ֵ�&^�e��N�u�i}ʑ0!��B� ��H�N�#����,��?E�J�L�	e�4�|
��M�	2=Vn�΅�wR;cL���kw3�[�[ � ��
3� �<	��m<���nԽ�Dm4e���4R�S��f� �'�F�����oV��zMw��4-V��ITj� �%
7��ܛ>�=�܈]�Z�k��A^Y�&'��.��
��uD�q�U�%��s-���<�2ƚ ��c�D�K|�YyB
������!±v����C��绂3��O�pf���;�/����,�L	�a��P��4t���0�E��B��!\^��;�k怯=�6�����^]���
� �����& c������3��5���3�<��L�x�>A}.�7����o���y���h������ 1���?Շ >Hqu�YՉpa�K݂�L���{:��x�`ICdz-��>�/�m��re�����'�*_��\�:&��+"�z�*�������(�7[R��,�h�i�E�@f�ƻ��OMiI^oN��.��F�|R�E��+��_�Eܟgq_ZH|;�]2CS���A����'χ%�`�O�_�_�<��P��Dņ���P�><甏�Q�ښ�/��uM
�
���䮗���s�G:�Y1�B)��'�Ȕ��.���d�R�jKf����X��]HLױ��!.�p8����y�Y�tJ�̞�	u�"0���)9VP`�MB�>f_�
��?�� �@��ȝHQK�Y�I� �m��A�D�������Y.y]ʠ����W���k�V����k��y_c� �C��!`P�*�H_���5F~x
�q�u�\����L�g:����np�E�����(����/A��`b�cv��iy�#��&NN8a#�18 �A��V?.��t~ߛۛ\�I�ѐ�,�e��@m�;��+-����S��k���'�)�Dh�Sl��>�-����N"���v�]�NQ ˳�1pܓ�q�:��TN�O�(~�x| ���;�б�xY���KL���a�z�i�7���͞��<�,�]�|�/�d�����|��8p�����e��C 9W�qx�b�#���%�ZJ�?y�?��&��j�c����@e�ě������g���'0�e�> �����K$`�[
#Z�d��95�z�L��|�iZ�-�9�`��Wp[RlzA5r���٫�:��=�ef��:���j���8ؓ��W�����̾�ґON�p��1�}B,j)>�����Z��Vi��_6R@�'�d���өo�5��	ۚ��q1�M�NX�0��t ���� s�[�9u�����B|��ղ�q�2��rnZ�VUJA"G�T�Ks���Y,�+���J�d��E��"&j�J���e��4����z�����`m�V�_,��{�칋`��A�0��gw]|����E����ez� %OV�-q<~���>8F���_H
�ވ�輖e�i��j�y3;L_���Ն؅�w~�����n���;n�fV�^0H6��ַ�Ь�ommJn�������*��r�RQHnx
I��h?�β|�}�	P�}�qh;�R,a�Z�S�ӎ'�	�[ ѥ�:��e.��?qh�;
����"��*�me�
��%�a��f�L��-�gv��9Fd�Q�-���X]����e6�сNǷ�|�:*����9
��d��<�X��W7����F_�~���	.%g�rW���4���#�@/52�1�����F����f�3�� ���d�@�A��v�/�}�.��:%�d0��|8`�f�Ճ9ϡ� ��ʺl�&'��6����k�l��*�Llۤt��^�.Nn|(��,�|����#r���!#�p�|<W�,��i?k���$ź���4î.	x�X*���C�K��+�^�����u��!����x���Z�/#��X-3r��EA�%��%(쯈�?Ē�`72�����336$L�}�s>������` h����(W#]{�
��3�&J!޷z��iZh����|���,@�)P9F�D��` Pӎ՚-f8.T3��Bo5��}r�.I'�TVqC���[�y�#t%2Tv����t��)��	�NW"&|���KڔN{���D�H�~�2��
�c������3h,�=zL빞Z_�qK �	I���OM���F��9ַe@�9j<��n5>n�Z�r�œ��f���.������.�yS�5a�c�(ϖ���?���P`ma�G�j��1��
2�`D.k.�6�7�Vuf��ũ3��7�};f��}���#0k���S̷��.��`8-�h|]���#�j�2G΄B�~9o�C���V8\Ԡ��]?s�<#�mO�'���;��6�������vn�{���7�S�>�`a;~����Mx�'+�IZ�}Pk�>��FN/e�-�j�QE�֗�#�i`y�1����9\�
s��BZOe�~m�uC�A�Ӏ��j����xq��A`i�Q��MS�rŬC����0�[�f����0�@�{��s����Ha�(H�s��FQ��	bg�b���A�B����0�^���_�	����z�qHx-�S�.��,�@��� �V'p�C�eN$���G�;�)g��	H��>ư�D�(lV.��C	�V��X����b���Z=lGu7���v0]��#�Y�\"�'en^�<���@K7Fpy��r�:b�i�Is|��^9�摢�I!���7��У�����K@���Ne�pz��bF9�Zk ��đK��W7	��,������V���`_�!�����.@����&0&Jꍴ"�"j�
��S��w�Fo9���+5�*c���v=G��Z�)@j�Or]�������*L���cM�:�ٜ���D3ω�6c4��^l(����B(����޳W�)���X�k����p\�Z��xq���2�i�#�6��~[��%j�q}uP��:��C<1�Q�D�s����C��u����2ҝ��R*8z��x��}[[��n�fZp�x�v^w4N\<L��z0
��{y�L=d	��1�/�Wv|�0t������J)�!iߑO��;���ݷN����C��ĳt�w|��f�y����
G���u�Y1�#�GR�]��Ξ3K�|�= ��R�{�o��zTv��p2[�0�-������ļ�=~�і%Ҡ_V�x	���l��r�^5^�J�M�;g��	jI�f�n�e;������zS�E#���"e�
��.�:�7:�U��'<m����5& !��)?)FFR�h�-�bhG	������B؎]h����u��5���F��6p����x.�`�@?p��w�D`��M�]R!H��P^;��C-��2hJ+U���~��S��Ix������X����emTS����tܖ�C��0�Ƶa~k�������1+^�\q�x�33�#N�ٷi�y)�Q03�|+p��8hGSJ�d�)Dv34�������^�������Q�a
��פ8�F{��L��3^X���?QM~���&�+'9=�߱�1���)�L˗�ؒE�3s>�Cw8#ʫ�^�<� i����ϥ���R]Yp�3����\�Z	�2J�`�I��%�bz�;�!ef!��c��_��Dߡ}Jh�Q�ԧج�W◛г�l�u˻������Fklۀ6^5Z���m�&�J>�"b-����G�Ǚl]��u���d�0er�~F"��֯���G�+P��|�>ʂZ��i|�_�N_��.�RiU�Z#�[����jz1P1N��3Gb��ek0�'>��� �m���
�|⃳!��0K��ɴ�p����3��@"b�	 ��5G[;Y��L�`'�L^���7id��n�	�P��רs/^�Шc����4=�bc@��i�bȠ"kO��h��B��wd�tZt����1T6P�y���7b��KI��_ ������(Y~��"@�s���S�w��̄��A���p���qf�E5�U@������P�._܁����Z(o�!�|	�ܟ�����^���2��5w�;�%{u��|�� 
�w�;���nEGP
XH7�H��*����3�"{�m�2(`� f���9~���n���8���O=E�N�:�\�����J9?���uM�ï�������͘hC��D�/nC�0�U8>��0�j���(@�CM�IR;f2;贠��/�Mh�Zl�r	a��JLwG�P,,�S
�i�a(!�zp�wm+���!���y�}�H��ޕ���V����oo{篽�OZP<�ͻ����>��C�r�h'��9k�(g�D�f��&��O@o�A��E@Lh�x}4��$z��pͳf�&c�&M˹W�v�L��	��7di���v�~
ú�5�����48ʡk~�Jm�T�6���6�<:|�%?���*g궺�	������wD�
���"�K)����j\��>���1�&^�za�zkE�0.h7Y���I������/R+4x��B4g[�����ά��ŉ%�~��^KO�⒯�2��P��'��ѷ������^�M '���/o-����}n�F��B���k֫k�M��������Z}(��	�t�!"m��&�U�1�t��J> K%���:��^ن$Q��L����5 �ePJ���w���k�� ��o�=��,�F��/��*Q͸�<Zi���@��,�����;�4)��E�b�iSr���AG�'�a�׭����J�sG�KOv� t��&x�&�}��<�n�Ϛ��T>Jf�<Q��Dj�]�Ut�d;�To��A�����Pɍ�5��e�:"
�g��۸M1�@M�ƶ.�QI����n��v��jMZ��/Qk4�����-�:���~b��:|B����IM4�%4�ɡD�!-�`�J켕S�З:��1�}��k&��ҿ	�)!���m~aZs�bKY�<e*�IR�&!�t���2�����4�����c.�տ�(�N�f�,z
���<�[���B�Y���!5�=I �	I��>X�6��+�[0>˞N��F?*����"l�B��u���Cs͜�?������(��υ�)�̎U����>tv���d}oR��g���"�����*�i8$����v ��
�'��K�]x�N03��t׶�)���Ч³�	Q��f��S3�1{�	?��&�Gd�����W���ě�|���8��ۤ�DG�{<�N�l�َW9+=s��O�2F�^���*p�:<�{�����]���#� ���-�.�:��F������~�ܱ���M�G�`�F�Q%�P�:�Ճ�a_p���ތhF����u�B]ի^�0uu�(�j���r�ct�GQY�o�F7�?nOX��׾ol��)�4�95�;ﵻ��� ��%;+7iD�wP�����'�0��l�P�Gy%���}�6�H3zb��R�!� 2�*Ď[��������!���d��H�ki� 1�8�tT����[�R��G�T_Q�� �׎̱̓l����l64��r�
E�Nu�,��2�*�nc�XJ��Եa�������?���6̂����&������ʒ����ÿ�X�L2�,�< ��=~>��r]����J8ӼՊ�=�⾨����s�Ƚ���=�:Ԁ�tL�v-���L���I(�/X�b�C@u�R��-D̄��\�m��ꤙC�*)��6g�^T�#�<:��6՜��U5�� �/����J��ƶD3J.J���È����͞���j��3�I���f|7E2������?�b��%��u���aP�F{~55�)J�-/7��1�1���_���;fv#�?ikck�����R�r���{���W�9�|Y�i�WA����q�SH��\���r��q��E�~�[�0�c=b��K�ɍ���R[�=�id5�?�[BSv�/��W�x���L�����#��V�L�#�죥S
���2�d��u���֫�Y�~	�g�e�OR��/Y��5z&-��H����w{���G=7rlt���`r{�3:^kNf��Nj3k���y֬��8d/	>��w�nHv���-Kq��]�Ƈ����C7��_U�\���{�}�aĤwN��̸z�sC<���0:h��� ���'~�g��$Lu�e|��5�Z��Dь�6�>��,��-��i^���#D���<57M�1mUZ��d1�i��I Tꄱ&?\��ui�i�ܻ/�=<����>��,��,��z:"���,�{�8I��k��B�p�acwlW����A)j�oQ}O�-����(eu���m�r��#]l �Hq��CO5C�� ��g�_k����,�g����T���B�w��v��.���ko{�,zh���v&#=	Iya�+�?y��h/�iQ�;}�T�-��D�Q"����P��S�Y��J�X����(�yb��悍.������P����M��;���xΝYK�۟4U�y�V���ϲ4]��]ém_�M��eL,&��G�����)fS%)���1�����+C�D�}`������Y�@])��}L�  �{��yn)��\ݻb5~6��f��63�4�WJ�8ߔ�,c0$?ml�X ���<g�1zy�W.�AQ�x�0�s0� ��"'@�;�p4�R�����^:R��ߎP�K��F�UU '4uD�ֽT�Lv'�jGQ��zϡ�C�ܑ4ۡJ��+Rq�"��-j��)�����&n�~n-VD��jq�K%(	�m�E��( �=*����r��Z ��#7͉E�FAz(ɤ���s��v���$�L��%FK��)��c/����D�����V��L:5=�(�ǖw��׼L��?/<�E�a'���-�
��7V:l��r\>{[�b�T�uXa�p���|pgA[ax�~JN�;�X�[D�T)��ef�P���T(z��?�6�a�I���Ă�c�D�*$E4V������y�����ЫJ@lT��Q���� �Y�Ჱ���ѷBL�ڹ#�o	]��LK�o<�'�z����y6n!��>)�~���玟��D�%?��O�GO��`�x�LTl���gst& [�M���c�8�!��P�|2
�W���Z�!3����5Z��[�c�os1zcC�����_�R������F�FK�*ǃt�֊���g>IS�Bo[3��W�џ�(D���|���xJBF>�� Q�
Y{%��-���d���<���f���]�s�P�� ��8(T�%��7A��ì���A�~/�w�� �s:�R�`Bx��Á�+ %��I�4m�U��h�����jVOHD@R��F5V������|'���Q�۰t�X�K!G��ya�w�n�@�0/M{��6t�o�`^ ��}W23��m�)bv�I0��+V��/���5Ww'6�P�o�;�|��;V����g�Bb���U�����*1��g�M��-��^Δd��p��	#TS�EA.m���,��jJ����j`_)tSUn�8��y6/������~$��|,�aA@�}aM��5�\��z��PA�}c����?�ћ�S8ݧ��pB0���Z�(�䐯ځ�T9��;�ArΗs(źR����e{2����hل�e"���L0
�:&e���(�$6��s����7��~����r>�w�-�+��I �#���v�n�K���S��i�|Ϩj<���p�;҄�}]	R��a�ks|ThƁ�@�T�BH3��\j���7duFSH{3��n^7S�����;HQ'�x̱��O`ʔT���+w�{W22���m�'ۗ��*�~.l&�M��6:�4=����X6@�����{�}o������켦��o�С˛/�����&�s-�/���gDhV�(% J�Տo�� ����n��U��/#�����lJ@8�4���}�1RIN$b��� �͡��ڰ��9�WṄ2�c~	V���.�u�6�E�����yG��؋��Sk�]��s�F�0S�(�倍ւVLƾ|�������ЈD�&@���/�˼9F\>,d�+h��'�H�f�M��F ������6	\�@�ο�c}��>ϑvog��Ș���N�7YQF�\m!��dw�0�ِ�� �Q�B��/�?��)��\��߈�H�+��+���jWqIH/�J�p�r@�Q���J�c�����������m�jI�[-ߎ�[�|�����n�7��8I�2�5��E�9���.�a�PRr�F�}s�����j�o���H��'a<R�q4�@R�P���\��hcٮ�"��^р�;"=���9�l�^S��5�Sw��qvMo<�'���`F���{jl��k�(��Cp��r?.�>��oD�"�a����+/U�C�\��V#�ٗD̗o��H
����h�ˮ z8��[�3myAs7�ٶ��U��؆x]����!`!Hg�Z��sBU��ɋ���Z�r�E:?%($g�^������,��?����f�'�	�i0�PΈt��� v�h�2��Du�qbM!��:�A	�A��8p��_�YǼ�b`��5�p��^a�m��#@m.}q闛�O ��q���k�8F>�Ps|�� @�
H���[o��n3aO{ o�`%�耐@�����N��MvQ	Bi�3�PTa��~��v������O�ƻX�`�<���	���$�c��p�~��0LVRb��+ۯ�׶Ռ��Q� �9���.�N�͕��g0�qWu�RћL-Ä�4��D���R����?M:���j�R)���)�ӐͿ��x�3	��J��S�(\�H$v���"޶(�K=���/{A����/�C��D5�8�!(EH�r��G�&�������he���4���z_�����3Ž�J����?L㐨}"'��p&Mw�D݁&!�7�-#�Li�`'Bf$E�)��D����SMk�w��G#��2��yHfQ*��������~fO>��k��5�E9>$�d�Y��~�|��D���ֈЪ�^f	�tc�Y�����äb� �5:�]ڄ:�uM�(R͞ú���b�B��/+��Q�	 �����%S/)���de��a
�"(@` >�hH�ɡG�.����!b�I��c���wT�$�9Ka`ŕ$� �u��bU��*]�	��R�G����`L|�&!�nY(>�6�N�=5݃Ѥƫ�f�n7��+��,1�$��X�H����'�����	�{��~�A�hYX��?�޽e>ɛ:X�18ZY� �ԯ�q��	�oɢ B����f�?��ĭr�9�H#�E�]��ԉoAV�[O(�)m-bQ*q����C^x��D�~�Ʊ���L�nڪ�τ=G�ς�S_�LX(�"a��&]t��b�ɩ�i��50����j0��Y��1�9�0=G\�ӝ7�D2����h-=I)�-u>���A�+h���E-c�jsz`��D,p�!�s���%�eUlw[n���jLĕ6�����ǟ��ɇC�|혯�&��5�K}�af{S)�X�vEW�,w�֬�j
�,{�GqHS��A�P������ĕ�Gb�¢�*��T���ä�����d�A�[��3����l�=l�h�<4KY@G��'����ڌ�d���I?+����L9�#�D�vf�������XCd����g��sB'P2�5&���6�0�We�s�v���J��a�����8Z�Om��cՂ�o��;����&��I����U�s�I�ZT�@ �6լ�vFv����v{]MEd�i^�F�N�	��X<����>W��ҵK�s#�������("6��'�JQi�bT]�ꤵc���*c�e���@62,��������Y�����z ډ�(�(0c�Q$r�}u慒��HU��yqt�� ���Q���v���*)���4��%􏠜�2���I�����O�ބ�Z�1�{� �ё������_	�^�(����r�SO!'u�Ё��~�0�+Q(q u'�*m�$���\��C���q����=O]�qHB]�"�w��?Ge��E�}m~������j��&��̃�O�
�����C���Q�2 ��'�_NT8�}��V	M\x �n��rB����Y���xGT �7�Ȕ�{텝ߊfi�b��Vwڱ.׶�̑��[%8$?�7�,��nz�#%����\���WA����CbOٴ��|��^�5� A0�XbH��v�s��I>�{����OF��6�h`��:K�z;�[��A��]tL�Z�����o�=0p�忻�6ob�iB�)��I�!���g(__�G�����Q���$�F؊dL*gy�G��C��j��,<G�Uل��!���6�VL��ac�u|���Ji�)l�6��W�k�AbT-���̹������sRZ�{)3;~�ϧa[����k�R�-�=���B�_�r�p�+�0�xu�+٘����CՒP��m<*���I�����$M�C6��u��0;2�1"p�4�᛺��#�8�{A��&�ɰ��T6��B:�@G�ow'!��� ��̥�mS��`
V�*�P���\��\h9� F5��IE;os v?;%�Okة�k}�����N�GU�����Y �Ĥ;���d ��l��QN��M�lM�����o�3[���p��z��[���yB�黳��)$#b���!��3Nz�s4U��ha��m�:봬�� �P�i��q�C�ē�碻]c�����d��ځ��h�3�*'^	���[���Kc-m�'޿�=��|3�O�l%q/k��� H0ȹ<�h|tk�\�C����#������[�Hg�X�2��Ɂ,�\�0'���>���_��H	��▩��{�z�ƒo��1|�2B�Rz;�Dz��(��@Smx�JbU&
�O=��u�NN�C{�{���Q(�ȵA��V5+ˌ���W�@`�}�v4�f�����
o��8Mfѕɖ[������2G0�>tӐ��ۂNt[$X���zG������{���1p��qI��;-u��#ל��(��@,+ޟ3>OB0��t��%�q�Ҩ�d���|Km?aYA�o���?Wp܀��~�Y��"F�����U��,Q&�]p�,s�����#�,��o"�I}�IQԃl��s�k�W�����@�x�3��AZ�!��GO(X�(@�W�܋,�bQY-�D:B��:�ܢ�g/.���i̎������<*�ǚ��z@?���U��C I��HZ�d	�I}�����vi
��S|�<HE֕W�m>M�3<n�Sf��i��`E����}�o�b��v��H����/��}���幁.K8��c���O88�u��5���M�e��!�Bm�ƚ�dz׎�1�ꆶJ�/�����.�l�|��wK�qf�c�ve��߷�u��S�r��;dc��zbX=j��&+���l��f"���*�sk�i!�,�{�g	,`
���2�;�$�BjH���D{�d��x�R� ����y2H	�X�9R$|l�	 &Sr%�=�(����S��q#��Bz�{G���_�*Up΃���`�b#��Z�����_׍��e�D���O x��M�#��N�˜'��y�$wuyL
�	�Q�,�w@0L��.��;��|>b9y��������tnk�f&>��[u4�`3�@e,6b �˜c���9)���T�ϳ��w��L�5YqY'�!��*3R��2X�s�;$~�3>�ў���-l�P�ն��sW��cƱ��zO����Sn$9noi4�=̶�F��:�x�;U^dp#�И��4�5�+[���ϯN1Niƌ�P<ۥ;6�w�:�$�a8�$s���\��z�گ��l.գ�x/;�ɸc����^��9��69$OӃ�#2�@�D�۴h.
�5�[��Y���9.����3Qed��7��N$�.k��w���DjTc> �:t�2���o��"����Eb�	\
ZM�@�C'�(b[_�BMFHN���De%�*K /�����߇��o���g�,]�I�V�${�z;_�m�O�L�Lj���.˸��9�0,�Y�O�ȣ]�+�ޮt@��I�9Sf؈�O�h�K߳9 �����¤/���˝���s5oO@�ն|�%��q@�R�
�r����,!d�W�rc����[���g-���2@��$@�+��o��!j����ߥ�Ҁ'eR'glC?��3
�������Ph��	)U�	�w�E��F�ڹ���x�#�g�=�N������԰�qՙ��.{� 3h��3���xGV��4U��3��-�ڻ1X��l?���:lH�bO>�yI?�38}������A�OC:���b*��p@�z�op�9!�y�,�y�(�L!^���5xA]� �c�:�9C�q��z�;8w�����9�1)&p�_�\�1	(�!��H��~�z�*�?���E����s�&x��u�[I2�|E 6X��3�PpOt�>w� ��m���۩Z��֥
��<#�����ܫ�_kҲ�u{��ݣw!,C�K+�r���I���1�S��`L��ɈZ��1��bCf%��y�T�gj_��B�r�aɵ����K�����k���:rN���tؽ!#�U�tU;�c�,�����ݨ�X�:���i��_+�_�C����14����#p}�.�
*�H��{QJ���x!32VP	5_���|�m��-;Ъ5h胠�D�;�W�>'ׂ��i<��{�	Q�̽	p�٫t;²X�UI�T�^�ŧ�&�֕[^���{���79N�v�!ɴ8�8d,��j�0?]J�q�v�����Nm��^K%�u<�������yr<����F���K�D'��<i���b3�qm
�B0��-�S��&�O��{���������h.Ї�>���~鉷��e�8l���y�,/w�"���y���{R3�H>�X|US�>x�n���`*��~~3`�\B��1b:��1n�7]�`.RxR���/�f=�PԧǳOI��%7'6(K�e��=9Y��'��a�[1� [z��)��b�߽j��$����%�=D���y�9�,�y�Uv�/9̚s�aC
%��ƴ?ӂz�omo�	.���&p�n��2�����p���y��C��R�"�I�B���	݅��me��dCI��n��_Z)=r�=�y���%Y2��i6#.�2��J����J%��w��{�?.;ޝ�V9��Œ�'K�<Y��n|�ɟAQ�a8&�����|����Gd��́�b�3�/K|t����[�O���y�3j�&�Z �]_��X������	�����nh��
�]�(1װ�sRe:�Ͷ�<��J�Y��������{<�c�.~��@���3�7�g^=<T\����F�/&r:�S86Ҁ�t�k�ʅ�N��v�h9鍍�~S�A�,VO��d�Ӱ�ih���lG�$6�����Z~��mS�ߑʬUʶ�|�#�;�X���BH���g��^�0o��
�����	��bpb8��c�ّ� 8@4��<?���C���� � ����Z����Hs���.
��>U�EED6���+�H4KxG�EMb��XE�������A�]H�u8kc�)�w��V�����qz�������� ѻ���+�c"��i�7dg�V@�1��k�d��p0$�\��W:��%[<hW�tGYv��l�,
W�@M[g�2��Y�r��[��O�E�)���N��1����{2$�Ӽ�h���L��ٰOp{���k*�-Ҵ�A���o�M&��z�J�ѐ�NN���A�O(u��ME�����n6�P�4�3\k�X!�uq���v�l2��&��0#��X�ϗ�v�q��|qW���+,��K"�S���"��
]�\���|g���C�G��ߑ|���w��;���2��wWRC��6@�q�����։�.=FΩ����Sa�Ue�z»�P!�X7�w�C���L_��xK:�>�	T�
�U���d��KR"�.k���J\����۩C4#�sO� Y��pA)�/�[U�>Λ�������Ed����\@6&W<'�=M�5�ai�c��cZg4���
�7�58 ����AN��/;,��gr*�� V��3s|-�q�#��ɴ ��Ad��}3�Z���<�@}�����GKx"�&��Ħ�g�� a�SxǹP�^�A�����
U�yX�U��ɋ���[�k����lUïj�C�CtYuQu\�'��� �D�B�ވz�$��r�#,��� ڦ�$���v}�����T ����KN>Id�^��:�e !i�q��z��!S�O������:w���n�\�� ���!����n��4�殣�P˔"�/m��-`{N��C��)Yaq��	s$��.�<���p�WH���֘��È��rJ"�8�����?�k!z\Qq��8�[��̾�:q���;x���@ᘭl�*N����>��}��`P�խQ�&�S�TN�͖�_�i.�T(ZV}һF�`��N��H������& l�Mc���7���������4��!1F �B�]��d?����t�ܦ�h�l�Ԥy�*8Ou<�`����4����v���D��a�	,hj�xy	R&}��Tl�A�)�M��b�h9<<��ua���!�1r����r��RՇ�\��L���1I�ö�ɥ���v��]���˷�y��ܠ��K��,s�JR�l�
nj��{��V�N�~8{���N�k�╩G*ga����{ɇ
N��w%#D-����xU1ys�_ʶ�ʢ4pe�6������I0���
�s�UQ�ӥǃ5�
�\:�y�=��^����������Axe.��B+�Dw�|�m�7$��֏���[�F�B����PM	��ġ����\y�!8���s��8ʜ˪^�]oWzU�OҰi�M�Չ� M��Ц�W@��+_�!N�Y��|u9�����`�c
��CU��#���ڵ`���$b��i�K��n����1��U�w���szs<��^�L����,*�&)���]����H�|�;�3>�?.�7�𝴈 c1�����Q������E�O��鰤����C6�H~I����Ե�eĦh�h�s0]�y=+�@�L��	�ё7G^z�������qp�.�!D��	��bovp$�ׁPk�2��x�kR?LY�o:8�Y�g��nOa+��L�Gzn�d�h�=����yc�����b����7������:��v������gx��k��N2�贺���os�*���Mk�s��n�~0_8���Ζ�`k��������z�q/IlN����߆I�UX���ܦ�4���1>�|M@�r)���M�ZD
�$��>bF��y��V퓒��'�گ�Tw��)����1�} � ��x�ύg�{����=���Z
!1l�O���KI|�@hC��+>Bh*�Y��uW�Ăp�B�߄��#����|p���|v�!�0WΓv�?U�bk�j4:��1'��3R�G���>�߿A�l������Zo���E5�B\8 l~�9�Oc7��I��㐚(,�Y�N��4��[?t�0Hm@C���ø�xQȁYaM#G`�v/V�{��npw��c�����G{�i�ĺ�xз����AJ��uk�e�,9�B�����wז��fV�^
 h}=�A@�~�0A'��)��Y�ܚ=��/�(����R�N�:��X(0_))MS��"nW۰bv
k�>�9uc�z��C"A����z��~{B.�n��c��$���Я�5���;����+;|t���+����cZN.f1��:a�����@�"b�*�,�/e�O�U�wW�m�{`"�~�98��	t��C3ǚ�xR/A�	6b}!��M��=����a�v�쒏��{�
��ǡ?z0�����g��lY|��E{ԡLo��6�5.�Y�p���̝�<W��K�R\`���	�V9f���SL�� 8���O����c����"���М��ħV�|j�M�L�Ql]Tz�����>�qH&��K�}���k���H#�,�C��}�yK֋����)���`��c�\p�n�4��pp�쌠����-�������4џ�P��wt�*i#=�& $�gX{�T�zRW��GlG��Ψ������|vr-c{Z��6���+!�o���k5S�k
�jzZ��%�Lz�s�V��3d���(�\BI�R���rZ/6�lalP���I�F.��]D���h����nڵ0�D����P:�DA#[���Ex�r��������<��P���^ё q�f�$�ɾ�=��XK��C@�*y�Y7+�������pw���Ic,�Z%銮eu�-5���s֠43ǥ0�������g�6n�-�.����|�G�΋O𵍫���E ��\��|΄^]*�T��si�u�4������z�\�t���z:�r�z���瑱9Y�-ƐV
O�+�AVF�VK`٧~��u��N�5P�=:�G\� ��^�E@ʞ���Հ8l���L���#��)�'��X����-�?ܷ�޾�?=YcU�mD$CAi�o�{���cY:,���� 9$�lJn��:�q���A��` ��ۈ��}�RB��� �L���~pB��c�ty)��E�ǩ�̎�����LU��x$��~�3����Bg��1�x�e@2��ގY��wV.����ON	3�`�{L�ˈue��p��)��1���$o �M}�R�I5�,p�561$����kd�W���;�b�s:l�k����Td��.���cYg�IG&��nO{3.�>����zK��u�p@PԾ�pee�1a��D���kWs���C��ЭH����`v [f�9Z��+�}��S{�M���ѣ��6k��4�Pz�Id�i*�>��'�j�r����e��䒶�3�7��O�N�7<��R��C���[R�C���C�Y�$��+9���5Z�2^"���<��)KY �w2��m�
�0�F8�P��cC��{���h����j��l%��ol^�x��=��{��kLWAC �3�8��O�����;��A��Z�~̿^�U�ɮ�%3/Kw#T��-&1�jn)z��:��v�Ḧ́,n�29�]eט
������}��<\@ȧ%���>��R^�A��Z��Nm��@+W���3�Cd��A�s����"�%#Tr���EQ�ة0�H�yA��}�6�]�P~=|���\��I�L�R�מt]M�;��o`8��O{��|��g|��3�|{:0�x���G{�"��	i$�muoAu*qΌ-�wW�G���o����'.�,���f�~5_	�d����������M_��m.�=ʮ�6Q�Z���B�F�68�*�o���H������=�V��?O&�T�a+j�im�������{�p������{P�P�A��YS�a�f����L�N�E[����1ޢ\�T��A����hj6��f�?�;yBQ �0�^�]n�T�8��ʯ�-�I��r�KcЫ�$��<R��M��lZ.��9�PyӔ��&���7̰|�30���FgO�-��3ZF�{O���$�n�mzV��-|��@�k�W�ҴzWN�F�Ҕ�i��KwW������zГ[��C��a&�AȮC��xި��N&2�K���=l��̄+*��A�)��3��v���Do�R�/���ڝ���V�����
� �hf܈�$�"KҴ��g��
��h�P��!H��g���O���fӉ*���a�)�v/iH���B6с٨|��XL�U'$Y�+��s�E�������f�!�ϯ���mY�/j�9�^W5�0�T�7yu�s:�7�mA�8UN�5|�	�Y4�����;oo�� ��������f.D��@nHŶ^�|��V�2�@x�cA�V)D�EP>P�a��V�8�a�Mg�����'�7�]rn�_��a^�RL�5M��wc,�8�s� 联͉GI)�Z�0��}�̎B���\C�rNŚ�9��"���\M���C��։�>U��>}�0��i��+�	>(�W��@�IqMs̴nt����t�v\��G/��v8*�����c(.�i3�I�<�O+��^�jn�{��<�aQćI��Z)�:GYs4�@2��A�W�Z���W��L:���\��J��^O����ì��6�^�T����ວ�V[�-����Ea�?�|��џ~-��Sp�톟d��N�UyH�`'K�df�T�q��!������P[��@�)!% >�^]S:g�j��O8�^:QO��r��x�o����q&�t�W?�[Ďs����%��!]@�&}��=S�=n�#�N$��;T#�� 	 �{g�S�:�{C��TA�}�5`��)[���@��V����FW�m�*:�����-*ʬ�������]���U@�݁����b�n�,Jom���}ݠ�����KI⡑���^��ᵕ}��x��4�\�Ua�|&��Ee�N�i�H��Q�Luv��z�|���A+v��"�u5x�kTK�~F�yi[ۖ|�5-�EU��N��'�<�ͷ.��^����F����R2-���o���SQ�ٗ���J�a"�|�w�������;�8��=U��.�̝v`.�\��yl�G���9��h��lb������=;.h��rc�-������ ��.�dU�z�E�l
x���[a&�b#nr�Fv�k�����������M=�"KM�q+�i���5w1�F��hG���\��k�%y�]� y���&r�ËL^9��_Qk�a��c�uZo�ħ�g�Wa��;Xϲ�|EdȺ�d�^� 3�����?2�T{@C\u�c��`���q���z�
�2��F�\0�g]y�)5S� ��_��+�j9T�7�_�A)O��-di��O�;�9X