��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� ���L�����I&V~u~[rR�C�XT���o����۟�V/]�@�!ӁUټ��)����؊������I�Xa-�w�H}�T0�me��|_��������M��)��H�BK���G֓�r`6��Lg�6�ދ��׌�ŵ�G�0�2�!�J��c]Mw(�C�����Af=�Эh�c��I+ݎ���O�� ��^1��0s���=9�߸K�V}9��^��*!�S�����p�QtVx]�����S`�)|e�_R ���bd���_63Y��UgN��l��"l�����I�Gɏ0�4��<vT�5���m�༇�µ�U��H��z�4�n]����-R������ބ��I>��L�� 4):E���V!����Q##^W`(�
�P�CI[q���Y�ӕ��Cp�5뿳�p�3� �agD oa��EčgF:K�=/��R��MV�ٳ P�"�:����Zk�Y �{��W��ϗ��ݟ)m�F0�XFk5 ����V�ӹ���:>�H�A_!��K�� pxH���КϿ''���H���%��?H�} VL�Wj��	[��WUt��6(2�"��M�2��d�)��*>\o�䝮6g̍�u&���;AV�{joНgl�z�-{@��oߕ�����W�S���i�f��5+��l�u�Q�vdy�-u��D�d�~�W��QX,_�_�IZ��E�]���v,Ik�5R̅<	�{�B�v�ū݄8��Nf�x�L��_��amY�A�A"���g�.��0U�8W�Y5sgVu�e��s,�	Ә�׹�+�YŅԘA�����n�'� j��>�d��(�b҃g��X#Q<��\�dK5��t-Ո�x!�17�6�=P�tDAb�\8{��R3�#�|�wb�����%١�f����1��_��yz�Jx�W����/��8��uܨc�3+��R�kW�P���**�ȣi�s ��"�f�Ҁ���K�M߲
�>��G�%P�:���#O���t������l!BE~gz���G%�wlgV��Msq�X9�D�v<��_��b!�~!����#(�;��C�;�l���7wt�C z��3�b�F����R.���`\�h7�.�e���q��4�K�qg���<9����G�K�$cQy^=��� bJ�=wD�����H�걥�5������b�>�?.)�l��S
��]�7'���d߅#Gn^ϥ����u����.��Qn��^���� �-H�
�4@ͪ�f��Yȏ��++�0'|9�e��0=���$\�=���W�M�<��_d�>E�QgY_��-1im��"� ݌��*
LJ��,ۏXI��q}��Ked�qE����� %I��E�ӽ�b�*7�&ᗯ��U~�lXQ�	�!��3�c�n�Y���Kgd�m�I
���yh���F�2(��q��ZEL:u}��W�������Il⊹j�8$��3�b��W�ݰ�U:��'2􍰱�������6Mo���i4��ZF���Y�7C{7,%!�8l��l: ��y8�W��Oi��汹�G�/�y6�:E�s��ڥD�V�ؒ��������ޙԖ�{�:��y�wJ�PsQ:�Ə�F�q�8M���I��Ȋ�L��4��{�:M�O?ut���{Q�	y[W��w����>z����޾�{y"]'jr���@��]��Y���ݵ�X
4C~#4 )}ɋ�	lxj������-�ׂ�5ov�	ۊ�����i4�;��rՊc]�t�n9O�9�-i?
	�b�#a�,%q�TxR�ų-n�
6���﫚��/��X���Ȍ��j������dqcDk�z@D���lsU�Z�H�T��2v�ڜ��f�N�Ds.?�"���0ӿ�t}bHG��t7�XX�=T�񫻻��3%�(ÉR1e>��$�����ajI�W��������-��!s�͛��.{���J}ր4ZI]1�5GT����.j��ǯM�D�{�6l�eR��Fƾ���b��A�[qX,��A���_O�J���aΕ���5���2�ǜL�tr�Ze���^ 3׬�, ���(v�hT�K��~�C�b��* q��QA�t��]:^:�%�b�~ݶ��
�C��#���ڄ,
�ʿf��G�F��"�H�?s�~y
�}�Jb�DV)��xf�:�i�-Q�`�.�1��P.ؔ�B(��N��j�ח��(Zۿ��C43���|�KdR�u���X��j�$R���`Q��:��V-� j��>�T�
GZ01���fbp2�i�u��;���*�޴���9��i��+;��%��Qt����C�_6��[<L*��2)իO�E�&>�G1��6}�V�n���Ɗ�a��S��ρ ��yԥRc���Ǭ�jw��Xk������
  M�Ne����H�N� ������ɥ!&�8tV�<�7��<G'{�f�r��A�8ȿF���&�agqV���o<�K:�	|&g �g\�_���S���n ��p�W���<�����1���4�B�yvD���u9���Դ;}\塌�ܧ�vj��;��c1ݶu�T�U�(Yu�"~+6��)F��b}���J�X�����}��|$Ƕ��(K/K:r8y` h��*j�aqE*>��x��4���Y��`M;�;�u���h(�Y7=?���n����U<�0t�Vb��B%#n�?'��tz���d16�GV�ҾX�"5�y2���q����tբ��U��2�:<�D{Dd���c�Պ������6-�p���"�i���z�`B[Х�s)�����Z ���V���[���"�_���8n�ZH�w��
��oף7||�i:^Y}ٹ�5����Α�r�9�«�G��L_�B� W�lDȋ�q�+,v�>LL��U��*��I������Hb����,�]}=H/�X�����=��bޒC�0���5��HB�������qg��׈F1�C���
��r��Y���Ȉ��^e��`!P^�y����w��F�i�^i�%�ES���\���F*KDe��k��v��,��"���z�N�Ӓ��v�~a]�!��4��F��`�
�FZ|t?��'�:Pt�,�I,}O�o��̉T!y�����<Tq�>w~,z���5>�BZ��A-�ׂ�j�z��K�>	�x���Ξ���U�M,�t�j�j��K���dc�4J��u�.\Y$t��r��	nF>�F�&��a�_��j���$M�l�DԽ��y
ň�a[�M�����F�-�p��J����64q�~?�s{އ]?�Y�I�Q��JE�u�,eĩ�AՏHXO�F7>[0F�jv^�J�L���]�
�㳡��/������d��e����DU