��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|۶��-�E��ĝa��v�O��hG������g9�ϭ&�;�C�hf���=����V���K��1�BVS?�ם�Aq�I�3������|wW�!�b6�f�[#�� #e��KF��WQ�>v-w�KNX���;������!�z�QɈ���Ҕ�#���hZ���K͍+ď�t��@v��ķ6_���7�B�F������Ɏ:�� �(�%J��{{�t�`��/�1��,�d1�쩜m[�S��^CY�_�b,8�/��>��e�|)��_]��uYn4������l�[�ʣ.��`�#��D��S��2��^�J��V�շ�"-1��ùS���L��DgZ��i0BWE��� G֗��/3h�+ ��~DLNSAm���ڦ�ŝ.�� ��_r�+�;ɒ����6_�j�7Ħ�W�@����(�IsZ��^h��p?�̊G�/�f���"�	_l��&�ԭ0��ub�}�Z	{��R_�|�DKB�a��X&��I��&�Ax�'ʧ����l:>�U�ez��{4>�Ӓ�O>%�$|��g0c���|�T�#nqێ��(���H���������O��m��������X�Y��x��wQ�"����+?�k�yKyw��`�Mͅ��G(2�J�$F�zRd R����)�Y�/�����A���7�0�4C�I4I-JJ��X����������-�t���*A%K,��;�;%Y<��.�o�z��++Glq�zK8��.�B+�1�wŘV�o��c�χ1%�*҆g�����M˺t-�����æ�?U\�b�4�1�����%����/
�N3��K���#a7�4sE+W�j��X��ˈ�����s�f���.fE�q�K������B1�"�O�H^۰T��#���.mo�` mvT(��|�%�w@�:��/��~R�����������8��2v����u
Ɓ�p��&q˨[/$r� ��+i�A�7@6�c�"L��0ϣ����P>ɺ4Y��*�5�q�c4W6➾�2
�y�� ݖ�<uͣdo���`Z�Xd���zG5��\�L?Zθ��\{��P��z>�O���݆�|����RYxL��[��������u=���1y_���o}ZC���F��\�Kަ5睷N���e[*'���p��Pm,�zY��1�d�/��dG���D1
��4������;YZ������4�h���DǎAAd���~��i��8�Ld����w�֯l��N(w��PMUv�7ġi����R�I���հ��	�frFX{��:�����E`ra�ǒ�=�K�7vF����'(��K��z�s��=��G�r)L�L�6SP)r�l�Xv�y��Ԭt;��2�RU��{ᑐ"�h �b덀�U�R�N��a��:��xbu���,���3U���w©��o~���bq��.=�E7�E��9&CL�Lދz/s2r1�3��Š�*��M�:~��1�\Bv�S������i�2 �K���[ۑ���=��HS�UwYY�{l�iTK�m_���Л���A��d�m�K:����U����4ˬ�<H��StͽI�<��5W#Y$E�$/VE���h@:��A��y���;N}}@�# ����s�պ��4��]�z�_o|j�E�D�R���g*V� u�G5	�p�9�[�*�W5Y�e"��<Bh���t"K��W/��	��T�K�/�f����|b���LEPt��\��B�wQ�L���G3ǭ�P����i1`�f�V�i*�<��fN�xl���-jweL�al��n~�+3R_i��Zݚl*�BiW8����4Ǜ��g[8��
/fԽr�	��69Ŗ�'��q��>;�D��le�"2]X^�@W�W{} ������`���РY(W����.�ۏD��z�2�@�����v/�'�/Ŏ�(����Ǆ�-�+���/�;YA�r��G}cX7���(����Fy���*��g�0�Wރ�{���\�9���3g+���{	_�XCz�4~[:�����{ *�" Ǿ�)�^t�J����u��ý?��Kbc�A ��C	z+��u��#~�A8R��/ǹ�~�Ӂ�^Y!8QR��̾ ,v0��X}���:�Do���A��\V���~�ZC�/#j��n��{3���2&�cZ�5G��V�W�Y��
�Viϩbh#�$7�G���t�/�g��a�/�鰳���6{n�'^��)'�;A���<�fj�q�L��]���.9��_����q(�A��j��`����V�^�iExbq!�CMD\g�������
ɉ��d�u�Vyjˇ���K%ps�U�ߖ&�\%����eX!��C�:�W�3��@�&̹N�y���dxT�a看о�d?��j�G���������Jc59�J#�Y%ɍp��<��<{t"�5�ϯ5���� �ᅭ��@�N�ώ���0��?�J#:<����6�k"(5?J	ͯ`@2��?����Z� FV/|ښAHE~#<�#�� �������r�� �|�+�=]p�ny>�b���	+�6y{kq�=e�\J�j[�H'���p��=�\0�SI��Y�J��9<F�s��^��;*�-�g53��-��᪛iq�A����z��W���R�>�?k��%�H��.���)�4�aw�zo�>V��.<����\#kXn�P� d���{Q�K��7����˛�D�MS�}j�*ﯺ?������D�ب;»fnZ�3���F��O
F�=M�!P�����;�9�АG.�-�Z��WU*�� �Ŏ��0f>�Bw�#5��,�X��Ӡqr���č�/}���q=�	Q��
����j�F]�$Yi�,�@%�r��:�XWx�~��>�nO�>jX�ɝ�U�~c]���,��TT�����eJ��}�ᠱF���e���L�W�m����E���g�݇�p~��Y�[W�j�D�}X.4ΛK3��d]�x�����G?-�$�'����b��$@Fw�H���1���KO�{�
��W�_�����Kǥ>�#j8+��z?��x�pb:��j��M6x����=�ݲ��h�xW����/Е/y���d��h������C]�ܬ�F��gAodn�l0��Ӳ�f���(����䆡��!�F�[Mr�+Okk�|���F0HǂT�J�8�ճ�Nű��bS�n?���T�V���j���з�O�c�^����������էrZӏ���2ERɊH!Ur�gݴT�
�k[��2�Y?��:�B�'�D�܃�!�lM�p�Q�_Xװ�r�z3~�C�5� ΤK��Vkl�?�4�y*;ܳ�#�QC�;��Ż&p��fK
��wpE��]�1f���í,��g�K����]�F�V}p�����n�/?=#6(��CyU�/�d�����~�$�ȋz4𫌧	IVG4o�%�'s
_�`�F6�z�A!�7��e�{�BTNڜZFE&�.��� 4����w���c���\�EjiY��H,��XѲd�l���5{�c����i�$�4A%�[�ɭo�Eϩ4�L�e�n]��&����ũ��(�ʖK<�K����=������T��־Ò8W42�0�>4HNLһn��춥��tF����b�dVf�{�������j�L|�'�Wf^�*G2r&ĕc�M7 �UV��x��q�4;zԶ�>��ݫm��6�
�=�[��<�L9ݮ�����8����ǻ�Ҿ�Q�O�g�H���Lu��k���ŋ�19es������"�+���tbf]${d+�՘��s��M�[ƥ��E��W��}1g�q����oq２n��:������Q��l�+��ߺX�8�˨��-ru���L�&���F��25}W��x�_st��{��8�} �:;�X����zM��Em��[����:����f�,��~I��UnS����D3�d`������C�C|h�kjy���!3w}����225����.��������|�5=1�YH�|@ *����"o������N��E�4%���{F�j�B������`J����{���eK<V��z�Ҫ��%j7.l��!:fk3_=.��&g/��d�:%���ٗcW`��>�XQ`��0�9^%��4Q��@j����������G J9�u��y>ծхp�{�/�U�c.��պ|�Q�L�8`���$����$�KR�3h������>����&���7�6�!�����qW�4�6��k�d�5�.��K���N�
�Rq5�����b�=�-Mn��Ā�~y��.�9ń�Gw�	`sd�A��8Eϗw���3�ʹ����)�L�΍��m3�*8���_^^���l���"O{�?{�>s½��=|�f�My|��$���,��D%/�9�p$��A�rq����rU�%��ioS��3��3�"��t���H�j<J��=��ŕuHQȾn�cvO^�t�����޿�5M&��w�]+I��;: ���:QƯ�,:ڕ���	
�=�M��kGj6�1%�S}��\
��*�{�6���Y�"�����|O��_��Fk�e�S������9��F"\x���4�bI��/�#E.0�	}�{!��cY4�p
K��!0��H�/�m@�����3�-;;���y��.�t-6�lrVǽ��7�W�n¡8�=c�##X�cg����Z�R�1����`a?�oGG{�׮��<q��ÇL5!b�?�����B�/#L���Y�ja�^2�žbg�3���$cTM�{U�!(�����gxG��ze����d�&p�L�K�	]�I��G
���O'����g&t��J?*=wS9d�E3�z���lt!�p��e�wr���'	��[�6�(��h�$������oB������p�'�*�T=�i�I��RZ2ꌻ�/s_TWIX�@�na-�Cl���h��~*!!��ﲉY�/S4Ӂ�*!��YZ����2��}��
	��~���� N��l��#T��6�:�MQMz塚��;C�6��ب���	����o�l̦F�'d%s���YI�:�E��j����~֟�� �Z\=�"��Y�$X��)@�A�b��n��s2�6m'a=t�U8�0@�&�a����)������9�����m�V�3}�9�~�r��`6ȏX{,�G�'�'7b�$aks=|��DM��:���v)��L%A�|zGujL�;X���������]�b}�c��F�>eN�}��m5�+^�z]&(���d�|h��×�|�y����7�̄s!�li�cz�}��	k,��^	�x�y��Nm=ֱ��2��ٲ���\��%֍\a�������]���11���AIQZ�%�17���ײX��jg��4/s}�ތ{�T�����A4��O�7�GL��̮h���Μ���wl���^g'��;TF�X����{[����4u2U.f�*��O\� �����v�@d#���w�Y� ��*0�!�D�K���Us�GY�v��?,�:�7������*$��I+�d�ǹ��`����j�ǣ¦p՚f2�X�G����`�9kD��du��a������I%�Ծ�3�l=�ݤ��j�{��@@F�b8]%޴��|���<��E�Oj��M���v�-����S��e䉳HZ�����a�5��sI���BB��L �I�B���_��O�ni$��7�`�o/�׹u`�e�ǐ�����#-�L� g$S�%o3��A���VzW���赖P�Wu�:Sr���ah�����RըJt@L��Q-�X�j)<^����f9	-�ǖI�- �;�4���$�f��}��f��)*,;�`�#�3#�=l]s!���u}l���әȻ S�>N��%�ϵy4��8����_�����9���`�a�Ėb3uQ�����졠�qNOS�	q��5�K̩��������#�?�7]��FN��wF_�O��tK޶&��~1C]���J�ڢB��b!]?��m��C�cm�\�����!gK[R�zZavK�6�-���A�)R�c��Y舾ig®�r��%�!��ը�J!��5k�PY��4�� ���/�]\��� �H+�_��h�he�Nl,�V	zo�ߌ���;,)?Z=�m"�c�a�^���sI���.ޏc���w?{uRa�`m���;�����Y���硓#g��`�(�����6�ǸX=�m�?7�)����kx�WY��u���.;��e�7�^H�V�),�����x4������zW�2}��aA�l�,�罖��l�/d����Au3nM0k৥��h&����	�}�<���,�#�ꀀW�D1፭���{}�ǔ�饔?��p]s0i��Iu֣�n�k�@)�h:����+�[
È�q���v�6���Y;��m�w���LJ��c:X���6{��jy~3�L^m�|Ĭ"���"�=��<�缰d'лIi��L�ů�.�w��y8�N]�p�Oӽ�Sp'�������-l�R�9��*4d��N��>@�n�.�t���P{����~U�8^���w��<���x����5��>b�Z�z$�O��Q.4 �ڵ֥��i�ε8��-�C`&��N����@����e�i�q��+FK14��$�Dxp�ݹ�%�cOH'����u�+Bj���0����M!��Á��r�#�(8���1~+�$�p�,�Ɲ� �[g�r(���d�)���U��ð���&G �����b4z����sCw�ow�a�d���g(�e��v�y���A-�	�±b߈�Tr�OA`I�%�<���?~7�����N�#u��^C�����m�ͦ-�`��a�+���s�n{ҕ8��"���F�Z�V�z�U;R	� �����?��Q�#���d>@�\-M�9�2]�/}�=L���Y�X}Ӝ#��A^v��\|�O.YP8�Q� 2���E����I�@����
�����a��_�u��4���U*�!2 .�\X7��t�
��d�~Ii���Yj)�A֧[r[����6o�l�>��G@���lj[�R����㻰�mR��=�;^p������n.% ��?|(�r�&9|9&��+Qx�m\�����D�@¤&���[e��W7W���*r�릻=v=J��U�A2��
�S�Ľ���M�3��)ի���R��IU�* �LN�����L����(1���0�ۼ�	3�!kn�P���[���k���D�n�hfx���l
*LjnVzE��Y�Z֠�!e&�9ѣU�y�n'���U�X��V�j�`�-YV�C�������=�����#a����&�-�ݷ !��#�dB��b>y���n!5Z f�i�����X-�>|*$��8�Z����J����0&L������f1���3�쾃���c�nu�
s�f�N%ЕN��B�eA�v��ʼl�#c�-$K}�<��
~G����d�s`vl�8ߐ��Fv5a������
&��﷜����ّ��N�"59Ѓ��[�ٹ�r��Eu�6��gK��9�
���m�K���T7m�h֒����䇜�Uk�6���;��VZ��c��<�����jXc����Q��SpV��G�o%��[Λ8m����c�0�m �:��;gl}�#Tv�ܖ�%����]Kj�	+��{)a��	\�����4��F h-&z��g����L��5�/�2�f 4ԡ��WQ.�J6�*��d6�1�Q�`I1���#�0����R@���(�F:Ӓg��dq��w3'�y����6~�ڲZȪ /��.*	I�=��wq��O�k�7Y�{$�`B{�����<8��2�#�h]Ǒp�7.��R*WM������"��89f���%O��	��ˉ�o���o�^�	4��� ^��v���2��U`��G��|��б-kD�#�?'A�H����|zk�}i 3I��������(2bȺr��u�81&^��A���4ERK=�X=��)A9���'N���h�>q�X�F��a���W�ѓ%�~��-q��Z����A��r�>�WK$((yP�Щ����S������H
I�W|΂T���lV������k˥��Xm�/(�(.Ft�i��/�8�<k�뱄>�{{T��������!���T��r���\�F�qp��Q�50f+�LO��.8m���#����7`���{����z�s1�02����G{��d@W"�Q��/+�N^���fx�Zc;'8��3��ͧ<���zBm�Dh*#v�4�"=_�xH�}���`n_�ьK�a�;�a"�Z-�pd�-�D�_�9Q���[�����D��J�Y@���?�����@-hP���C(��
�o����r7��o��Q�ȸ����Z_�����Z3��sS�N:4J�j���M����ض���@����(h
Y���U9 K�7.vL�IuV��j\)���R`����ݒJ�n6�/�ԟ�Q'�3�(�o\����pj�K	9��)��;S��q͠?7�?�a�$;'�j��:�\�!�.5oQ	ni4�W�4|9R9�/�����P�}�t�����vYABz�]8Y����U�XhN�G�����s@l�䃲��\|��7զt��>wut��
��J�B<�~��0
�s���M����=E��}��<�F��~�Y������o�^�p����>���*���w6COe@�2|�b'�ܘX���U�"�\G�q�W��V�iV���"��	�!YR'���)%jyR�-^n��9Ηs�[5��J���'��d�2n%���S��L�d��"�g��(0.�QAQ�(���;)�A��>e��*�-J~e����F�&E?7~����h�_T�ܾ��E�n����Y�/h�X��R��F���&�t��:ѝx�$�<?��W��ѝ0��)^~�
F�x���F�}c��Q��N}':}�Zr�4Ι?���o�Fe�+�.u�CfA\�����^ y.����cx��!��R��88��y��^�%�?.�E� �x�\��UU ��O�R������sxC��I���4W��)-N�s���ȏXZ�̀'~�#R�����-���'��K��" sƩ.����+�O�mo*�E�a�ߘ
3tK&z�vML���fz��(���)�l��5��_���g�>)�)��[#���
3�a�����I��W�n�@�+�ނ��JY�y�5x��
-{J��"C8����R���\�kLO4QWn�ʘ�r��� �iJ���/w�rkT"��Bí�,%a�K��\@�J���Qb=�KfB��=T*Dm�yBH:s��������� �sfᨬ�`�KG+GŠgi���m��h�*��*kkEVǰ�N#"n�7���U�2�r�o��u`����@�f�Qr���� ��(�� [_���G�ӻ58���xQ���N�Ӎ���C�ӎ�� ���e�Y�[.#��{���KXM¦
�!�=�/���/�<]9�.�c�D����:ݕ��zh���f־uz����lwe�{.K���)c����;�#rd%"������-�ZD���Yr��MY6)F�m	K)�{����N��
{5娸{�����0�Zf	�d�(7�ЕsM���c"Q�&}t:H�7��ZP����&7������ia�����C����US	��5挛����Fs�\��9�9������"qL~[��I�=B�i�x�[�1�?S���d��J|%A��m$����3��&^-�EL%X���)�+c2Q�Q��Q�����	^[���j�,��j�(�K��Jq���6Gy��JI��Q�cD�����1m���c/��ߧ�_~sw����/�$ZX:P�%�R�)(*�����*����K�@��vr���#��	meTHt��'��EͰ�F	@D�Kd�RX�;����u�Z�в���u�7���k*Tc���Yhn�=���[\J��Փ���?�yWn�+Wb�&���d���p�wk�p��Ə�IPK��t5)��_\���y1{�ٸ���n��(x�m���'7�_[�x������Mz�ZB�hD��8�t��v�a)u{b�d��2�c��)�� �����H�ֹ�z�=���줒����P�����]��}P��L�C�տ�o�V����dx1�� Q-���Q����8��+�����hNܔ�_�]")��K��S�ڄ�O.���G�v��.� ���J�Ý�<��C�C�ϘZP�i�J����VyZ44�|^HQ�Kf�wX*XW��R��������]�kk΂�$������1.�s�79�f1�;�b �Bݵ�'�$�a����dsb�L[�v�ML���n]�����{X��4�@���:�x�&�C����YԌiSQ�{�W{"ʭ:7��1��㬛�ٿ�}P�䵷�)n��߭���L��Iv����T�
�D����.E���9�qz����6w?����ۘ���=�癟���$���?� hp�iW�;�[�E�#?tu���V������uH"m�5s|��i�.I�e1�hSc��Qll�����p��F������!��E�����&x�����`�I���˴�!��ݛ�ս��r��]Iۣ�+�� (0�ő!}#���-3=�#ˢ*�%+#r5y�6Mn�@o$�<Ѓ쑦����A���{?��!!I6�"{��tE�����Z��ԛ)L�:В�Q
�Ԯj#.W��C �ݼ"M��TR�B��[�IR�7�����c���\U��lJ��9{F�^�����j|Q�f1@��=�]�]f���?��A��jX��*q�L�5L�����S�������������Td0�Jhh���e�\�/���[�-'�}uP�9ĕZ��&��=�IKʅ���:��{�~��j�!����I�~���)����ܙ�u�'7���Jd����M�/�]�O� ����4��z����H�@��~-�)����`Z����\G���hg��fXL�`ۍ>ġ��2������.d|k^)B�Tl���2N�I�D?��c��G�"Ǐƈ��HI�\ݶ�\�02l�Y'T�3��\�H5��XYܤhHih�\�Ӿ��Z. O��׻�k�<_@��s�Ӯ%�5� 0�r���\�)���w��E�]A8$a-ʪ�i[oqS��.�j�Љ���+@�C\N�F�c�ʘ���<�O�*�@����b��R�Acٌ�Z��U�Y܌��j���*��5q����t�|h�u��nB.E}~	č���������U��>h�i"�Ќz|��̠x�e�_ǽ�	8�>,�9,��@+өW�_��=Q��n���~��S���S�X�Z��m�T;ᖦ�*�ڋ�zH
)|!H d�0�sT��P��R�o�s��	�8fѻ^���#�Y��8FXa5�ʭa[6�Y5مJ��؞�^̬�qb���'���Ӣע��jF�����lF�(�sP��\Yd���&I@��Y;�i��c�,�[�����!�hQGm���hZ(i��ViA�Z��+�$���+�2u���<q,Au��o	"q3)�?�u�K�g�[�c�[�H�d�!��*h�������� �Fe����(VFR�©6b#Z�p�oqچ��#��^�5d����IQU�2�fl�Ij�E�3Z�c�uJ*c���jk��m��͆A�����Ɇ��բ}R�)���8ŕF��v�\�)��+�o�f��p:O�:�⪰�*H��єZ�B�2�-Gq�|#�?f�\�-݌4�z�̜��[x̄�QF@`��xkXp��܀~�&{SB�s�H���\�$�N�_�qE��/�_��}x>�ωV�Y.�M³�K�C�IP?�i�Vv�?h�)ّ7W����`Մ<;�sh���0'��VN�͈�u�}Dn#�6h ����uE�޸��.]:��1��87��
�G�q,�Gij�e�����f���N ҇�N�}�\��7�����U�C��s7Q��A�]����`f�73@X����ܑ%M\�uI�c�E	��3�$�Cq@��O���؜�f�m�ku�9<��~���ݿ�&�L˰�#Gϼ�a��6b������%u�e/+��Q�0P��$D�O��GC�/�H4>e�6~�8_�g��R���4�#�Wan_"7MFV��G�Ɂ��"!K,f?%ڹ�W%�ݪ[ރ׽���0 J6� �R�����C�6$ ]�}�;1�p�f������<���PD�Hi�Їù��Խ�o����<)Ԋ]p�H��Ƶ��������ɯɒ���=H�����YF�}d���`�L�3r�K�!��;�p�>~Cb��k�'=�4[�,w��3��QC���O���"��PDl����qD��Ҙ����v_�+Y�M�]��?�����XJ��:E����h���Ae?Z'����<����^��CÿH�&˙��CJb������My��sY)�r�<��`�>��l��X^�zP������4=8�n
"!1c���i�h�c0�C��v�p}�>q���;��`��2y4A����~��X��Y���=;J(��l�M�n�9��U8 �;$�kP�ދ���ZK����|6Ao��*꿳�u�G�Z)>2�V��SӞ��2ޏ��l\s0����	Gt��Yv^��[�0M��ap8���p���t���A��Th�b�ChL�[n!E{�L�.������#c]m���KzR�ָ��N�O�k��}���ӕ\H�p;�B��)� �&]���z�>1�q�k+�[z��0�dX,��O�9%����}6�9.�������
,�4E��U^�Act������u%�r�kseH	��)X���ω��B|���۸��qNtF����i�ԟG�XBˍ���Iyn@�b%���
(Cgg�**�f	�� ��T�*2���S-�mݽ�ʲ��~�v���]�;O�e��"�
7���Z���-�!sm7j0Q���~N�u��,����+�� hJ+P�w�չj�~Fߜ�Ȃ���~�sa��]���]X����+�Q"9����P��؁�9���	��7pK4'-�h:���Ex��%���<"�wy4̜�(9��RX�������-����h0�gu� �ZC����^WH6\�E�}�������:#]}�樂�����́3�%?�0��:o���@T�I=&$z�;�`�l��������|~��)�������D֗7�-g�:j��`�N嘺�V�L��5�MM�Ӳ�J�tyR�7��'�*�'�+U��R}��>� ��!�j���,Yҫ�xF�M����+~�q`��KC�qAl?ᒘ�;nS���ї���I��N�������B�����H؎�Vj�-#/���Z��]�۴ ㇞�3 ��բ��*r� .���B���}�� >%V*6q� >�	���bOӎeՈ8�TŠuYP�/�W�TҋB��j?��߀�l(��mgSк�ŝc�"��DDQPv}m`��F4����D��q�Q��[&��
ˁ�I_�=Ar����w0��1��y#��0���N�U�p�1@�<�$viy���ƕaj��罅ŧa�O�|8o�O�=�U�\x�|�a�2.��@��l�kJ�j3k�TsPW�PM'���v�N��q�`*����|���t����-��H	�B*�W�:����]�(_М]��$<.N��:���(����\-=�	}fUo�O�)}^Rm!������	:x���|�PIj��/2
D�Ύ��A^>���o_8{�M�H�/�Y�D�+O����	�%���^Ģ`a�5� R�C[ƴ`e�{���J�� Ƕ��7�o`M�O���=(�o:�D��Nnd���LŹ�)�:G$ww�67Q��#�Y���EB��H�A�O܌G�mg5�8�NU�(�k�	�E�=~�̧=ֱ�ƙQ%	�-	qj
0�_����;z�QМ[�jݵ���4"�̈a����i�_��^v�"M�9����U�V����V2W��y�[!� Z�K`)B'��y"PSօ0��<6�gk~�a��m�ȝ�5p��B��n����eR3�둒���Rji�N7����}�74<g��Á�i�� g�nD�3,�s����dHP߹M\��E�DJR�m�Î��:�80����[D��dd�g��y��,��
��}�Y)o�9+�&@�'�XS<�s��t4lxQ��_�����Ґi��Wm6���Y�9.��b"��Rc�����&��Э�gC��(��M��`E�ʡʄ�d��r����I�|$~r&c��֍�W���yU�Z�n8��iG*��Q����)4M�_c���T|Y��@,���LwG}�w�;�+�@�Խ��م�л����R��rr�=���ؿY�{֛M���f�����"��許AƆ�\o��ח~<���p�O�X��$�C �g�_���/��e#�v��A694NVV�5�z�=(%M�u��Mǟ�w1���m���*x8�.���zMr��ܸ(K�'5ߧ9v�HS��װr|����`)jů�Y[{�q>��}�ހ����QQj$S�yc��L��nJ5<�ϗ|�ꐫgܺ7� Ͼ�k����� >W�~�)>�M�l!�����Q~���Ik���f�)�ͱ%vϋ=_uT�l�"�L1x�'���5��nE�Ò�*����	�bb(�aHP�u��!zD��۽Ri�)�ޓ5q�4�o[���<8?q���2�\
�:�pg��O�/13����3y�_�˝�Ɉ���� ��j�I��v>�(�+�Ƕ<�������F9���=�[r%���ǹ�r�<��\죲fS�(%�|�"�<�GdD4�{��p��l� x��������a�Be�tO��i�5�2�fHJ�e����X"� ����Sc�*��l%�4�_;9��܀�X�pO�@���3
O1�C�8?wːg4���7<�a��\�Kv�kn'�m1��D���2"�d�ssܰc�=���'Z��OY��<C�a t�"�Ӟ&�^S����~Ǣ�F��z�{�jT��t�@�lX��i5�u��5x��?g��G"���hR@��P�?_��j��,?��x���̽�e��5���8
�V\=��Nj��f��D�����!���"p�d�	vE"r��Z�s3:��7~t3��E�=~��Z�/�g ����Ox˄�=R�!장~>=C�=+ ���Q�b�C���/ ��7 2J,`Q'-�.��'"[w�9t$y���qC�T���^�J]�Al�xAw�����n�W�_U�x�o�7�u �3��p��L�o����u,�e�{�޵�oL�R�`�o�K4.^	Y
5cT��0�i��8n��Cj���tࣾ����w9���U1B����<��K,���RM1����x΄�Au~ �#@�fj"�PJ�8�1*?�2D����`fHoS�W"�S�Zk�Q�){Sv�=� xdwq��QQO�P�zt��`9��r𜲍XZjN��ň����l�9b,�w�I�bt�6����o���d���1Ҩ�h)@��7�7J~�_c�+�p�o�fŖ럤�ِǸ�*��n[Y��ԡXd�j�D^�����LH1���*�^�b�QY���]�|�Ŧ���U����%���no6�y��I����Y:ݘ�����υ�?��_�Y��OK'2�������矐�Љ2�'�:�-�n�N�&,�7^�spi�K%F�AB��*u�Hm�ZV���n�b���aO	���J��qJ�l=R��"|���N�Y�Qק��^�Z�88o�8G?l�}��/(��4��2�1s�w�{W;���l6�9��5���I͕���^��	l5�g��O�/m�m �Jf!Ƶ�>�����;���1��:��VO�:�D�L��|�g�f��$��@}?��|�X��'*�Y���hDigLl���n�+��6�\5�=Z@;��V�6:����T��>�jY��ĭ��1?<qj��P�j@�<�G�C��q�mM��i������6����s(@!9l/pZ� Of�3��*h����^��Q�SQ���1h�\��<��$Uz�K�Di15�:���^eTfH�Q�E������h���ؓ.U����NV� �x�v��V�l�@%��m�"�Yt�hj+��bѹ���M�{�Ź�C=jq�G`��&��������ܬa4')�F��|���9��vt��&� ,�?���N��^�6��8t�D>+n�B�SR*m��2�mF�mɍ���o�T~���$��[���[��X���8Nb�~,{�p
+̥���j!�G��v�	$�)���;|�)��e� P��Fܣy<s��\���/�i�N���H�p�\l���������D�,!��/(�Kwi���=�Y�?��̾b�Z������_o4)=�Ov'�l���K&� �87����s{����$>�8�T���)+g�U����C�������t\T5����OfF��-v�ܞ�Zm��텹[f����'o�n��{c���T�� ���)6��N^�`{��˷e�v,K����#���R�w�<��=��JH���?�.�{*6LY�9���Q�ЕΟ�� tȻ��rC��=D��:�o�ss~��s����c�+�{y���C|��U�;����8S��l��m��쒅�����t��!�l������`^����=�7����O{��4�@��s���s�8ܽ\|I����o��4E����/�?l۵�ԣ_.�ې��'��V/��Ϋ
�fB���Ly��	��,��/1/��uSp��P*N���%���㽷w�^�IhW��xq� ��f��hE"�l��7f�����C{l��q%~b�"I�"�,&�=�p�p�3��`���0J��$k>�|b�2�����@���%�����ZQmH�R��K��x~uy�:D��B���;�����h{�qa���m9�&�W��I � ���`�X)���[�u�������m���Q
��`"f�#��<f�ٕQ4&��.�ͦ����8(.�b.ѕ<jW��9��p.���YBKE�`�տ�Ud�§J;S��A����N3p����`z�ǂ��~��������i���!d�Ż�n_P:���y��K��2�k�H�Ӂm��\7��т�0]xۈB��O8{�:���Qg�D��{أ�w��1��7�$%I!PIj��=��T��yƻ��F�-�|��9���6>'������2@{|��~D`�:��g%F �ϩ:�>l�j��5�K/!�j4:�����Ѯv�#���~b/�܅19�D͛�;t�8�!x��s��E[�����7���� ��1gw�Lb{B��^�apc|��4��w՛�����v�ku��MY<D��_�ͣpd�c��_(q���&�L�&�>�M'6m��y�{��������O��N������S)�G�ݖ����m��y�4	��4\j�,��vӵ��з$י�2��� A9v���&��{�������.}B����ʮt!k,� ��k�r�ԿxY�\����]vF�)fx(@z��J1��KÉ��:���׺��v��W�y�)\��¥[V��mVբ�%��i�H���i�+�rN�K��!<�֞��wޕQ�+�#���=h���hkL*�<���}˘/��e���m9�Ɵ�2&����;$v��?&#uU�#�;�db�u������� ,��4P�8������B���J�������a��
���9�֋u4J왘r(׶F��K)��\S�Y4<��\����Z2cn��&$��^����|��|��c�^�}py������Web�N7����=����I�\S}���oq)���J���䯢��"iI�T4%���/~8�E�6�
��t(�Ҙ(��Z���ĭ5X|��u�of��]���O Ǚvͪ��[R��X@��m�(��.������c�����S�P�q�ځN�ME�������'�������L_�'͍:����\j�)7^�5cE>�S(a@�Zu溼�|7�m	d�Q�U�X+ُ��0m�Wm��e��`(�mz%w)�VB2���t<�m�G��E�k��w��~[hٲ�^L�>�x>֣�q�s!��J�8���d�D5�q�� �����ްm��/��;���l���F�9�_�.�,����HD^׬�R��s[ρ�o�������f���#=�[�K��i�E�R�f��n��x�76�:�z%SؕԐ�Ե�$���e>ѩ<|%�;zA?2Uyq�欺��-�\�� S��X��5��e�L���)A]|pN�\>�� ]���vl�E�����K����U��\���mqoF��4+c��c��KS͝��7׭���R�Ǖ���gh/@ü�ޛ���;�)�L;9�/���'}lIK0�^�0��ν��3�j`�'kM8]��8xJ\GV��t���>�ߔ����esf���y�� �Q����|q[ɝGd�'�H��Y(��`Yۆ�p����0�,�QE�m���7���ƛ��q�^�ӊ"�U���,�>^/����w��M�I� m[�e[�܅ܬ�*������׮w�PZ_ ��r�Ǐ�7ⵜ�a�]��ks"���ڑa"q n���'��ad�Ht�p��e]u�BX���O��~���Ms�^�������F��AC�#�Y��dV���2rve�76u�)�x�|��|K`k�OwSz~�
*���S��v2�PG����$-������ۉ*� �����1�@�S/NO`E�/�TK�'yC�?R��'\E.��&Gc�Z���(���2<�IK�C�q�U4e�8�����2nF��a3���[	��������KT<�?x����~Lw>���sui������R,T�#3N.�D�\��'�+�W&�"��3b>�\D�	F��� �m�ԩe8���Cw_n��7�Q������u4�i�!�m�}�4��u���Q��n�(;��W;E�v�krA�P��x��v��3�@�3�("�N�q�rq)�j�#�JZ������d�/ȸ�#�:ŰWDS�<�pNn�U�'��r7���o��+G�8a	�{,�<U�?p��&��-��/�W����qQM�<�&�?�+Mp��6+��^+�������,��w�����#f��.ZV̲V
��M�gߟ�} �f�ɧ��X�����D�r�u��HH�1�� $��a�lf6J0�j��r�U1�u��t"��af<Y��-+4�>\#`Vz��Ʈ9~x�f�"�y۞@���C�e@e`�	ZHĘ�ȵ�����xw	ݹ��ij#��h�k�W�!��^�� |��ıS� 0n���@�v�����m�]):��V���aD�:ٝ100��:��Y@sx�|)1!;��a���)��vX�D\zx��Վ���~t��sw��ۀ}�/��M�d�*��&z�a}������:?%ZP����:�ρQ�w=�['w�>"�s�g�����j�#FU�{P�}�Ϩ�T�o3� ��'7��>��z�܉Jdff�ׇ(��)�9��eGr
�6xv�m#M�:���b��Sz��W	�^&nd��z!�}����=@��{�m&xU��0���u���J�1����s���vK�u�k����U�O�IE��hn�����i�O}r�aȹk�����Hۥ}���S�x"@s�V��"��M�Y�>UU��K5pO�n�	�m��k��=�������3R�2�8K�y �g�s����XPʔR����ǝ٦��;���$���fJ78<<7�e�oEX�15����q�]IH�w���X^�3z�H���?������R8���%��X�1f�(��Y����+���ɩ2��������p���	����K
��6?��������X�?��301�=��A��=Wr�Ich\�A�j}Fm����.���83�Ld�YP�y���hb���+#82�"���I�K;��n��V6��o�/��� ����	Υk�����Y�$���}V��R�i��i�<+��'�M�Yd��J����~��������e/F�S�H�In��5�p^�[�It	�uZ�!i_R���fl֘dCұ?�Lqd��E��$4��^I�/,N"Ԣ��f~�y\�;��@��O�����#�7�ı�d������@0�?Ƈ����Rs@�&\��m�b��^����Cb���m1y ��'��OA��?:��b���X�|�J 	�/�lN�)��`��ض�-h���fhJK�`�G/�3����X��S�>�Q�	(j�]OF��5��\�:^���~
�wC����F���pP� Ç������y�zkc	���~�D��\SG������O��r����#�s�ԑ��2�_�`�#+�F�����hwJ����`۰�""ZL&rf;9���~aL�W�Y|m����h��'��$�p����=;�\�OD�E��I��f�sS�6=1�
���M��$�!1#��'�{w�<��5�G�=O�kaUT��|��^\���%����-bF�ژ��{�fi|���j�v���&6�Lh�&�.���$VKė�8�6�o��:)-�y�3%�J@��Gh_�4��>m�#[h�qm����Ҫ�����3c�g
AVhj4��{c�aC��Cњ���HP J��Z-P?��a8<��Y����O��� ���A�ho���y)D��'�ܬO�&�����%ދ5j���μ�h�͞�#tTj�%d[�O�B@w'W̀?N����6x�SG����|���P�;[�Ѻl�X'wj�_�Z�>JKaȞ�%�]*�qh�48o\�f�{)f�B�N-�z�}�F��;b�s,��_��������jm�+�*�y��͗s�!���Y�L�W��7�/=�u�q���-<�Lz������[W�E�S�S�������q��c�?�G���y�c,��;�B�,��;ͱ-���~?��y�3�L�+;�~2�jks�z�+rL��?�SusM<9"�kbv�Q���$
�?�D
p7؝(/���m�a&��d��Vn�����r?��E�c��
e2�Ѧ�̩��nw��Baح��K�-�����d"FE�X�露��/7�k̤�8#����e.������rX@�������$�Rf�((oc.�ܡ�l)��E�n��(���4��
�m�t-f�S�R���� �z**��ي�*v�j:
5 �4&=Q���?��U�c񩪜հ����"!r��y��0ˀ�yݳI8��A��f7P\iYz�=�-�b�2=f�������U gE�c����5�Maġ&AD.�-	]��7���	!�e�28v-��$?�ތ4"p��s�8?{�Ag_�����mb�=L�}ʹG=i��j4��8ǃNq"�������Ǌ6�)��oՀ�+X�^W�Ӳ���7�Ay�H��z�9�J�H:��-�qTo�V��)*�L��p��:+7�]���)�Q��P9t4i ��!�~�{�V�,K<?��2B�D�ƨ��z�R�4�i�3�`��B�9���
N�]��r�(��ӟ���.��2l;t{j��i���p���Z�S�����; t��Qy�;�~���%�G�YF���z��]��ɥ�2�f؉���ڂ&T)�э݀ќéH�zV#�d����,�nǗ�>���,��xKn$�y�{��]�ǈD--1]�ʴ�SLr�!����d�+���6���fՖ|�s�؂���76�jUnf�e���
&�7uS����WiA�O�����S��-�UF��x�����_v[���ւ��/���I| ߓ�}KKKUK~�HϻoC��S�o��$)��l�b�<k��'0Q�MY����c��*�x�J$���K~��i���TR��yF��1���I��D�Qq!�9� ���{��$	gL<��zV4qp��/P�q��N
����~��vO�t����qE��U92�}a�և(E;'3���P;�b�~H�(r��c���'{����T���`-�aD��cY����neH�!�6��w��8n���CrV)�H�I����2���G���u�%�u��?)��w���G�u�04�v�/��u3��~~K�;^�%^q��1�ر��N���g�y \��$C2��T9���YS���i�p;2�A�SMY�Y�2j�=�v��'Q����� ��{���G�@��X��S�w��힥����I߱u���>�����m���3����Wڮ���l��ל|��Y_��-���g�h�;S�ż���5��5P���`�9��"��E�\f��������F�&N�H���fQ�t��<	.�N�v��]c�ٔwk�t�T=qA��5B"���"���C�?*i��AJ1�JRP�w�N��@��<5;��;��Դa��9W�2���0��~��:\����Ri1�P��a~W ?�� 6����21d������Sי%ȞaTS�<��J==�0$��������SAR�=��lADt�ғ;�#�OA�Ib=�`�):�DX������`q�+��Y;+{D+�8X�p3@V�Jm�e�� �":��R�����0��lǿ`�L�����4\h�7�x5�w��2~��Q�KG�ڊ�Sܾ��8�&��,M*֎"�u���h�@A>�p�h�_�K)1X��� �w��P)�n��5��6*�.�j|}�h�!���RR��@��q#��F/��.g��EV�r�)��� ��t}�EI[�6��!����9Rz�GO6��c��4F�m�����]�*ߌ�4�ʖ4�@'aq�md	(�c$'�D�r()����\�����Xt|��7nfF�\J't��J���Ѡ��Zu+9�$C���p���;-��C�m~��3e�]ʄI�Ȟ�Aʣ��&v���v����:�з�O�����cL����Ë�+��7<���^0 ¬���a��Rr��_�.o�廈q��� 9�@�ʱ��)����\������D,�3�C9�ò�%NF[x��sv�{����X����E��"��Qϭ��6�$`���J{�cR96�:�����b�J������A`��+��b�?��}
ɤ���X�T�����$1<���ǁ�^k锶X�ܨ�CZ��73�
nBh��,�	��a?;��mN^fD��W-�N�qj)	����-4�~D(�"wgr���Fؠ" 2���[�P�
��D�5)��	w����6�-r�K�XR^�4��pl����#ZU�3%�B��w�d���b�#!�g:���>>T��g4w�|]�z߂A���Ēh,'[�lv�w�/����xL؃K�w�h�pM"��m �Hf��`=���1G���%VaƇ�F�p.فDh*���f!(�T�l��k���t"�E&մ��t8h&�+���������5����10�у������Xv�<Q��F������H�����f^gn�׸��!�ݨEJ�
�P�I��i��q������K:��
��y�GM�(d�F^����c��G�v�O9Y��P�Rn+T�<5N��tC��i߉��,�d�du�����d��d�=� 
����v���[˾ecw�v ���H�����tWuUoX�:�W��gLO�&�M��֫>|B@n�;� q�5Ʋ�We&�~���.�r �H+�FdQ;�ҏ�"�2�K9N������"�X3���t(�?��5��h|��-<��2{9�R��M/�p�3b~ߜڌ���E4Ɗ��2CJ��r��,J�'!�����dM�U"�_G�p$Yv4�
Q�}488�1ƜKbjDS�Za�GΊ^,�&l��E�jR]?�Z�P_-؎m^���<��2������h�#�1�	��c���p>�"5/�ՠ#٤�Qj��U�yۭY��i�$�7l\��6�n�Ϩ��I��" ��F.����(3�@��W���zqϋ `I�b�cm�:I�"�Q��o|D���&b�i�K�J�n�o����"��+�)U��j-�\��z؉��W��z�9����c�H�!����wœ�<.�lN�)w+?=rD3̂1n�o+���
����\뚾[��4��@���#�Q���4|�=�\z,�� A���,9��jU�2I�0��VX_��_&��b�����9���O�^��a�g��Nv�j�u.(J���u7�CV��b�C�4�(��B�a��!�:��J�E��ZlN��G��T�O���y(s���<k u�ٞub�[�\C��iq5��|�6�Ⱥ��m(ģy�����3��no�8���^Ѵl�w(���Z�{`g��f��Bݐ	���51&
�h��xie-�R�4 ��������U��,��Gqח�`�A�?���Qa�a���n�WƲ��?�F���vv����	�R)��ى���#�.�!���I�
�9ݶ�|iI��N�Y,;���~����WxuTd-����:O���,п?�ǽ(�$%�+�ȢȁQjT������+�d��r(��wPX��F곻ѯ��0��E�,����`"���S�?ʱ����dw��щ��<)���|?����J�m��	��#��|@�}=����ͱ��\l�>Ns�:r��em�O�I�<�<c4����$@�6i@�N�'b��L�<H�<+ogc�jmLA�f��tGaSp�9�N��?y��n�Y`����s�V�|D�Ww�|���C�ެQ�r��e;m�J']��R���R��Î�ɕRᄉlE]�qF�<�i(����W�_�Ð�����!��\&f����{��v_9%��(��G���\P<Ӭ�FM��Cy����],��-H�+1$ߪ�M<L�FB���!r�G�CI�5AVhu^�ɏɠ![��q�����E,urEk��p/�y�5ؤ�ϼ.
~%'�dM�@�D���=���U����۸1֨�����cc	�S�#���)����27-���������<jH*��	�T,1_J�衊m���\�t{;f���M0܁ǕZ�N2�Cc����vi�[�ܧ����y?3p+���P[ �[��%�©z ݰ����iAEc�Z�?�=>b�l�y��'��1E�;��Uc�_�Q���ۼRj0:��i�!�u�Meh�sd򏦖������T��IIɡ�@�?o�D�)�xW-�o*���v/-q��w��$�����شv�s�3fe&|�NM��t�h��z�R�K�+n|J��
�G��5!�a��� E���펖)�[w�5Z�̖��J��9��W7��K�-�/�&[dy�SI���;�]8���_�	��	�x�>�U����ץy�h,o��!��d=����Pu��gS��{dW�h�+��O~�2nd�7K�5ߗ�\�n��ɨ�N����2w�h��������t�5�+H��.6��|��N�~Ǩ�2Ra����ۑX�J��B���U�UX��;�DUqQEg�F�)r����1cZ��)�*�&�4�Q}>��Э����R	����n7��Z>��Sʝ�L��q���F��y�M��Q�r��s�o��a�"�e���!��|˦ڼ���N×1��$��hv�?�L��k�����t�����:I#�>k�x�L��}dt_C��$,���\�.����"�P�Ҏ3g�!ֶ�Atb�/} /V�d�*���X�]
���å�6jn�o�����,�7^�\5��Ri��x��I;�	��!pT5u{�5�]�� K3�&��s?Ġo�&���tA+қ���ºS���sQp������c|D�6�\�Da#)�������q����M0@�ܶ��H�5x��aXB�S��	�SI���L��x�Y�D];�(���M�X�(GAGb,��^if�; p�i&��o�IcM n�`f�=D1�z�>S���m�BD����愾�wP���a���t1��c��Jku/:|��p�g[��ڊj�蝕7G��O����*�=�0���@@���	d�ln�n����lh�MQ�f���q.,؎0/L>	1�h �
��F����ϢU̐�1�	r�� N����q��O�h�@x�_�t+��2=�[�:�sO�y/��>.�
6Ot��R@?�JR�4��o-�g����e����΂��v4���m�fm7��{G���R���>&�I�P�M��#�"�ûV�a�^��P_�V��13����]'{'���[t��	ݳ� ��lۺi�-���F�P���ػ+�x\H��
G����thbt��V���Ze�2@�EgP����Q�1hoA���Z� �F��߁Qv�Mz�,�Fe�8������F)�XT����ڡ���I[ܩ��hg� �h_?
�:6��a5|C�.;U�yzDޢ�,��[0|��@� U�Y�_�s����Z���qPT#r[�Mk�ώ��;�f���W��8x�iP����DEr���Sl����� b�U��>�����f��L*�*I�c����QbH�*T��{[eoQy�X������F�8`��=�Mreh}�^�N��b�&��XZ���X�x�4aV������Mպ8)K��X(��5ߍ��/=VÈ�`��H4��/�N��b,��� �d��$��a������t��i��r�,���һ����ab��L5D��A���E������t��Ȯ�k<�w���)jQ�Z�AB��T���x�,
������SX�HN��X����7�a��>���� c������]��|Հ�A��"D�JJ��Yx����p����t5-U�>�r�q|��o\��p��"k��2l2&#���Ѷ�\�gA!�N�_%{��hU�X��a���p���T[�yE/n�����	�Wm��6�=�e$����M܁m��Y�lC}R�fb� v�@����C��p�28���E���2U���5�������
�ECF�Z-yv4��؈_G���أ���C�4Z�7=i�|{mLh#��]���Z�.9��@ޠc�Dv9�#Q�l�$�Vw�K@CGȈ�/G���1Zt�#[
�طlI�����)X�!\�ڧ[ۡD|��������t����#Í\9��9�9J���y\�����KdH{��+�*�F�����8��)�I{a�?�a�2Q����,�:z�<B�L����RiX}<ɕ��O�B��K����>��U��oJ�>���7�L
�/�)��p���a(�v ��x�V�f�q���VEO��Y�k�bQ��*k���]l�]-Z_��3H�����^�s��r��0�661J�܅:��ۭ�L������V,7i��	��h%W�7�jr�
0�8��>���� s
�]���B U�eHz�R\>��$�(���J�*
��L�vh�מ$O+GN�h������ǁ��e���*���e��$`Nx���D�˸�R��ZJ�m����Ɵ����NO4��Ǌ�p�<#/
�;RR�̱���
��9v�F��p!��k��P��T���iq�t�S���#MX�<D~*�B�j"b�g��g��;T��3�@��f��W�����S�"�s� ����!6J%I]![�g�<�����fnx�dn��I����<�k~�DΏ�<�Co,ع:��1eK�2�S�=�������ﱥ�������/��1B�-��Ks��������a�j��F����}��A�W����!M��X�����(���t~SèA���ښ�򊀎Q6��o��fH�X��S�����#��Yy�� �s�k�43��*���~ 
�wj{w�츒|es�L��K{�bR6"��p}2Ѫ�Ciܵ�S ���
�h�"n�yA�u��	�>�Lk�m��A�[W���mu'Q�4�\���o������o��Nf��+J��"1�%t��������*S-C�߸7F�{�GV"Wp��=xFep�{�j�݃���6`��b5n;��F A���f�p���ا�肔5-�uWS���nJ���m?X��Br%� ?�
a�A��[b���(G�F�}�5�=4+��YN�����g֋��#N�w�������kM{���Ne���>r���i�ia�I��[<�G���pzʦ��h&sU����u��{gN?��>r0�|N�ڋN�{1נ	�ܹ�!�l�MINpYZ�!J���;��J�6����n"��THn�|����!�Z�b��*؞i�Ө�#}<�\�j�tv����H���b���HsZ�+̖��8>������ڸ�6Rz��Z�
�����)'$�%d�vtK�n�U�9�-�h���Q����X�݅�l�%�#�{����P���/E����\h�����x}�ÜI)ƞaz4�D�_4{�����^�x��(Leݐ5�qC��KRs�yA&�aX	�-+��:��WR�� ���m.���b�(�Ҳ��kR8��(-w���F !A������YvhD*�L�ύ�ҙȳ��d�7��d�C�T#
9�WdzBX�Ί4<�I�ӓ���x=Q�dJ �pN7�"m۞`������E�s�2��B���3Ýi0>r�2���������A����i߯�Zs�	���8se���ގ&]����~���	�z�lc��s��$��\DK-?�q�t9BL�5���U��	�b>�vK~I��-�5�N��[������2g��2���ڿ�-����h���.m�D��a�]���F��*�����*q�̘�m��`�{'>CzjΫ�
bM�� Q��da/އ�v�����wr����Hs��1K���?T�����b*��Ŵsa.٢n�����2�Y�-�������Ca���?Ջm���/qݔQ+��_�.*�EZ��� �9�ߴ�5��E����=u�v��l>ka�K��H�_ܒ
��L��v�G��3��H��n�]����_��A�q��Y�z�6�m m���\5�l�s���gBH#���7�kXq��l$`&��_$�;|�N���P�
�o�W2��{��6^�H1z�}���@��:�*8]�{-?��2�$?�uP�Y�߸h���^�[��,��]���[q7xu�+�itH�����o���}m7ο�.��*){� �"Plͺ$pB-�pOl�"w׸��`�#:�_f�}FPpoQ���ߊ���~�4�\��`7�}[h�4@YIܬS��&�c�Ч�ӸX���IԚFY� C�|�ɑB��N9Vƞ ��6	��M�˜�żbRĨm9ۚ�Dyk#%Bԛ,_�О�����	Qp�!����55*f��J��R���U����(gA]�T��x�M,�ȩ��1�|���@��39X�VM�Q�E�0�����$O~���~��^�������'��q6'(�<e�zl	�朤�m%Q$T����?�n��c�Y���ᅢ\��)p�����3�3�Q|��l~�܊�;)"~JzOV'?�d��>ytH�;�k(MwF�6�l�^�FJ�9��|4�qG��igM��gM����1�>S� w8��}C��q�2eֵx�
�2p��:��h�kC$ ]��x-s�^"\UF:�£����*��ǮRP���g�yүz��^$�z5�P_>
�w�D�������sCIˮ��еF��f�S��^Wj6�К|�sf�R�{#�>܍���Y�v.{��2dg��6��ҿ�LK+l�jg#��<�ʔ�B��y3��$�����O]�����ss:m<&T�vIpxa&�$ n����&��n��ch&��-W�Z�@��;\B���_U1` ��;�n�8�<NM���L�c�7�0Ǵ�F���=���� 3������-;Vԟ��X���\���۪X��*¼F��j�;~$�ÆF/���g�|���rh$�_��֍�Խ�9Kk^b,�Wɰ�g|j�m�#�O|i!esK�I(k7��E�}�(�l����^����"��-=bW�2*�"��s辺�*�A?�Y�P���*��?��������f���F�6m=��;}Z����<�3�\�%D
Y�_�ԉZz�k�U�����j��ݑ��ފ�����׮X�=g��E(��R�Jp 9z�w3��x3�ŎV�B�o^u[AI1u�r�m�g�%n&|�������k�}�G�/��M<V�][qk�S�߇�f'�eCb�p�͝�X��UVB#��OUNu����~0�`� Ӄ�J��6�8^:��,��K�|~B����۴�l�Si���{#�]aeQ��N��"����}K��{Y�L���Jb8�c��q�5�T�Ī��)	���7�h��D�j�$���A--.w�x��G֥nr
ЃOoS_�-���e�[�t�ׂ��[�/�1-�^}Z���I����a��TmϦm)j/]���f���֫Y����xA�y���9�1Ke'}��(��m����9R*�2,2�u�W�x��2��V<JN�����øE�����GPA�D$�pn,��qS�tjmL�t�p�'�#E�No��_�=D>�g�˴�����ڱ�qy�,�j���KM���j��םKgD�����W�2K��.���R���=zw����&�H͝�z��J���f"����kC�g(�Jh��	oCy#:��o����g�a�P{�
?����&ep��J%'O� �_+�����υ�xRD��4"}[)��_��l
o�y�e4��2rzf&�?�mr�"$ǩl?�`�$��;!9��������O{"�҂k�8�A��R)�� �D��%r��ǡ������#��4��p���Apo:LHϐ9�

�K����Q��fO�&��&^ ٷ�vQ�#MϦN��TO��0ar�^R2�����<;�v�_��c��ʚ?���Zq5���5*Eb����%�#R?�N��K�H�2bQ�taeX/7�+��Lsg���V����1�T�}�NE�������xl���������^�}f�������!�sף%z��֨�p/�D����>����$R�L/�-�����g�����ᵥ���;���3R�G�O}_�ch�%�;�r��!�o��P��+�XO+%�Bu��sM�Ł�p��(?*W�jGfA#d�����#}]��1o_�o����]�j�|)�CPe�|95��	-O'��1�YAҠgf��Mp��������{�~�1�o��4�/��tzcds)� �����7��g��[���+�6�N�yC�o:4�gBK���@��S_Ah$��{�ez�;��ǫu��&O�l�Ą&�T�ף$0/!+�z�F5��{���6q���0�|��9���&F'|���/&�s�j|/��\/M��@�|�x��@6)S,�S�A�)�+�D������Я�3����C�eM����i]=�L���y|o�T���p�^Ó��s��+ʱ�X��uo]v�δ���x���T<��s��8Ȳ�����;�0��hY#����vO� ,�dK^�W�o
,��[�V��D�`䞤Q#:��#(!a,	��!:P�i��gwწd,��� E�Of��x
4+�����薽N�6��v-���aWO�ǟ�a����6,\f{Q�J��63��W��;Ĥ�����B�\�_E�0 q�~����xh|[�����1�EϺ�)����D������Y^�	�ڢ�hM�K����/5f t�f�E=]�t�O�%��l;��N��2����z�<JKFD�g`t~D^�_C�?r���Su��Ү�U߰C� �µ��ȑ�O�i���袜��U�i�����]�B�� �9�/-�:7rE+)GA��9f~����1߭=�} 3����-%�r���@2N�6�Q�q�y�06���%8�q�%)�[��uQ��Nb�uR�#���v_�\2�܅��W=��kfͧ���u�+��-�S�R�~R�@�w�����'�*����jV�����')���ի���}��;4|�sn�T�>]\���\F]<$F"��~���V�O�ݚ��U��洲;d�y�ړ_���!S���a�gq11�Z�(>>5"�9�^�@�WSs�/�ǭ[�gB[�&�\�����4����ޟ��2wq�@���	��O��癬������C�,�t����"�l"���X�I�W�.��dML{i��8"c� ���)��\�LYqn#�V����>�Z���L_u��"j�2���n��s�ǝ��@�Fxj��:C����7l#��`4�ņeN�I3�C���6�\���%�s��N�Wy%��#�@o���i�L�p���/��y��x&�nAr���B�e:�-��,���7���n�a���DF�,QtI�O�r��^�ȐW�B,����T��g��w!�W5�������p�/�U���va@)�oL�u��4�V�f~:�Xe1�(uv�p��kl�x�������-s�d�d�E�̈́��=��]oGZ3�l�L%�޾,������q�^,�*iV���4�4��J-\	J�F��r��r� ȭѩ�a(�aێc�Vٲa�O_R<	�L�� ��<�)���׎|�e�v���AiN�g|0d��X>5B�Piϣf�[i���phI�E�k;��:f�WҾ@Y��i!�a�1Po4�x}���A8T#�6�����f0Jʁ��������9�qX�n���R�U���WӨ$��@k� el�&�K���.r��ČhE~5���Ը�,���P��4���Pׄ�я���J���j�`�Y��W`�'���s�~[�r/|����a)�Gޛ��R��f�>!�ס��|~q���~B[���E�P�ŏY��P���S�	�h�=������ӯ�h�$	r�5�I���g���iWM� �W� �x�'νm��^%���`Ɍ���b{��"jP�?w��֬Ƀ4te	��AҾ<T�/�ힻ��D�`,'w�v*ƀ���جqEM	�$�su��k!D�ˏ�KUL�r!igA��x�A��E���N�ɳr��	;4T�̼�;���������^���=�R$��i�'�j��/2�9�)k3C-{)V���ɬ{�
�_�*	�K(}����l++�tN�7�s]�"��T��6x*W�m��2&n	����z˸<3F����X[fbFZ.�uaqt��.��h9%�� 6�~�b;�7�9Oy���0Ǣt0y?N�g���4'}U��Im;�Ț��F���(-v-�Ɯ"��rz�>�9���)��]bL]�6[��Ϙ<j�#@+���+�L��c>��<��
`���(����z��f, }��LR	ᢇ)��j�26�����n�
�`fJ�����2»p�	�����16��m�UI��EIo)��3[�����=��l���tw��ęMOY����y�?Vt©���Rɏ���G������ƨ&Û�,-q��hjg�l��/N�x� QRg�\�A�A�
Ӗʇz'	����N��3
��Viaϰ��DJA���E��;�v��uy�<ʊ���2�=ʍmZ�'�9�M(;����,ыҸ��|kx�|MV%�O\�EK�"l,-�D ���']�@*Q�'���H�c�LK�y����0
oF� �+�ˬ��}T#���JD�\^�����7�^������/��¡)���[ܪ��4���b�^lFpCW����ï_el�}{L=��;��Whm�ʖ�f&��~v������(P/�Ā���Y�����Q]h1B�1|��6	qF(h��r�x�Vu���ݯ՛ǋ�hI
!ı�g߅���h�#���j
M��ټ��>q�Z����ܠ�b����p���Q>ď��3 L���Rt�~yp��bX��N���F!$�E'�����1m���1��]�/ ӕY�]�~i�I�A� ��r9�O3��7'����W^X��x�NW���k�uX�l��IC����X��d��	��A����׬xn���L�g�֚��7�WSob(nm���9��,���:T��_�Y1��2=WpZ�7]Z�'�!���������Jm-�j�����`�BV���.5�)QaJʦC].2����بiĕ�AK��Tl� S��}�;�RT�����l�UJʻ��W
-���J��}�3[R�9O�˶U�1�[�e��_ aZ��wf�������.J_�36������{�Y���Ԧ��Fv��V�p-\Y�%�d1ޞQ��=&��ܮ㛷���~,����^��G�Do�£��.U�(E����|4��z�N9g�_�%{���S�ַ[��!V}��N�k㝌z�n�L�(A2$b]�����fa�vwB�K�=;��r�a�q=���ڃ;��� �q�X�/�!㻮���v��&by�V������M,�c�A�c�z�s;��%j�f�}�[��xގ�~���},�jq�^[Xc�����M��~m��O���2)lB�iTC����h�d�c�s��}P|� ��$A�鞘	3�|(������6(P!��B���	�Z�����"�9F^o1]��x�6t�{�49Vdr:��0�9��	�?�=�q���`z,�y;</M�6�m��ʘ�*�\P�w^>�[�So�) ����s����@F<�?}��m��'���ߖ����3[E�]��'7ݯ0Ǳ~-��?�.�@<�=,!� &�v����G�.^^��ø�S�8y�ni�z7漐:���^��n���ڇ�^K.ۡ�o pE ��w(h&�8��a�k��u��~L-��9���b5#yu4Wk�{V9K��?�3�Sދ�.ӝ;���-+/��^�m���q�-u!�*o�r��Ԧ�|��T��l�nЖu$��υ���|��:R_,Z�8�NA�|����p�(;d�
�	=f��V�o
�@T�Q�2�]2F�K]����^�o���)4��s�8=(
٤���:l?UUi���ռ�.7$9�u��1eR�kS\�#g.I�>�b`�C�x�|ۥ�i����i��Y�Q0���,�I�M��/u�
=�Rբު�ȡ�K]�����<� S�T�p^:/iJ�8�&kbs��4���}�.6�lӦE�$����q�
8rz���r��w�/$�,9K߭s�q #H���@�-��&� �oc��Q�]F
f���#�=L}�4%��?�<aLц���
|Rd��#�1�w�XQҽ�'�ZG�.�uTݹ(j:&蜆��gmQ<LM��rj�V�.�]���f�)#y���B�֘��Է�XS����w:U���1��l���sůK%��=nx����{1^'��z˟�l`~z��~d�N�5��x��Vw�����CqW��*��x��0ng�&��*#m�M�s���P�J�[p�'c&����>���_����7�.�T��8��V�8\�%
~d�xW>�}��S�.��sn���m��wm��9�&����9�E�˽v���Q�q��K=�����>j?����6X�J���Z.�@7̤�PP��O����������ܼj6�(A5�H&RV�U�	Ȉ�G6�@�P��]����4>y��/��9���n�K>���K�V�"�'|�@��]��6�W�`�i���xy�wo�6�2�<���Iٺ?�
6'�������J�~�c8/��j>�/f���R�""�ַ*���[���@��3mQCH�2�٠�����0&�F�ڙ6��鈃�h�А���|Y�.2�Hi�Hw[�Rl���M\����3���k�mv��-��#c2�_40X�)i�ߛ�D�$%��5��ʉ(G���i��A;el0�6�Y�԰�6��i���3�'p�̊�r�4�aZϰ��㗓q�J5��ίa�����5� Y
�y��:�q�� 3 �F�f������fAHjq䑮��>��񺮰_��d�ĕy�3(�m���e�;��¢Qlid�l�A�B�=�	���7�^���y�-R��-�iP����Z)��I�kF[��-ƨ�%����O�K�`��M��-fӋz{��	���z�[z��#�v2?Rԯ� ,���g�'2ɟg��W�S��E��̚ޖ����{3Sa3�Y�ZQ���4�A�M+-��ϫ�#�<g�ht�c����1��-?�zw�[�/��;���|\A&�`��Y��1��u�~���~�S	�놡 Q�C����93+a���/��֦52MP;�Yq4�]�	�^ ���-�a�vU�B�-nm��;���I-8���1j�3�엃��+�5�y�\�s'A'�r��b�9�r�X���<��d�맼�ु�B��q9�Yc��_���U�o��)���R�L�<Բ�r#��C��O澖w��kH=1g�.��ج!I���T^��z����^Q��%��=k��>pi�)!���n֎�I��^��q�M��)���A�#d��s8��XL_ ����]�Ů\B�a�ҿv���wT_`�#�A�LTRq-bA�9K'|�Pd���03)=�7 �d��eJ�&���uA^g�ܷ"�%�^�� ��eˆ#.�^/�L{���`1P�  h����4��*��2�{�J��p��he����æh�|���Ĥe�h��R[�4W,��ݮ�3�JQ@蹷ɩ%���B!*��>�]��|� j篾��^�)��+KS^%۸B���x�-�v��q��|� �x�V�}
첽�"�yB�����h:�:�5"���cF�_��K>\�^��Ȍ<�;u�3��2:)��Y
v���S�2Dv�u�U}Tn�M������������LOѓi��x
k�̹�c�sRNX$��Mpt���ׄ^i����"�x��H���T)�#ˁG ��ŋ�Mo��"<j_�".�&�� �#�e�oJ���"$� �Ԋ�g�ǣk/����C���$^,����:P�o�_�FDBrI���*;��������\���.�@%��N�ȓ�<�c֍}:'ږ����D�0��)����I��(������uB�H��UM���	�J�8�}���,���V�q�nH�g��5�ʅn��o��u����rnlG�Aͬ(�q��G4;�����f����U# �^��HV9�����HF���MvR���'�Pmx5���Bu"�������=<�:r����)���K�`/1�jQ���H�����/���P��ě����"���x�ƕ|�t�c4*�x��_���(����%e�w�[n�e·�
9��jL��6�	:��� ˀ��0˺�p�X|H�:�a���!�p�&�5�-=�qu��	T��������u�xS���s�v�����;��i���w������J���J? B��t�K��96��ek�VM��˥�PX�|� �V��V�|�E��]�µ�\N��@ˣ�F�AE������P�P���b�*ٕ��8z��
s������]����Ҏ]��:׍��C�IL��9��p�h#b����	���'�,"e�7����\~B�W��t�y�ss�k�::�b�9�i�����1�ѤA8��R4���p���
^j�F�P�k�����`���������K��u5�:��D9�h�L��e���xc�g �$z���@�bvm�!Z�V��#W�ϴ&�swiAc��|�)��j���m�$;Y�����`˪���s�q2$���{?�sㄉ΂Ȩ� ��NQ/i�N�	�ER�b�����4
���t�KR)KB��s����� ?ST��&P�-,�vfmӸ��he�G��Ce2�l�=/�#S-��,��5��R�<I I�
\w�t	���$HJ?�����#���A9�����~G>���+ ����/��.R��@��j֖�_`�T7�Y[�X��>ih�*���e�HPH��/v�b�ѥ���1�ϡA=��)��pv�D2��w���0��{��e�|%��NF~�;�k�7H��\�?w�.��{yOy`� ����Zb،��3�3�����]�I�,�������<.ַ���V��n��_1�U%^���*�[N���.�_����^�?��g%�*��	��\+ZN>*�B(�U�I<��`量�I��@�x���1e�5��Z��*���п��|����� DO�$�oॼ�|�	~�b��Atb��q.͟����9� X���'0B2�Ӵ�	��eϼǇ=˄��uvcUE���r-~�uP2(�/T�a�Q�A�UN�X�#��I�jڛ�=���J1��D��/*_�u��8~G(u*�����:M�u�N�@GY�a��,(�6z�]�pre݄��Rh�JWT��蔽g�h�'�Kl��;CD+jʋ�����I~y�
T0r=L�������B�;hJ6(���a3jKI��a�Xs+�vz٥��L�0����[Ȁ!ᝩmV��o-���З_�}=�����Ш�r�������
;��j���ͱ�ۜ�⚥Ê�ɿ�S0�T����E!�~L�0!���D����8��u�p�5*{����")X:A���{Kue��ط9�j��w���!.�k�S`��kg��n�C���?gC��EKJD<��l�Kj���^�O�H�ތ��XU��0�L��4?$��[8@���T|,2%���|~��� ��rAt�us� ��4u|��TZ�$jyZ	*k/��ɵ괌qNܛ�]��杯�c�g8�Ү�Y�z��~`7�������h���K>}�rł����H	�G�"�^.��ǁ�z��"��46S�IB_�T�ސ��Jı�y���GЂ�����M����EX��cIu��z���|f"�o���|\���!�����Ĉ�§k���E����67p�BȸsvWs��B-�����u7����!�Eԅ7b���%��2iA0�S���ݳ�KG=p�CZSQ���OǄ��j@t�{ �eM�`�����/�����@�n�`�~����]ʥ�Hr�:�ٞ�)1�5۳Oϸ�,��8!��Eu	|�S�B@�
P�	��,��m�%��x�;�:>�����b�ĩ���<�&�R�����1���c�>ٛvV �Ħ����=���#"F�+��l���"��������V���/��2�<���=|��/��������c�R2�n��?��x��4�>DF��'�S,ѯ�6YP?�7G�)gDJ�Q��%
�������oy�1D��5/��x�A9r׽'J�a~������Pw�4M#3D:=:
���� \!�1��q�A�ȴT >ɐt�5�����}�>k����J��5���}��� ��z����<{K=����-��R`��k���ag����oO3�2�V����Ӡ�+~:]�������Zϕ3��_�.%BeTV���dcMc93�ڪ�e*�De��Q2-��:9�4���r��VG�y&�Y���(���kFN���/L��d�����s����h�M���x۬��ؑ,�g&��F�~N/4�-�h@�{��~� qL+^t�&w�P��6N;���
o�����
�=ZO�%w�������HO.��%�S��/��-��P���Z�/O5�+�>�5�K;�.�a�5�x���ɓTk 3dG�xcIY��3�Bv�������Ck�Mf�J�t�n(����9�h�O�/td�@������Q��z�Yc��2�7��S�v�0��g���;A��e� %T.����3�'Vľ��_�uM��"��L��P��0�^��?<��zJE�5��[.z�?� ���1ܑ������j���#�4J�ާ�&L�~dd��u�@Ƃ�,C�B��