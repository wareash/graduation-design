-- filter_50_1_4_GN.vhd

-- Generated using ACDS version 11.1 173 at 2014.05.16.13:43:04

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity filter_50_1_4_GN is
	port (
		Input  : in  std_logic_vector(7 downto 0) := (others => '0'); --  Input.wire
		Output : out std_logic_vector(7 downto 0);                    -- Output.wire
		Clock  : in  std_logic                    := '0';             --  Clock.clk
		aclr   : in  std_logic                    := '0'              --       .reset_n
	);
end entity filter_50_1_4_GN;

architecture rtl of filter_50_1_4_GN is
	component alt_dspbuilder_clock_GNF343OQUJ is
		port (
			aclr      : in  std_logic := 'X'; -- reset
			aclr_n    : in  std_logic := 'X'; -- reset_n
			aclr_out  : out std_logic;        -- reset
			clock     : in  std_logic := 'X'; -- clk
			clock_out : out std_logic         -- clk
		);
	end component alt_dspbuilder_clock_GNF343OQUJ;

	component alt_dspbuilder_shifttaps_GNLZ4R7UC4 is
		generic (
			WIDTH                   : positive := 8;
			NOTAPS                  : positive := 4;
			TAPDISTANCE             : natural  := 1;
			USE_SHIFTOUT            : string   := "false";
			USE_DEDICATED_CIRCUITRY : string   := "false";
			RAMTYPE                 : string   := "AUTO"
		);
		port (
			clock    : in  std_logic                    := 'X';             -- clk
			aclr     : in  std_logic                    := 'X';             -- reset
			input    : in  std_logic_vector(7 downto 0) := (others => 'X'); -- wire
			shiftout : out std_logic_vector(7 downto 0);                    -- wire
			sclr     : in  std_logic                    := 'X';             -- wire
			ena      : in  std_logic                    := 'X';             -- wire
			t0       : out std_logic_vector(7 downto 0);                    -- wire
			t1       : out std_logic_vector(7 downto 0);                    -- wire
			t2       : out std_logic_vector(7 downto 0);                    -- wire
			t3       : out std_logic_vector(7 downto 0);                    -- wire
			t4       : out std_logic_vector(7 downto 0);                    -- wire
			t5       : out std_logic_vector(7 downto 0);                    -- wire
			t6       : out std_logic_vector(7 downto 0);                    -- wire
			t7       : out std_logic_vector(7 downto 0);                    -- wire
			t8       : out std_logic_vector(7 downto 0);                    -- wire
			t9       : out std_logic_vector(7 downto 0);                    -- wire
			t10      : out std_logic_vector(7 downto 0);                    -- wire
			t11      : out std_logic_vector(7 downto 0);                    -- wire
			t12      : out std_logic_vector(7 downto 0);                    -- wire
			t13      : out std_logic_vector(7 downto 0);                    -- wire
			t14      : out std_logic_vector(7 downto 0);                    -- wire
			t15      : out std_logic_vector(7 downto 0);                    -- wire
			t16      : out std_logic_vector(7 downto 0);                    -- wire
			t17      : out std_logic_vector(7 downto 0);                    -- wire
			t18      : out std_logic_vector(7 downto 0);                    -- wire
			t19      : out std_logic_vector(7 downto 0)                     -- wire
		);
	end component alt_dspbuilder_shifttaps_GNLZ4R7UC4;

	component alt_dspbuilder_gnd_GN is
		port (
			output : out std_logic   -- wire
		);
	end component alt_dspbuilder_gnd_GN;

	component alt_dspbuilder_vcc_GN is
		port (
			output : out std_logic   -- wire
		);
	end component alt_dspbuilder_vcc_GN;

	component alt_dspbuilder_port_GNA5S4SQDN is
		port (
			input  : in  std_logic_vector(7 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(7 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNA5S4SQDN;

	component filter_50_1_4_GN_filter_50_1_4_Subsystem is
		port (
			In15  : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- wire
			In7   : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- wire
			In16  : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- wire
			In5   : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- wire
			In4   : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- wire
			In13  : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- wire
			Clock : in  std_logic                     := 'X';             -- clk
			aclr  : in  std_logic                     := 'X';             -- reset
			In2   : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- wire
			In11  : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- wire
			In14  : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- wire
			In17  : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- wire
			In12  : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- wire
			In1   : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- wire
			In9   : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- wire
			In20  : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- wire
			In3   : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- wire
			In18  : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- wire
			In8   : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- wire
			In10  : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- wire
			In6   : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- wire
			In19  : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- wire
			Out1  : out std_logic_vector(36 downto 0)                     -- wire
		);
	end component filter_50_1_4_GN_filter_50_1_4_Subsystem;

	component alt_dspbuilder_cast_GNYXW7SHLD is
		generic (
			saturate : natural := 0;
			round    : natural := 0
		);
		port (
			input  : in  std_logic_vector(17 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(7 downto 0)                      -- wire
		);
	end component alt_dspbuilder_cast_GNYXW7SHLD;

	component alt_dspbuilder_cast_GNRCC4IV32 is
		generic (
			saturate : natural := 0;
			round    : natural := 0
		);
		port (
			input  : in  std_logic_vector(36 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(17 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNRCC4IV32;

	signal shift_tapssclrgnd_output_wire       : std_logic;                     -- Shift_TapssclrGND:output -> Shift_Taps:sclr
	signal shift_tapsenavcc_output_wire        : std_logic;                     -- Shift_TapsenaVCC:output -> Shift_Taps:ena
	signal bus_conversion_output_wire          : std_logic_vector(7 downto 0);  -- Bus_Conversion:output -> Output_0:input
	signal input_0_output_wire                 : std_logic_vector(7 downto 0);  -- Input_0:output -> Shift_Taps:input
	signal shift_taps_t0_wire                  : std_logic_vector(7 downto 0);  -- Shift_Taps:t0 -> filter_50_1_4_Subsystem_0:In1
	signal shift_taps_t1_wire                  : std_logic_vector(7 downto 0);  -- Shift_Taps:t1 -> filter_50_1_4_Subsystem_0:In2
	signal shift_taps_t2_wire                  : std_logic_vector(7 downto 0);  -- Shift_Taps:t2 -> filter_50_1_4_Subsystem_0:In3
	signal shift_taps_t3_wire                  : std_logic_vector(7 downto 0);  -- Shift_Taps:t3 -> filter_50_1_4_Subsystem_0:In4
	signal shift_taps_t4_wire                  : std_logic_vector(7 downto 0);  -- Shift_Taps:t4 -> filter_50_1_4_Subsystem_0:In5
	signal shift_taps_t5_wire                  : std_logic_vector(7 downto 0);  -- Shift_Taps:t5 -> filter_50_1_4_Subsystem_0:In6
	signal shift_taps_t6_wire                  : std_logic_vector(7 downto 0);  -- Shift_Taps:t6 -> filter_50_1_4_Subsystem_0:In7
	signal shift_taps_t7_wire                  : std_logic_vector(7 downto 0);  -- Shift_Taps:t7 -> filter_50_1_4_Subsystem_0:In8
	signal shift_taps_t8_wire                  : std_logic_vector(7 downto 0);  -- Shift_Taps:t8 -> filter_50_1_4_Subsystem_0:In9
	signal shift_taps_t9_wire                  : std_logic_vector(7 downto 0);  -- Shift_Taps:t9 -> filter_50_1_4_Subsystem_0:In10
	signal shift_taps_t10_wire                 : std_logic_vector(7 downto 0);  -- Shift_Taps:t10 -> filter_50_1_4_Subsystem_0:In11
	signal shift_taps_t11_wire                 : std_logic_vector(7 downto 0);  -- Shift_Taps:t11 -> filter_50_1_4_Subsystem_0:In12
	signal shift_taps_t12_wire                 : std_logic_vector(7 downto 0);  -- Shift_Taps:t12 -> filter_50_1_4_Subsystem_0:In13
	signal shift_taps_t13_wire                 : std_logic_vector(7 downto 0);  -- Shift_Taps:t13 -> filter_50_1_4_Subsystem_0:In14
	signal shift_taps_t14_wire                 : std_logic_vector(7 downto 0);  -- Shift_Taps:t14 -> filter_50_1_4_Subsystem_0:In15
	signal shift_taps_t15_wire                 : std_logic_vector(7 downto 0);  -- Shift_Taps:t15 -> filter_50_1_4_Subsystem_0:In16
	signal shift_taps_t16_wire                 : std_logic_vector(7 downto 0);  -- Shift_Taps:t16 -> filter_50_1_4_Subsystem_0:In17
	signal shift_taps_t17_wire                 : std_logic_vector(7 downto 0);  -- Shift_Taps:t17 -> filter_50_1_4_Subsystem_0:In18
	signal shift_taps_t18_wire                 : std_logic_vector(7 downto 0);  -- Shift_Taps:t18 -> filter_50_1_4_Subsystem_0:In19
	signal shift_taps_t19_wire                 : std_logic_vector(7 downto 0);  -- Shift_Taps:t19 -> filter_50_1_4_Subsystem_0:In20
	signal filter_50_1_4_subsystem_0_out1_wire : std_logic_vector(36 downto 0); -- filter_50_1_4_Subsystem_0:Out1 -> cast20:input
	signal cast20_output_wire                  : std_logic_vector(17 downto 0); -- cast20:output -> Bus_Conversion:input
	signal clock_0_clock_output_reset          : std_logic;                     -- Clock_0:aclr_out -> [Shift_Taps:aclr, filter_50_1_4_Subsystem_0:aclr]
	signal clock_0_clock_output_clk            : std_logic;                     -- Clock_0:clock_out -> [Shift_Taps:clock, filter_50_1_4_Subsystem_0:Clock]

begin

	clock_0 : component alt_dspbuilder_clock_GNF343OQUJ
		port map (
			clock_out => clock_0_clock_output_clk,   -- clock_output.clk
			aclr_out  => clock_0_clock_output_reset, --             .reset
			clock     => Clock,                      --        clock.clk
			aclr_n    => aclr                        --             .reset_n
		);

	shift_taps : component alt_dspbuilder_shifttaps_GNLZ4R7UC4
		generic map (
			WIDTH                   => 8,
			NOTAPS                  => 20,
			TAPDISTANCE             => 1,
			USE_SHIFTOUT            => "false",
			USE_DEDICATED_CIRCUITRY => "false",
			RAMTYPE                 => "AUTO"
		)
		port map (
			clock    => clock_0_clock_output_clk,      -- clock_aclr.clk
			aclr     => clock_0_clock_output_reset,    --           .reset
			input    => input_0_output_wire,           --      input.wire
			shiftout => open,                          --   shiftout.wire
			sclr     => shift_tapssclrgnd_output_wire, --       sclr.wire
			ena      => shift_tapsenavcc_output_wire,  --        ena.wire
			t0       => shift_taps_t0_wire,            --         t0.wire
			t1       => shift_taps_t1_wire,            --         t1.wire
			t2       => shift_taps_t2_wire,            --         t2.wire
			t3       => shift_taps_t3_wire,            --         t3.wire
			t4       => shift_taps_t4_wire,            --         t4.wire
			t5       => shift_taps_t5_wire,            --         t5.wire
			t6       => shift_taps_t6_wire,            --         t6.wire
			t7       => shift_taps_t7_wire,            --         t7.wire
			t8       => shift_taps_t8_wire,            --         t8.wire
			t9       => shift_taps_t9_wire,            --         t9.wire
			t10      => shift_taps_t10_wire,           --        t10.wire
			t11      => shift_taps_t11_wire,           --        t11.wire
			t12      => shift_taps_t12_wire,           --        t12.wire
			t13      => shift_taps_t13_wire,           --        t13.wire
			t14      => shift_taps_t14_wire,           --        t14.wire
			t15      => shift_taps_t15_wire,           --        t15.wire
			t16      => shift_taps_t16_wire,           --        t16.wire
			t17      => shift_taps_t17_wire,           --        t17.wire
			t18      => shift_taps_t18_wire,           --        t18.wire
			t19      => shift_taps_t19_wire            --        t19.wire
		);

	shift_tapssclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => shift_tapssclrgnd_output_wire  -- output.wire
		);

	shift_tapsenavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => shift_tapsenavcc_output_wire  -- output.wire
		);

	input_0 : component alt_dspbuilder_port_GNA5S4SQDN
		port map (
			input  => Input,               --  input.wire
			output => input_0_output_wire  -- output.wire
		);

	filter_50_1_4_subsystem_0 : component filter_50_1_4_GN_filter_50_1_4_Subsystem
		port map (
			In15  => shift_taps_t14_wire,                 --  In15.wire
			In7   => shift_taps_t6_wire,                  --   In7.wire
			In16  => shift_taps_t15_wire,                 --  In16.wire
			In5   => shift_taps_t4_wire,                  --   In5.wire
			In4   => shift_taps_t3_wire,                  --   In4.wire
			In13  => shift_taps_t12_wire,                 --  In13.wire
			Clock => clock_0_clock_output_clk,            -- Clock.clk
			aclr  => clock_0_clock_output_reset,          --      .reset
			In2   => shift_taps_t1_wire,                  --   In2.wire
			In11  => shift_taps_t10_wire,                 --  In11.wire
			In14  => shift_taps_t13_wire,                 --  In14.wire
			In17  => shift_taps_t16_wire,                 --  In17.wire
			In12  => shift_taps_t11_wire,                 --  In12.wire
			In1   => shift_taps_t0_wire,                  --   In1.wire
			In9   => shift_taps_t8_wire,                  --   In9.wire
			In20  => shift_taps_t19_wire,                 --  In20.wire
			In3   => shift_taps_t2_wire,                  --   In3.wire
			In18  => shift_taps_t17_wire,                 --  In18.wire
			In8   => shift_taps_t7_wire,                  --   In8.wire
			In10  => shift_taps_t9_wire,                  --  In10.wire
			In6   => shift_taps_t5_wire,                  --   In6.wire
			In19  => shift_taps_t18_wire,                 --  In19.wire
			Out1  => filter_50_1_4_subsystem_0_out1_wire  --  Out1.wire
		);

	bus_conversion : component alt_dspbuilder_cast_GNYXW7SHLD
		generic map (
			saturate => 0,
			round    => 0
		)
		port map (
			input  => cast20_output_wire,         --  input.wire
			output => bus_conversion_output_wire  -- output.wire
		);

	output_0 : component alt_dspbuilder_port_GNA5S4SQDN
		port map (
			input  => bus_conversion_output_wire, --  input.wire
			output => Output                      -- output.wire
		);

	cast20 : component alt_dspbuilder_cast_GNRCC4IV32
		generic map (
			saturate => 0,
			round    => 0
		)
		port map (
			input  => filter_50_1_4_subsystem_0_out1_wire, --  input.wire
			output => cast20_output_wire                   -- output.wire
		);

end architecture rtl; -- of filter_50_1_4_GN
