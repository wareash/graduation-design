��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e����d���f{��@����S��>���4{��ת�AO�Q{���X��F}|6��ϜׇL�O'�~��E�ʆ����΀�����I�+N��~�2����(�Ϝ*��BM2h�_�Lu��'�ɉkT����R�h^�d�+i�]�A��a�ڀ��2NN�ҽʦ�ț�n`���p�@�F Պ3΢��m+VD�Ψ���V�'��ތ<2:��.�wm�ղ��I/�� P�gF�[�9����������ig��4;:5KL1D>[�=f����u!����Yh��ex"LR�9,Ea]&�H�oE���>�H�S&M~�]��T�=�Yy�G9H�'f�TO���m���Bz<Z)n�͎����¶���c!Y�]�d��s��|N6Ճ4~Z)�Ap1���ի�� ��@���E��!�'Py+�N?���_M����TO�(ڛ�+H�`hX)���2m�3�:SSH|=��T1 �,R���is?W/�L��S\y��qR�B���[Gg��|��Bb�$��v�YA��A�v��gF<Qsq��^���r��tO(�e*��I\�Ĉ�//C�0v�4h��D�Q)�3=-�}��X��,}%Zқ����m�G�DX�s����W��e�L��ᨲ�2����eԻ^��^A�|Y�Xѩ ���
�����A:?�9�x���\���{�����+LbBU�����h�ӆ2gi�'4��%R�%Y��P��Ϝ�ܠ�a��~��qD���U�ȦD��@�_�b���Q�Y��N�郏�1���N��	Eo$��#��|�cN��:�þ�h(�}F��oߢ#���l�sD����z
%��r<n�(��[���^'�Pvn0��s?i��9m��d��v_��Q���m�+���y�3'��#4�+'#�b�Lt^uB?[�]�����hQރ'L��tͤ�1��_\�h7i��5���P��'gה����[��A:���:�I�-��� D����
����S�*���T\Ej9O�n[M�e�Ě��%�	n�%\*'w<^��~1� �g&�>mL �njB�蓫{Y(������Ax��%�0n쒻��S� �rn.���T�D�������x��ilE�\�Hfx� 1I��T	c�����'re�o�#��ZS8�B1Y�r��%�\� 9]^,^� ��m��/Eaߡ���pz]=X0	�>;���z��7��wZ�a�C�d=^��¢�/4K���Ӆ��t*�R!+;1 @��>,'/
4t����e��7��+Z5�=S�¸�r�6�� �I��[l->$�B�eY)g���#�:҂ɢz!���d��E�5�*31nG#^7{3B�pyV���$
53]�������?	B�l|8{������"�
1�z�Dx�}KW��c�]�b ���}��/&��lݘc�1�@�W9�E���WK�>�����W_���	��8��x2���B�������"DQ*��F<\W�q<4$����Y��mu0O�q�V��vM3�^$�c�t��~��᳷�����o ���Ȃ��/L���h��I�$��M���& ���9/Ż>���P��qX��Exd�0��n1�O�X�o�U1s���M�g��~9�|*�ԍ���+��&��"��I� }���F��)��%��oq�?�Ѫj�"���*�V��Q�_!^V�z% �I�`v�p��XmzT�l������>�;9d'$��`"yj1��)�\V�1w�H� ����:�#e�9�E��Oi|��r����kR9f(�d}�f|(�]B��xI��ԭꐞo�T��Ĺ�[φt%�Z����$>!�l�aǢ!�%�k���y��8�p׌�詿x�u�ϫ��:KWD��u�+�9�����6�g��l���c�e1��eeUg��'g?y8r�ax��&� �/����q���1�4qՇ�Il������y z��H��>,�1�<�Kq���c�����JH�5�N��Xc�UFWi��z���ȷ��.h>QＦ7�f��=��(."��`�rt���R�C��9���iߨ�a�j�}XwX4��@XO��u�r\[ew�t�TQzn6��	��y5�e!Ɏ�V[[��W������oׄ������D]�1�9��VVwX��<�/Z��U�W#��s�T�T�+�����	�� 7����(�4�>�0��n�H��|����:O?�H�g�Z�9h��)��ض�ɬ�yV�ퟝ>�2�F�: �iU�"�{̉�'a#�<��^ytB�_�������p�xJ�=;����<܃׽�!㱒�K
�.��LqD�
{�&�`A���M�y�bɴ5����l^������|�i���WZv)��U ��Q�N��~N=�b��0yˆ>�zB�S_d��TOHK{�+����۶:�xg���<����)V�(AliB�	�^�}��T<�Hn�F�֣�F֧�,��&�A�~f����Џ��yaE+��a�;��d�����T`�ٷH*-�_Fw]�*h����u�L��j�����:�0iKO5�b��RT��ʧbF�%������MY±E�������Ǘ���f?W��bp]DX��8�ġ���mX�ڂ2�k����4n��l�����?��A�O�<rH����p�n�9���:h�}xxS��q�)�Ƴ����Ȭl��xҤڎ�}ER߉&���&����X�H[���<@�[���]���F���z�	@�h�p�^9��m�
(�lX
h��|V�l<c��+���BM�cvY��VQY��cq���_���Nec�ԴC&��J���JFq��m�� �̍��!�r��QI+d[�NŬ���h�-�t�Ѷ)�pt].���!TZ�R�W�v,�g��z��['kE �L���2��5�T!w�����it3q�
�W��������:�JnApG�'Y�H��"�������зB��p���˒$kW�1���QE<�T���j�T�@tk�0��R�YbX��S2�}�6��:݌�Q�� r��K̸ۜD�Fǯ�N�]ú$w����Bu|�����1Lk�W�a�r&AY��^ݼ2�k���{�l���g��(s:3�?.x���a6FTO$�q�JԢ��������.�L�?R@s��o`Ku![h�������"y��mnt3�{Ƽ�Ĕ硄�1J��@h�Z2�$����;�j�E�7�|���S����K�v��ɠJ��-���o��|���e�� �����]21g宁$ל��	H������mdN+}�0�b��Y�ቤXw�a���ŉ��ٹma�Վ��51�3)�o�e�9�b�5�����V6Q��'<�E��I��6Y���)di��@�<���]�B�P+f�6ֱ�QbQ~��c"93������=Z�~zM�	���i��\��1����w�Ї{w=L���;GP���Ry%��vm*�v��T�A&�nێ1�W��T@5��pB}Xh�������4���f�L�C�W3�I�wL��aW%���BUBҬ���ϡ�]������I��ҷ8*���ʃ���8l�FPo��/-#"�,N9Trg��6`�
��SiyM�M�튟C^ٛ�zxE˒��v�v�-�C�cl�h�Yw�l���)�{Z��O��d��E��+�r/b�B�Z�=G�l�6N�"���?Cg�DxoEт�V�(�=���"m�ϙ�r��"����KM��s}q�J�2�F1"�I��A��
q��Pr`"��$�=��<�Z�F��� ��ޅ׺��E�g��j�A�Ѐ5�S�z$�*M
��fQ����l� .�<
w��S� oo)Q�8pKaނ�\^!��*\/@������z�$�l�n��&�w�0Kq���Q�2a��{�6
���7��yy�؋�)7�����f'�O�;���������R�ة�*��H�D8&yŲ90���lu��|������|TB��M�>��?�`a�t�ǣ�X�Ϲh�R�]�r���$���6�s�֘��(��t�20�=�񦃠)����@�lK����n�#���,��������$o���~Ϛ��^8]�QV�[�Nk���m�P�-�]	Q��D�4b(Â��#_ǯW<m�2���f���
J�>H�S����[��jV)Tx��Ó=\$l��W,1u��Y���x�'��舩%��u��wLP ��ٖŖf�d؟7�y��{��O���n�,�P9p
#�&d#�.Q�������/��@|�x9����Ҽ�G�{�dVw$���Ro�Ӭ��=�7c^�,��'�ģl�aY_▱"b�[��M�8/c�
Yce�L��H��ꟓ�JofAfEP({�х�݁�6j�/�9ef<���MGt��B�����_g;�(`U�#�o�C��4~A�;��W�L��>��~dPG����P? 2�'�`�4��n�MYSO�-��F��aL:1�$�Ei�Z�vr`�'��e�Β
���*'�p�H��,��~��I�x�孼\�M(ڣ��7Bq���A�,!�jֻ؛�^�������ђtpC�E%�Pm
M=��B(i�\��;����y0P��'j���OJ�v�th�;��L���q�f�vߴ�R���3�� A���>�S�t 1������u�d,|��$ xe��D��P���l�ϧe�����ԡ�3��:�� D[l�"Ƞ�F��8՜��% ��_/E��Ĺ�]7T��t�m���5R$I���4	OU��u�Q!�@+ �x ��R�'P&n^^,N:.�fK,0���t���&���#������m���% �i
P:z.�o)��`�����%�}?"�;=Z
Y8�%<t���I[U��z���PQ+�����a9
8%'�D�a�K�Q˛� l`ķ�E �BSN}���N�o����[���X�e���P���"o3�q[�)��~PdE�2��[^�e�4LD���@ӳ�TÒ����V�\d �%���4�1t�E4�t�n�M\H�^`�x�����Z .;�W���3jѕ1�K��0d��hI�Xe�	z�G-�6���dS�lF��T�
pH�ed!�"��ƨt �i�]z��Y��'mQ_*�h,�y�99�e�	�xV��R�h�� ��l�d�!t}��|Kme�����ם줢��0
�zᜢ�R#C�"��@�G͢��D9���{v�Gh�^�N,�����ë�ӭc�lQ$F�%P�(����>�i0.s�z�#F��;�6�裻���Z�䄻xK����] �ף�H�������`*�@�^�	(gc��<�\�	��i��������$l���'��;|�m^����oh���B������Y��C�"��͂�^�k��Dd>ԕM�X��k��F� � #�/��1w
]�(�j�� [�j2h�d�܀Y��@���:*�<��m���K�-�&jѮ 44�qgb�Ua?1�5[[�ѰŽ %�#m�'Ik�v]�I�h;G_i�2�?^sw��Ͷ#S󀰼����e��]MH�7�'���{��T��u1*mI����a|���eS��aq���҈���5�1�O����} ���3����A�Զ�T���zj�&!ȣ��tгm6�x�F���p�J�[��2#T�9�CwCEQW�߅�9�*W�jP� ]wv	Ъ���_���6�乫�g�-���w�WG�G�̲��~C�y�d��M��?��l������_JӘ=|�r�y���<��g��-��*�]-�1lY��+??���v�G�z�r��d��JL�} k��|��tU�VS�g��B~�n�
����2Ԩ�r�+����݄����qGY%���s��봙�p�w<�\c��G�m�ԫ�:߻��MBn�FX!ήF6��Ѱ
c�/MM۞f�y�{sG�Y	���V��mF>�C��(g;�|��7hT�L�j�5o��8F��O������^�BWr�K��qj��]-��r~+?��E�g���#��V 4-x�@�e;���*��q,� ��.)v�]�{�����e�r\��\�L��ŉ t��������]ޔ,u���?"B�YŨIA���*��#��V�f� ��#|6y�^uCg[7���F7��(,�I��-�5Y�_�J|�%��a��9�?��M�E Ii�t��)�5�&/ ��M_�o�y]��/��q2|�g��m~P�`�e�����K��t�PDAraq��@@�=�Y^��@�3�_]�SY��ۺ9EDh�:�R�� j�}�C3{١(��P-�\���|;��N��ڍv��{��~k4��͏-%»����S���+�	��q�w8�@TP��Q�r(s��RDҊ�7-:=<rEc1B*qdV�We�H鞳��J�����w��т���L:�4����%��ءBߥ1D�
E��t���[��ỹ
'}�6�^�g"����0[!�D��'�o5�w	ENBԆ��T�������F�D��ض�&�D�]���6 ����A�`b�5��5�DH�̋^?a�\Y�իN&A.��L
e)B�ݻߎf���p�b�Vj"�%+�q�n9��%e4����;�no�kLZa�R�P�S�R�%5/��$��^�=���­[��e>��`7�l�*�0 �[}�Qr/?��h�כ��WK��ϸ�M"�z����T�hтu�ߞ�=~������m�ڣ�e���X���pë��0�g�h]��<Uz/��d]��=d�
h��P���J�HD
����%�M�����F(ם��Zr(��������b������Ϣ�ML���P��|?�'�y*~Z %8�PB�3x<�-Q�?���`�8}p���"5����CYMD%��j�q��r.��N��e�+��$��.+��&����鬒�.`�ݰdB��t���k�S8M`w��Yh�<N�n�1Xx��J�v�])hT��w�>C����Sn�3g�
>�?�p�	<NSU��'��n2
'�3az�)�k,�n��	c��4��5A:�����ay_n/�`#C]�+3�(=���{��Ĩ��򿶋|�g��5�6H�M̅q���Ie�L�f���������O3�9�0ݧ��t{���^P�SeG�Hf���B|�NY:F�a�'CS�I�<4*��J�w�壡��9[{t��.ؘÈ3��z�oN���z�
�94d~V�j�_�0��z�;�����`�:�����U��w[x
UvY��h��akq�[�<쁣i�{N��0�uuz�M,�T�!<C�������%s���������%��Ƙ}��^s�	���Kr/b>����d+*��ᐲ䎉H��������.��Ο5b�cu�����ry6�[X\e
�mɺ��m�qL�Fl�l	�T�1�Jű�RQ��ɦ��S1N&�L8M�H����h޴F݂�yi�����b���7"�����.��>!��
U7��{EC�b��\�SaU�����P�r��&�!���_Z��;-v��ý�8<��l$nP5����ȂP�p��/t��j��l^�'�2�����VEjHx8b�6.���x(��.KCA���8UZ4j�@�X�|(={TU��CM�V�a|h�lw=3	���"���A{�c�R��]6���	�Կ`��_u�x6������Tϐ1�T��먏�����4#oPz�9��i�1K(��������ch���E��j�!3zc���ˬ����\����ժ�G'�̣]�+}��C�	O'qN>H]�
��/'���虈�b������D���I,B+H�q)�nI�h	�+�$��E%"�k�;�_x��F�fJ��V�ṟ^4��VEK椔�Q#/�r&�U-b�5�ڿ�l鴕��n�|wQ���@wCH:�[���Ɲ�>����Vu�62Soo��]�M�a}`r�r�d��I����`��g߅���u
�GOw-ĴI�ߥ�d�K�N�.�Y��޺�c3&�L�����5��}'�h*^$tU���g��G�uPϦ���7X$dv���"��(�Ȅn!��Ĝ���:m�X>���0
@~;R�٧1��a��N�N�ph/���4�q��
O�e2�d����ܬ�YB���yc��J�a�w�i��70�E20b����6t�31�Fy�	�?J�����S��0�8]�NB�^���Mٶ�o�TP͚~�j��{)��x���`���~�V� ���V(�n�r�3���|k��9D*�)仓�}�=�<�}n�;;�kY�N=�>�1���h��U������unUpk�*Q��c,�J��� �2�a/iŭ���F�d�gDm�	�B�Mρ%|�g| L�"�_��lY�(?/_�b�v�s��EB@K�g�͇���$�z���ތ@����*�>���`����3�*��c�Ԝ�b��ehu$���v��&W��Ep��vH��q��5`�����aa{`x$im�d��[���|�=�n��ut��aCH�E���Ye$�I�-*���� 0���H���g��6��_���:�k��4�%4�̌>��Y��AD�m0���?�D�䝘�_�tpC[Q>O��.��v�O�-Y@4��pra��,��������������CmD�����y��s=� ���0�֣�ж�nx�u�TL������Գ���){Cq���j��hl�]�6b�����.��Z#���S.��'�A]Ĕo�'���s�:�;<.�j��c��͖���FfR(�d{}�kS=-��V��Tؒ���)�";��h=rgox`�|];6��/6��O�7�y23�%�٤�0��_��]��ڄ���LY�Ú���ŗ�nE!��D9�6L0�<q��dYǘ�ŉ=h5�е� �{�;�%Z4e�3��Mb�i�7A]^'Rb�ƙcW��7�{��!���(ڧ������'% �䅙b��]	!fr �/5�]7^��n�@z������\�ɤ���W�n	Tl!KC��P�!a�\E�ɸ�e�@��i#�'��TҞ�r��k�B�����JO�x�wa]��.8���vQM�/ݩ��Y�@����d�a����M��X���+yF/�o��U� J���#�_㸘bZ�� ��|1`�.�ߞN�����;��ʲW��>l�nz^�� Z�N����b��ڔ��p�6Oo-����D@:#$gɳ�gqX����~#� j��<_�T+�,�f�KU]ms�)�-������H%j���$l�#��59���z�e�6>#˧��������f�g��@ǒ�Z�������/G
C�͟�]^�{A`P�hf��_����M���a7�f�]a�/��TF���f��J��ɀ���)�p�;�u������p%��Z�#���qf�Ԩ�"���冕N����
C>٤ֶ���3��F
j�lr��.�"*�FH7:���Gu�������XD�}���烙�A�oq��Ӣ���:���S4�XDs-�~g���2ip���hF���x��B�AC��#$"��t��U�ƨ�X3�<�dF.�M�E�	������G��t-��؇���pC�Z*|�&W��)2�6X�-����Po լA���z���HȘ��	�}�Oѣ�MoгK*�o؄9�������p�q_� 7}h[�\��J�� c�V��\�HXf������x��Wɭ1��Aa>Vr!6����V#oL'�Mno���1 ����'��V���.'��Q���t��þ-B� �Մ��]��QD���E��&��>����Z$[�=������
B�ei=����O
O���M��b"x!:�Uj$�bB�X�Ѫ�KK�ay�c49w-��ԋf+���uffN����z182�$�,�t5S`i�$�l>�0�vr)(H��+_)���H� ~�|��]Б�h�@��1����a�3�۴Y�@U�� ��S�� vU	��O����U����Z���O�%�k�q�L[�|��:R�z>Z�(/+
��j��[� ���	��X���<�i�q���Ho�Q�A��4��Q��Ԛ���F��>x�~y�M��I4�ھ��w� �xW�}��9`	|� ���Tآ���J���h�.:����!��s#of6'?h[u��!ɰ��
$}�����#m���p:�d'��A�pnn˷^nM�)��j��h����oi�K�Œ����<� Ɔ��U@��v����S�J\^�(l�S��L�n�zk�����Q�.$�����j�Tx�W��㪛�$�f�.�c��$*�4r}��������w���Y}����A�;�e��g�m&�?��66X�l0�xS1���[����{X`�ly�����+ZC��,pi�åv)c%Hc="�5N�3 �,\�V<(1����� ���w NG3[�WO�U��mC!��1nO��5��}k��\W�D�FK��XT�L��H�4���h/	�/�`k������-�tб���q�R�5��
�^ ��)�}��C��P�/<�ӥ�K���C;t�:c�J����|Eb��m�v�9\�E[b��QGPۊ�� �٪p�+��%`��t�|���7YMr�oX�"�H\�4�	!6k�����K{Wѓ��.��1�lN&U�f%b����-�q�Wu�L|���v0����\���_�r�6��J�<�^B��	*�:����r���S\s�T/���)l���B�zg���Q8�l�uz�'ia\j���2�(������ܹ
N3�
�S#� =�pmj���0v��
J�͔�90�ߔ��F{�;�|�Hui;S�L����#^\����i���1��慩�б�U�M7�+ƪ3�;#�Tu"��Rݗ4"�M&�X(�?$Y������A�Z���N��]��-��ɋ�󷠞[+i5�Ѵ��D��.i-,f �K]m"}����P�t���/U��g��9� w��;S�M��	��\�0��t#���ٜ����d�w*`4I�)��,�8uh��P���^�7\]�z�q�S�_=��^K�C�¼D	��;�]:�Fuuù��Y�W׵��'8�5+,�$����i�v� K��a�u�>�7�X�G����U&��k�Z��~hR�\�=5^�K�W)�m��΅S��́�\���zV�X��r�ؼ�E���O/�R�zQ��Ko��@*زU��٦��)��u&��j�$��m��2�X7��+r~���e�=��B3 ����=���Oȸ
y��v&�<s�Sv���լc�����5"��'GKQ؜�5oRH�{��Г�D�~x�U���(BJ�.�f��X�hvu�"V��M1F���d�k1�`[' O�[�3��e~� �c���a����qխʗ?<e�U)��WH��=�Zsa\��n^�y���~=�)����MeI��1+=��b�.��k<��0PƏ#�w�(i���<D�<ʌ(k�֍������:	ɋj)8H���ϻA�U8�j��$��dgOe����L[���,���-��G��;	HP�L�N��q}y��7>�WҁIܙܰ��L ��"l��]Z��'��_����a��  �mQDC�%ܵ��d�$�V��,E���,.b�!Mb�¬�c����'���V�@�]ؗa=��s�K��)�
�5�Wܨ�q��%�N�T?ep�	�s�	�D�ރ�m��Mt�h��ʠXO�Y�>&o���$�Ͳ]��7U.5��>�DO��(�"�%bo��*�����b�,��d˼F4%\ �]!`�F0�͟l>����Y��.m\$����1�������{Z�����]�<����7"~D���Q�y�!�-�Ve*ܗy�ᴉ�C-ʎ�2��(D��E�̰��!@W����t�q�Q�U8�;��~��q�G%9�؃��ӭl��y�U94���~�#�	%��^7&/�B��D�� �HT�����Ủ�`��wq�e��ʯ�e�t]$���o 'e��m�J�V����9�Q��u11��S� Ye��FFd���n����s:I~�[09* qI���<64@�s���]�9�˦��
�bI�,Gg1�V��&��V�2��i��ˈxN�CT�r:����H���Y����)t��AU��5]@Z�Nާ�Gۂ�vD͸7���:e�2?��ڀ�O�"��xvf"W�Cx/ɗ��w8�H�^ǜ��@��{68�Ғy�dͅ�VB���Fy��:�T��c��+9g�.�Қ{߷�~�&������ϪQ��L`ξ4��q�+�Hy_�bpk|�e�#�^����Z�����hæ�K)�!s��1�\�/��~C#P����`*X�1�DBt�{
*�$N$��c�́|2߅�� d��Fq�Sa�4;u<����F���^� �A.�*ڛ���_����0���y��'�{o�����q�t���Ą��0���O�[+��w���ZK������(����� �����R@�P��O����}S���1�Ɛ'/�B�/��zzJ��u�l}F��l?��$��!;aE6�C�L��e�=@ٓh���[Y��@��"���x��?Z:a��@m_G�3;���]w��~Y�(ր[��5k���2�W+�F.���oi}b��&�5�%&O�> �@ aG�M����|`���6�A8I9��[��*��؟u>1��tF�h�X]�V��U ��H�w�y�I�������x�ht�����9z���q�E)~7��\,�j0�V0ZxO�+�B���"#'v3p��e�Q�r3�HNÎ~���-��Xy�c_�ʺ�s��u=�_�7a�$vgZUg���`>�(��>V���c�ɲL��X��E۵��3����Aݕ��p�cgQR�w ְ�ɵ���$��l���9�V�&~��d!J5�BYD��|k���Zt��]c�\;�+%��U��Qd!�g��:�P�Ű�`_���7Pg0aJ�%�Kbl��#�a��&y��!�V�s�Q�̃�/�^����D�=����(�$3��[�&��I:�����m��)­]y5�� �� )���� ��]����Z���kTo�3�r_e��)�4�W�� F��/�ے��K�%�:q>n �U)0Q9��|ߌ��%�0U���
�%� 4�3l����$��)a�cF��@�@}�U6%��G]�ea KbnJ�����'a�Db�RĎ�"��l秋���ovĆ�ъ�P�N����R�B�wpG������D'>y�ɬ��nw��X�崡a�G�'\�*$���zP���(��p�$��#GwWK� ��5�L����o'����6\���LǽF�H�B�Z��F����'����~�l�u)������ج�޹���<�E ��J�w'��PEiH:K��@_-=!��q�O
r�+��c��31rle�+~��J/]���{���@!V2w�G�8�z��T�;�������(;���֟�����㪻�2��[�S*7T`C������d�����������<�"�����V��I�Ұ����Q6��an�p}�5��/b��w�!O#Ť]w͖"�'P�b�w�b�G0�j�$���Ï�^-c�q�C״�ˉ{�2K7[������n@�!�;4h@<��'���Y����j��P��7�R	'���o�ͺ�g��a'�|"�U$be�l�ai���C���j���(�X
j@~�G�*��6����+���
���uFM�B>�����3j��+p%.,�.����[�B��1����qo�ꂪJ��������Bԇ�|L|��?<`dS�����*&|_\��az�1� 6�U���|�W�b����:Ku���7�������, =�u�`��E9D�ͷ��0���D�i�\���Ӭ5xxU���nzM��2��v@�Y7�.�5�>�L<��y��]]�[��_#(wZ͜�K�	�O�;�?K��/_�`�� �+@�K��2"�$P��A��KJ��q�+G<�����j����K��83�+7��%�a>ո���Ȝ
C�"�B�^)���d���J9$�LJ��h(���hs�~�1v"{i
�����PGP5mm>��I�{�a�T���L�v(�$J)I�q�MX�����r��������J"��]v�[�}M͂3c{Dꑅ��HJxE���u4�e>v�-O�^b��NYo�TR}/������Բ��N������4KM�+@��ul^�����+����u�����@]�h����^&�C��O�Nկ�@!�Uw�ADv��I���F��T� �Y�Sb��K�BW�j��rd���ƴp	 �2��ĺU비��l�Ώ!�qk��aޟg�:���!rߦҽ���UX�"��ij7���߁5_���k>#D^�����)ǬZШ]{
�;��'�/�vݒ��F�q��i�\��pe�j&�V�q?���"Z�1K�!�ܿlb8xD����խ���J����b��ֶQ��>Y�j� �4�"h��]Q�򩠲�?9����zx�Ml�i��w����&"�B�Z��j?t����vi�|Zzk�'�e@Sh.��.�ߜ�Q;�Mu�L�Z��Al}"�+<�OTs���v��c��{A*�цiNe{�WY�>�n@�"K\AMU��zwx��/֚Xi߮���ȱ��Y�1�� �s�.��j�n��M���Y�l�R�i@�F�O�)m��d~�����z&W�S=��`@��8ou�|�س��lǨ��y��/(d���U��4�,�[��ӳ���؜��D<��]ġYҧN=y$���(>K-��ݲ�ytʝI�s)Q2�4D��'�S�FK���Q�v�z��7�n	N�YE�|Յ�k��G�ǭ�w)�G�)�S� q���F��{��C����kW��wd�H�zz�>ׇ�Q^17S�N���jO�.v�45���������]�2�����C����,]m��K(2Uۀ�z�@�OA�>�X��c�?7Ȃ���P���7��\ĄOp����	tyfq[�dR)�X�%����m��Fu亥�H���:E=20���[{�Ja�i�<	}�k�����'�t���D@η[M	����H��w#�OU� A~�l�+Xa����S�i�Gn}1�;MQ��Z��l��]��vym6]Oct'�J�tJdk�0m��dV���l����B��x��@y�;��m�˴���S��h���=��f�|\d2��<,��
c�d�<�� f�y� �2滅h��n8��i�< �a��l�M��r0,�hvR�0�F�4�
�[���?6Y��NG�;�����T7X�� T�e����ƑSp�*������X�	�~E3�v�L�
_�(�.�Ƌ��F�C\56�4�����d��]�6~��/?ą��Q8�4u鋼�����{ �|��`�1�?ϝ�٤�����a��,��͒�=Gm����jw���]�ҿt]V'7�T:&-�A�g,0|ߊ�×0�I�(<���`�Ф�t�U�rE����&ܺs���<�7�)�����Q�]c!�3(t{о�Qo�y17�#`�[EG��4?�t&��'��`�|�õ��Y6��ym�w0����Qw~|��XYw5f'���.��H�pLT�ʭM݋�ꒊ%�4�|*�[\���4J�7��ﯜ�gk(��x6�;�H���k8~gv�{}"�4��^!a[{hBB ǳt��_��9�I�t�;�V��ğ�±��\9 �Oa�]�����-�7���W�p�h���ƛ4����RBL>Ob�6魤4���I�6��m(�U��[Y�P!���U����0"�&v&�B�W�K�c�u��q��!����9�_R�UK�-v�t�fn~�bb���C�BW�{��w�GI�ř���xl47^_��}�y�h�C��܈'�
����~!C�S�`tkf0;�hx�g��R��e�Db3������\��׍R��X�V��W[U^r���4hx�;3�+�\@r�F�l:yd�6D�Z�0�G��MJ�����U����ՌD=���N�M��寷Y��v��B)�E������
���;C�o�-��د��,.��9v�m�ae�3�"Q��S����<��-`J�a_L�C��{tY��~�co-d3<ß��;��ش�F�~TO`�3�L�&Y��K_��v�ՎK�7��Y�@��bL�1w5}��l�_�u������GV��w�R�˯�0��� �a��yqՋTL��s�d�=g���Њ�6��"l�oT��̗����o�<�] �yY��U�k�o�~�g�h�}�.�=�z	��h���
�灊6�Ո�)6Gyr�S��sr*S��ζ�[����x���ȯv9Yn�v$���K<�+�$��m�<&lZB�q��v��W|M���`d�M;Yak<��ZZm���=^�'�5�q쟯�<�쿙3�`�$>L�}�����sό�(���v�(�p�:�U0V�7�U��R:\>f2�}�q�bR�\{�XQ�8TT��՝�3�0���Q�ќ��jig�@�����晌��'��׻��?7A
?��2?V�0�)S�b���(�r\�(��[��璍�J�>�o��M��A�cY�!���\s�̩���Z��y����>g��&T�A��G˅�6���V<x��7J�gδwTi���J 49fɫ�V٥o����Y���'/.ջE�ne���Ks�I�V{����kU����D.���o��b��]7�y��S��]f\��V7��,��^*+q���읙=�јp*�m΋��}U �D|.�WT�9>5H��	d�qZ��~�P	TWN�_{�P6z��[x��$:�|s�<�`]�[�E�ZG3l�r�M˩�SW�i�0�ԧ��|nC[���Ҫg6!��uc	Ϭo̡�EcJ����O�PRC1��n|�W����{��{��f��1N����1c���6�z�Al�'��ǩ��8�Pg�I>ɹh�\���,���Tp��`��?���7����9%xG(��MX�ӭu�����N�@�Z��ޤK�  ���G���a	Zb �! ��q�I����D��#C�w��f6�w�c&5�����2��t:�L*
i�4��� ю��D�&{�ԅ�v[�:m��1 獴H�l�t��,;R_�������m�+�xDO��=o�	Ȱ��s`/��k�X�H���Y��i��'cBG����ỏ��N�,�N�3ȿ���G�^�6|k�2��o�z��%����!�����a<@�~&�����~�m;<�2�C,7�
�v�4(i��D��vJa��Ks5F��@f���9���nq�z��$3q��	F/�sS�c�z�QX�I�b��u����UN�8��Л�0W.}Is���:��K-=����3���9����.v�c;������q��x9�L�0{�a����)�ycV�`x����`B�T�����pZ�m��}߶o��-0���K��Q�s��VP ɡ���j���-USs�m��}�L�5��+�	��nJ��nVp��K^�����k}<_�P�:��{�AMQ�S[�Ж�`qڳk�@�2r������\��h5;z\n���}zԶ�%�����5�:��������G���uL�{�u���#��6�qi������x����m��")�>Z�e�%�	���h��Oi�T��:�b[��A٥|͒�l�Xt�k~�rdď0�"�b�|d���8qylN	R��nBi��{셯��X�Tʦ~P�.�x8 ~�r��8�\tc��SWc�=ogҼ���������s��)�I��N����1��Q´+t�>��6��Ͷ�YyI�B�(�8lI��x�BoC��������o	�+laI?����yަ��XV�в1]%����Ie�޵�|��c��1uH.� U��rz]�Mb����}0�+�����&k�XCW�'��0����|���K�s�s^�v�"�h�t�������Q~���2L�G����P*?�V�uL��A��r����4V��ۖ-}��Dt'������6��̑xʯp=֯�fbe(���z{AT�g�F˼|���;�W^dd��B1�9b�cn����% ֲ��f=h���P��9�ѩ����}�MPG�6h�F[��/�~krd�+�buB����N�s��6$ED�\^�*�s恩1=����bj 5��*d_Pض�.@/�|ѕ�ڀ�z���C0���k#���;�Q\7�Dhk�ܒو�� )�g�K�����+�O_�l��)�sg��%�l���XEǰм:����B[������j[�_�~12�_] ��/����b(����޵m/���o��ws��>����=�k#����
��"�ݛj����߻$j�xM-h8��+[�}o��(�SzE*�:,��H��fG�:1�9�+tUH�S#fd$�:�r���� ��|�)2��KNW6�]���p�E�`��o��Q�q��@z)0��H�<�"#���^��0r,pP��ES7%8�yt�B�� �|,yRNIo������ǝ`VK��	$��Q�Z��_�p^��Q�B�_|�_�p	ǩ�l��ˮK_[��i�A���4mD])'}�����D2Ĭ����{�f���-7xp�{�>.^�Y���N����G��U�T��$X������"���k�K[j`�B��uؼ>��=���JbB^����[�_�:ہ.�E$+9R�WLiA[�a��.��R�T�9���V�Y���"��H����$�;������(��ODff�����6t�7?#��Ռ��e��Jփ	OsS$��XY�kR��BB��u��!#2F�m��Kb��� �:���?Qe��dm_��t��ߋ��Rӧ���ۀ/k'���|�߰�=«������׸VhpaŘ9�GQW8䑎m)�˨	-�C��Աۇ�{�w�A%@y�
t�]��خث3=+ .�҇p)���K@Ro3�f\FEت>�z��CE�'��3���(י7[��ƭ��Z��-Z���+k^��x��ݱ��W�>�I������f4�[�"��ɉ:a?�Z�����)�a0;���2�fP^f��9#�_��L�[�Ф�