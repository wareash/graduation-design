��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e����d���f{��@����S��>���4{��ת�AO�Q{���9��p����S'&�������8z	]��/��X��~ �`a=�\�|�?�W㒽7 �Gp�͌Dm��ӧ[xu�z���aS�&M*���~�?O�5���lc	w�b�`�(�,�p�'�$'��	�?4;�L������+��W^�Q�]7
�_�V�eM��)���^W���p��Du�E��z~޲L�.�9��;�Gh-�}�u`�sg�MBކdG��7����pFO[!��ϻ"�sc�i$+4K��o$7V����+����	���Bت��
WMT�?��fBf'��b�f&[�zf�&����#�-�yO\:�t梨� �o�Mv��h�<���7܂�=SG�)�W!��⯁�3*v�	�ʚ	To��g���ɿk#ý�z�N�T�f8|��$��Ԯ���UPX?Yd�<��2�1�����PW��Ø~	���70kou�7P����O%�5\Z�h����ꀵ_%la�u}hRI�M4Y��n1h�?rΤ�-����
yS�h������g' G�2.�]bd�'�@��F���D��ުg�\�>��]x;L�����$�*���@5��������}a���"�J���+(�Q�D:�<fR�M��_m�!@1<`0%;vxowK�L�8ȿp���Q���@�w��O��*
��e��x8����aB�v����zY��Sŏ$��D7�(w�J��۾�</)j�>�����
��ST����j���״�$]����k[|���/��!@���(�*���hU.�ά���į#"u�Z�v�#�[�����5����o8��<�}(y�������;Uqi��<$�Ԟ,yx~W�ɲ��äH (�DHB.���1�$�Ha�!q��'�R������E�`�T�]�#�s0g�3U������J�)����b	�o��.i���7�����	�{?��g��`�0U�l��{�a��i�T�?�?V� 51� 4�d2D�F���nH���RxO�6�����X���!D$<���Ȥ��!�,���nV#k8l��o4
y͕oA�;S'��Q3SۤJ���ac��5�r�cy�櫞�� >���f����e���m=�V��u�R�L��.��ܪe��
��gy�)>�0׉=��{��C���L����+�5G��ts������Ƃ��l�(bg}������zpm;zuW|�xu�j8��}��{J�n�02b<�n��}"_3Ք=�%T>2����~���̇V�>������yr �\��p�����H"'x
���鍬�An�!��J�\|�Ȇ�/��M����a{�/t�h�l�g��� �hPXO�l %�� YV�5	; '[ԭu����rk;:���jKI��`?KB�Ju>�����o�y����<�df���I���� ����/��35���3�!<~�L"dv}�JlK�Q�m�}��dYUQ�����qs�=Z	~�6N���!�#�7���"F>�b�I|H���/�[x�ب�K$`���`$o̓�(�Za�!�o{��-��@�>�J�+�u����bL�����(߃��s��r�.f(��l�0��I�uB\��H*ن�?Mjc�ǨH���_��t������I�H�� ��dT��� ���d�|�R{��P���x$���
KV�=4���P��(^N�����f�"'��2{",�K{=
�S���������p�+��U�p�m��/�[�Ֆ*��һ�
���HEq�l���Ol
6昞_6�ԵY����<�s��.d�� �L`Ħ����oܣti* �Y ����e���Vņ�餹�
T+���Vl��k[���(�P���Ӌ��P����P��:::�h)Ü)�2!�|ڬ ���&�~ԗ[cy����6Y�ݰR}�t�e��Y����W��c�U�S�)3Ll��Ɋ&yS�ͪ�V�Pf��e�`�3�}�/g�ղ�]�h�T(�KAE*��(��d�A�"6�>������ZF�>Wĵׁsf8�U�|oA3�����;���h�`�% �X�tØ��	t@!O������◪Y�~����:�K�4uN���2�Vh����G�e֤��O��[g���Gh�_*��F� ��Kfg^00��0�v��y[���t�'=rt�����5�<B�ӐG���ϯ�n�͋ R�;IQ6�>�2n��.�z���>��٘!��+|�t�qQq{���X\�m�/�w��_81��<�.-R�nv1�G�a��R���YM#K�~��u���|����Z��U�l/�����>��c0�7C���2�*�J�hk�����T�\������?����{|��h�sA%����Dw����wPC��ҫc��}�%���t["cQ��.��X��&0���5��8�����.獴�ZٓKZ��䖎�V���{*�=��|ez��2%��9�$<Kupi��24��' !$Ğ#�~���t�N �C7Eq5R>�7�KK�el�N��	.�h�+#=������Z�9 �mZ� �ᡜ���6�"��j�og ����ۯ� IA����IO��m:�?�H�F����u���/��U}P�j]J��&ͨ�e�Kfp< F��j9W���aN�.��Y=.�j'ߑ2)v$��f[�a�Hkɉ,�Yq�Q��S��LJ��zGi(���q�5�!�ˢ�G"94o+/�P=���[���=��~+��?�wK�l�}�:�������aY��#p�D���c+��#�=n�^�_�����>J*9c!:t�fw.ybv.��I�o�U�d}g���M|��=���32��$p:�5q�� ���VH��<%���|��Π;@LtCp�B1i�H�As�<ٔ��B�8+
I���f\��� !D��3�ˡ��w~&�EoK��s�W����S�Q>t���~-wv,�CU�ĺ(p)G�l	�jAܓ�W�W�^AX��3 ���d��:�فD�k�6wSl�MhW/`V'3����;�ۋ��C%?�`1K���2@i�Fp�d�D㰙,�mnJ��e��Q"�}��:���{@0䝐 ��\�˛^�h�F��X�Pr�JF���_u�`����a$�|�C;Y��qW�f�|ݎ)®���:��MV%�	2zZocq}~l Lȱ���s`�>�#Ե�XL�j�{��|� �P�^ez+2�G���2N�vc�!����%B;x�d���qϸ
:xe�)�	�i`�%�K�ʑ������
�<=^]f+(�kg��ܲ�OW�:G��:�n�d}��e�~�_9�^�A���i����d'C���P�+x�~�ge^J�_u,��d��� 8 �d�����������T@	!	�&Wy��0�҃��^R�)7�����Z�{~:����Ē�_�m��>dt�>x�MJ//����M��U�T����:J���l 4�aG��Ǟ�XL�h���1PJ�㞄\��m�{�w���T����6��������y��iyw��xE�K��T9@��ӵ��B.��k���d)�˴ז���d�UV��-B�_������2��(v�G����5ʉO�����Vȳj�oɷ�9��.ųuS2�o���*X@�i��,��`�G�h�Q��c|R�>)<V*��:B�"t�d!��=8BZ`��O]����4�&���S��Ú{��¢ř�`u|7�87��6��+{o��Y�d�3\��r�P�������#.�g�p{$y��;f��ƽ���-QvN�7�!���> �Т����1�}�#<���	E�lq��`�=�a�絔ז��LyW�
�(�Qӎӭ��$�, f�+g�_k7~I"�t�w�P/�k`�^��ߙ�j�کo3��Vt�L�wN�X��-A�D���q:È�����}�2�k2b�-�����M$������
?B<��QAb���,��_V�l�T����7	[���q��~�i���k��|2a��ĤRd�$�e�۠�,ث;�&�� ���_���3�w.�G���5������-�*�vqH�X�hQN̆(�ʂ�얄�_�R�vT�3hG��HG�D���Lc?�A�#'�C�VB���CU�{����\����h ]�-�˺l��U!XS��,l5�ѩ>�k
@P�f%^:����PȤ�:fw�a!���.��4�M�ǘ�fsW����{l��B�o���Si���A��%ʎ�AJ��O�ܙ��_��c7����$�gz���(
m�Vp ��ȑ.�EM���<�ۆ�s��s��'� z��3�ܚgQ�j�����[ӂ�g�*_�[��KDɹˍZ�ו�2<�����\K�����Kd0��xǻ�b��0֔�[r�OT�(7^��>X�"��R���P�BW�����i���몆ُIݴ_}�y��u�POC��m�L��gt�-$��!o���Ҋ�������2ŬY KK��h�칩�_��"��5�3���S�hG��P��i�"�s7{�����e�O�Ȃ��lz����(�׿�� �,#���pRFVef<�_W�in��3�����E
���Eu�+�1���8ُ�n84Y�FS�y�2�9�Gj��XQ�g�&�F�4��N�5�K)�K�O
O�����x� ­)���t�3�O�NU����H�%�6*�`B�8��,��[?+@�Ʌ�d���#�I?��Ho����Ί�_�'xiU��l`�G����P��3=D�0sn᎟�ԫRi�H��ݚ���դ�2T�B�ޗA��RKZ!dǌ�'�����@L��
��M҈��OZ���GO˦-6k��"���V���V���e�3�� �n8�$G>�i�A����ƥ��Ɓ�	�N���C����O'@���>�
|A���A��PȂ�:"��gd:�C�G|���.��GcYE�,B�$�sA)�d%��i�yZO���I�B�[b��X��-�>%$ 
�3ZI����M�K>�ј>���AL���u�ҩ$FSb��j�K�,�
N���kܘ�6w-f�ci�Y�և
��Եri���à�`��<ƭ!����b�"%2��2 �^����k�^)�>_GZ���9q4��;y����k)��<D,��G�=_m[&C�5Im:�p�&PQ{����80���FHM��y����J���W�j��+�+	�%��BX:J^o/3�������[R�=Ų�q�����;����(~�"�tA;�5598�@��uLt��*Y��8�f��xD:`,���ZztNliV���� �K?�r,��h�!j�h#����}>>e��{u��f�s4�`]j(�a�ԫO�����s�-�{��`�_��ƣ���.��9T�R?�A/J�G�b8����<S�L�u�i�O1'��A��_N�����d|����%ُ��
6+R2q��H~����V���^��6Y����Eq��3�u򳍳�F��3o�D|��"GA�-�T-`��ųXd�������ɖ� �Sع3`y��f�|�OM�Jt��tk\�m��4�Q��[{E��s�����w:<mo�%��@�Z��`>N?.G����Y���1$�#3T���<2
����}Ǌ���H&ʙ���\x��9
�ŃEܜ��-;�K�ӪcT/�~vW�[+�G�E�I�`��d*�8�=޳R���u72ap���,Iq�fY$��iө��B1f*0B@&_=R���PR�١X��?�T�|A���x-
�fb�p�����d__m�+�B�Y������R��������NE0�'�b^!tJ���8�<)X&�LV�l��qh*�Uω �hK�s�o�[ĲN��֗>!������LY�u ��F��O�����3��Q��QGKA��;�Џ4t�&��D �|W��ȡ� ��ݸO�n��F!њq�˙��=����2��i$�i�\{��C:������ ה��Ϻ&I���j���-�;����OOrB֔��s��cl�/�����8F	b��6m� ���m�ި@�Vo��Ͽ�r�r�W:����g�\P�1�N�%��J�q�p����+�n��.@�Ͻ�|0���=U��s�(Ԁ(�V}�K���n�R�'���b&�ܦV����s��H �FB����=����!��}<�Z���~;Gf�E&�,ļ���e|�|��׾9�%S���a�x�R0��
�i��=�WK>�;�
A)���-�>��s�,Y۪�O'�'PMN8���]�}�d]�%���k�VEVSg���~�ٓZ�<�Ia��?D;����,�-k�1�â�m���N��mCz��F��x�v�Rb7Ӡ����nB���-�AL�-�\Kp�wԸet�H`=K>�Jי,R��4�������)ㆃ	7��;�'������A	8��v9yQ��?��nl���A�1�m�"{�vY��xB�6��yM�.���{~Ių���)j߾f|�K�~ʘ&�f������u~�;��8q<
��Թ(���8��w��o�V(��wH~yT���_����)2v�vN �s:���e,f+��1�|��}�v ���'���m�`k�\7k6��q�1s5A����DD�o��[l�I�\�\}���q�[�=!�`R�"��Umڷ�j���e?'hJ$�|Sۋ�I*�#4MX$��mM��\4{���.Y� M���+B��rC;�åワUN�R�uT��a���b�8{����9�[�&?d�pӌ$U�T���c��OK�����1A�Ζި���7
�����H]l����ouH�����Z,��.+�:�}��Lw�K�+�7�Z��p�]8�����N��g|ўMZ� z�+�V�����|�
o���"�jXB�A��=�i*�����4�\&��V�'
����{\q.�@���J� E�6����;��c-T�(TZ��1������_�ޭ�,��Wi����֜����eNOq�yk�L�׏x`�-��Ӽ�^���ŀ^Y-Io�a����*'�^� 6o�R��^NHݳ��7FGfi��R��v�U#ؖr�
�e�p��p4*�7�k Vph��0"�Mȳ^kW��'V�bZ�Y�6���MF'H7y�|f�~Mt.�nle /�8N��O��=�5�r˜�0|o}]��%��g=I�|���Ge�Qv?ɓ�!�*Em� qP5�`r|�t>pE#�/�n�'��5mq��u��S຾Ԛ���NY�����_z��J�XnȶY�8�1WEQ����a�����lC�E!�?q�2���eW��~h)TJ^	����AP��W��> ^�G =M�x��^���@����a�!�u���)&fA��׿��?0��������Ww�,|ޮ��K_'B�������#��>�����$��{���@��A����J(T���8���oz��X��z*&Y�za�"��-2v�/�^F ����v���lW�#����#��F�W� �d�LNk��4^�������'�H�|���)��`(�&B��͢!���DK��Ġ��T5RwӦ��j�ͦ�V%��Ӝ�6}A��:B�q3������
$v
�&�-�Ϥs��.x��I�q19ʫ�A�w�����o�%�VK񕁬�*8ʅrra.,�:�O��]�8�T`E�5������	{8���KB���pV�Y�D�a�t����먳��"h!�����)���O�$9�[Y��룜��?��Ji���l��.�M���q�Qn�!�cx-�(�����w�^�ͼ 7f߄L�k�:<������%�.Ҷa��:~��sic�b��Ȭ@��Ԏ���n0��~{p�*�( ��ذ/O�"�O�c�c�����|T� %_����-�Oǩ	}�Z(H߬���뷦�f?��P��!�5�^��Y(@��ԷKW/o��v�T�2�L�:ff�����w)� �o0�c- ��
+s���T>�@���c�˂x��X�`��5��|S���@�4(�;�/��WВ��2x�w��,S�n�^#'��8ݵf�2܀�� �l����FSG�Ɲ�bUIN ��FR(�<��LX��j���%�֛�8�HCy=�d��w����q\�ً$5(`�[6 nJJqYC)>�"^]��]���Ε��\����9�Cu r��juQm�Q�H����i3#g#*���zm��@]gmV=A�����Z�2���{��\ƟaF�OX�~����U'��z��O�K�s�����w�p��A�&&);��jC}=��pل�="Pai����S��3)���TI%P
�f=�ra��lq( �[�Sv��p��E&��D"0����>�
C6���I�<m����R%�\@�Rf�<Ξ�*z�;���#�5��xb��?_�uú�AEq~͛��Mw�>w��~���w9����F����`��]�zQ��֍UD��H����M��6��-�dB�bI�Q~�qvO+X�Q�	�O��`d����!J����g묥�4̵��'��Uu���<�f8Ew��]�fi.C��P]�\K&D�^ڮR-��]���<J���.� �M�qw��z?n��/��6��c��;�0��p�a�@�\�b~���̠����@^�]kբj��7��鶘�f���0�#ݥ?}���M�f�Q�0U�^����dA6E�
e�tM�L���$p<�|��ݯ��1���;^�l�fU8.����iH�
�[K�0U����"i9��p!w�M0�
�{X��!o��Ž����31GO����0qt���?
�B\&�`�
�&��{����6��g�I�'����9��w�Z_6c�3�d%�����M����:Y�J>�sw�v��dZy�s���r��Xaz��r���VWқbf�j�<	o怓P�%!�YUm����'�g;w���T�D<۠,m��8|4�:��f�Ԕ��Ț%g��Z.��ϙ���x�0�B6��kU�*�ε&{�&l�'˄����'�瀭�y����/��HR�ѯ�陌��uKi�NB 9\���������iF,��hۺ*L��5�'��+춟ʄ��"U��wJH$l�����V���S�>�8��6ꞥ6�6��C���e������![�m�w
��z�!�hZ|*;�M��<}����[��=	�`-��yO�>`ayD�B}cu�<I� ,$dd�.����#�u�����&�W@mf6��8Pc��(pr^��ߎ���wG��Rh�'�椰����E��LԧE���dв��*�[Χ��1XQ�F{���E�F�M���{:�&H���	��B�^A1�'�k]w��m�Tѽ��Ƶ��^ì���)����6����=?v��L�O�#�w(J�f	���U�{��O�%ؐ\�:����R��TɜG���UIˬ��Kظk������*�^�+Tl~��)8�t����\}p#����ZZ��|�bw�;$*���-�(�e�|1�x�Es�r��SLhl�� x�P�kF�#��>�q^�3̛��=4e���i�-�j��6g�Y��f5B���3�\�\���{����Z�`au:?�P~L�'���� @Kсc[���9I|��sO���/��o2Dh�S��b:����.h\�d�n��#h�t�>�N�Uo}ӧOՒ���^|��z��$�������m���dMElRV��K�K1c�$��P��f����,��?1G	�)�h� q��ߔX��_뙋MVi��zN����0��O{m)a_t=�9~���r^�v)@t��q2�����I9t��M�Ǆ�ݐ�og@���a���6�f;k�p�s4|�3z^N�0`�Z��PWF���
���2Ns��lX�� �����?�L8�qI�#J�L&n`[ꔓ%e״ϣ�>.�E�2�V$0����W��$�7�gn��@c\�ٺ�2�%��y�b��QK;Ȥ#א���V���2>.��3�B�t�¤��g�p�}㓭amf�:���& �{<ؕ����Ü������������@�N,ԂnZ�<����ƙc�5�kXu8��G8l�p�s��e�pNCst�@�vh�qN]����m6&"�M�N�X����o���no��������)z~?�H�nO��	PG�	;1x��� ��`�3ڃ:|����820%B�c"�JN���\�r/h1�K���z	O���k(����>�ӝ��+�%��^�l��_���Ӈ�<��iMߣs�|T���/𗷳QL�)|��	X�!AB7ĭ^�F���4�>M������쒎@8���g�H��W��������܂��#����=�N���ٺg��@�=�r�^�w�����`�A��Y,	Q�8v���+|�*�"1���'�U�R�����C3$rQə.h$�2�N��q>[L3"����� o�3�Gئ��ꕷ��@��4lU��խF�D�T] �oIe1� <�
�n���|���@F6�sIrO�7-8U�6'�xF�#��sE�[n�!���r�����g�d�w��\����$b�M�kY��DmD�	�Zx�8�i����D2=�����-�����ՍkeJ�V ?�ј�
�0O憵�B��K�gÛ'���瘊i�� �eZ� � �)E�*R��5�Ф �jJ$���żY(��_#ҍ�����iv��5#����+ߺ����2&��+�o�!E�Bw���sͮ�Y(̠��_���-�EݣS��+/��8�u��X���r�\�� p�%f7��^�f��0�?¨����.DJDE�ا̳_�7*�z}�i��A-ʲ0	��*�ee��.�a�~S(�
��m��q������߰�:t$&����*B��)0�+Ԓ'��0�z�7�K#&H_���Х�O����}2�хUQ����ɥ�5��:^D���1Ͻ��P=b,��y(��l��n�{�4,�8�eAO��/󌎃�nvx� �f��e���V��LVRi�	(O�!,1S���c���"5Nb�@}��� ~x	"����7j2�f�2&�u闧�����&s�����f8�6r�H�&$�~�� �qUJ~IG�:~ђ��B����?�eh��A���g��=�7:�9���	�r�flʕ���<��k�L84tm8�O�Cs;�GԔ�N�F�;'���яHS�A�6��M5�5sUU
����ށ-&���Rg]��R"	��r:,��6�Y5|���Y��]���\:��z�1���ؓ�)K��
�	B���*젞h+|�76ܲ	�cX��/�aJ���з�`�/� �7=`�<�1(9�����%|�m�o�뷋ѲY�1��8�>�k}�0��?/gO'�Zn��� ��+H��^l��ڌ�l�h�ȂB[l�ؼq1(�x����m�0G��l$Sa�sJ����5b��d�p��cL����J��&(ٺ��Y��T� ���;��QQG�r8mO~��,�3�q*�?o�wNOYh�&g��GдK}�|i�Je�1�s��0|�ۡ]�㝐�>g���d���G���V:Fb�	H3x�M�i�3jCԟlB����������xI��\�ra`��qo_����3ڇ��@�`O 5�pc'��S�DCW�Q��p5�
C����E���q
��DW�ȣ���!K���R�H�`G�T���r	"��Xߪ���ۓ��EZHstas+Ncn����N^��� yn,�*z��(��d��L'` �Mq��s�b���v:� Y���_Ӓol~v>���݇��IZ<��7����ɢ�ɂ������N��B���cq� �ڷs1�_�bA�]�Uk��hsYJe�LQT焍6�܋'B��{��A1j�}�7'9ה����BQ��� gѸ�@C�3�+�/ 4-������ 䫽1��8S��� 	��8OS�����M>�H3����N3�g�ߚ�s��j.���S�����j���-��2o����)fܳ` �P�޹��O�D�t�D�̆�ށ���/�����ػۿZ�)6=r()�oȰ�r�U��v�,�����yy��N��ރ�}/����*
����z0uɺ���N���yN�J<����ZN6j��<�28B���sTu�[ef�^�I�)_02�~���&H���^�.YĿ���RZ;�J)��<�����ּ�����A�����cm����^3��(��N�U���}z~�V�WƗ��S�M�R%�id�-(�S�rDe����@S���D�=�p-(AW�FR�WQ�R̲�esmJ�l�1f%���Ң�c��x�vW9JE*YU�\/!�c��|>�8\:
I�ٍLrw#P�7 rkW�}=Q�[_���(�qX�25�	�;�w����r�n�Ζ1�E��L�pu����.Y-����v!�?���B�)�9�yƣ2����u(\�X����r8����T�V �h���������/���l�K��x��Bݡ���לgf~w�@�g6��n �13���l��9�F�7 /j�̏��*��-�{���ZlP�(K��Q�������"�$�|�}���U�}t���R]�_ʪ>�ÀY�9#Ɔ�?[/�<G}V��)�C9�ۛD1��%�f�̑���0���
�2xEYSm��,������&�����ħ���T+�"#_� |ʋ�5�V(G�o�ߟ��!��HNNAn�m�'�=� Xr���P�K��y�8�.\{�q$�0�����ʜG��^Ĭ��B;��������4V��t�s���G*��)���g�o��i|��^�rE/ Qe��So.@]�cH��x��� ��A��1(c�qP-wS����P��"���|7^6�$�a ܨ-X������uA{�=o�V�!}��o�.O��[+'��7$X�WǨ�C��v�c ����y��W���nu���$:�'E��G	h�|$�Y�˸�-ūu%0Ђ֥�L�<��8�N��}�o�hP۳Ui����=,33T�~H+a�F��&�+�H	����r�Z���'q{����~��B�c7��˛Y�W�>꿼�p�1����*|��F���&�fnm-�aG�s#�l�j����iW�)�w��rѣ�x�'���,��)�N+�A��6U�K�1��=1�bʀ����>l��~���j�[�
�YF��S��Әz�	vp�R�������Ѯ�p6 �$�����!�����0�����ȉ���!�A�MNl#?�c<���ڃ�k��{��̶%���`��'Ǣ	��J,h]�v\�s��P��>��9~p�O@��O_�$�Lj4L�s�3$6��OsA ��+��@�7�j�� ��W2��c��%pWO��Ls�0�3�Rfmw߷ٳ��#�i!��L���mDE��F<�sm�DN���#^�+�|cog��G*ug��w�^�j��F���V�t#���
t�KL��f��kP#P�5�e3TI���RUlސ~6��� ����5��K�����D��G7�a^�r�x�~�5%���3�i�-c`���t��%o�̠I���x�!������+6�+1��B%-��w@�(W�?��;c���<h18༕�V[ZpH*N�4�lx��Y�9Xv�D�iV@3m~B���;� �B�&P�V�@{`�^դm�8�Bbqv=<_��`�e�2�NZ˷7��N�}��0t7�]�A>�XZ}I�9*�)�# ���O��_��2�f)�'��jd�+8�I8�M'#]k���Z/5�?e^�H������9mɗ7�/�G����fh]Lo�	�9;�pz2k*"��h�_���g�V~(�����(�����Q&�}��M8�'��voZ��߆,yThh$�}l�P�k� ������5n�qd�h��K��j(�i�O�7Y'7uU2����B+'f���l��6:9	"+Vk��Kʦ��}V������~��ܻ�AMEqt�����rFT�zBu��*�EP�2<��пF܆���n��i�'��v��gb�d�{L����d���rWZ�rT/JN���˛S��$)s��c]�����>�ݷ܉i�˾��.�d�կ��n�Ҙ����
�إ�t �A�i�B;�x�"�n�z��2���y�����6�*��,�R�ܛCcٔ+G�� o�*C�����e���be�zF��TFÀ��R&�J/�j'�|���Y���c�� ;YPW�q���_�?x
����o�W�6&<��^*���p͏����=�|���i���vP
BrY��Ѡ��g�ިOi{��&Ĥ>p�l-�K��k����9��(�.�'�=u h���B*]��Sݹ��5-���2<��08䪈z�[�/��g�;�=��)Dި���4�[��N?�ћ��hq�~j	�E!�Dhx��G� �(P�L��e��3Ezlhx�4����c�-��1!�{ӓ�8MZ��K���/�D��g����[����6[ST�@,�i؊�KhQ�E�VU�� �%}�v���*l~%���'�f�C�X�2��ݲ8@�Z%�exT���0F�kF*Y]�eq�6zj�>7��2����t���k�v�H�҉{�`)"G��?�O�ŲR�(�.c����
h���fy��r?Ŵ��}!V���X���ԅ���֣���N����b�=�eH����#|��qj6����
s�z�}��8
#ZH�����N�F�N�t���b�0��i���" ����-g�I����S��?x�{KH����7^�|Oe�\�)��6��S���F<��}:n^�3U�c���+���J��?��4ڌz��<uA'�ųM\���K^'RNNh ���N/�,�u��I%�g�*���VGV,��o���Lj�o7�>����+Ep��h�<��5'�M����la����?C�[���Ml�8���>�H"	�H�rn��k��K�H��\8弜�u&	���!�4��囜׎�ۯ��TP����]���A���i	*$p�a@U���ԧ��u�o�z��&q����"�%�+���X�(Ǻ|pw�f�SN%�V�աP�6��Mw�-�fyp��l#��~�+����cX<�ߘ
Z��3g��r�5� �Ia�a���oУ����[�t��Џ�	2v�ҩ��B*'|�e��hD��
�+u�=7�7��3_m#���>o��E�þ�:gr����
������Fl�V��kI�G�d��y.�5#��L�<F���D�*��W����2<�V"��_=$y��O����	�zL�� xj��>[��²���n5v�p�n~D� }~c���8S �bW��A�m�Wn��]kd�"f]r�T�E����� ��f�i�_|ִ
�ҋ�DXJ�N�Tc�:�1Nb}�(��a���A�L�	W�p?�E_��T3�����К��\�#y# ���ERm�P >P.�5ѷ�A�����zAtMÍ��o�!�h��JS<��@�����T��`2�Ds�����v_��
����h�vI);��a�v����}�\����/D]wQ��bw�
���7~ۨ��|��e�xr$��0��?��3�3�Wʕ�{t��T-��5๗� H��.e�Wv��Xm���*Ym��y��$`��5q�|^��� ^�����ʶ�C�QM�"@�A�JL��9�[�õ�DK9'�a��ll�����/�+���(z��רW�w�Ũ�9J���1��Cӫ��,M�7:�)���bֶ]=��S�����G�-��.�����m�-�MЪ�Y�a����N�9w�Z�1]%�2��@���]��M$r��#t����ِvvŠ)�p۶�&������:�{%���\�
���6t��(D>�V���e�2ҩ�b�6e��w���c
9_�`'�9�r4�����xx�N�	�����8�$?Q���e�E�^Zo�q8/J�ƌ+���!ⱽ/�
g逥m�Pmܛ)��%�2u#��A�������
/ �p\k�[�?�(uѴ�>���z� b�a)T�Ф(�¡��p�f�}.�5H�`!Rc�w�!�Ng�\4Vm�g[�nwL�מ�&(��3wM2�{ӅW�베!,x��~I���6�|S�P�v���hh�m���.Y8�vCy��
��!��ݦk�v^|�K�ҐFW,
�"�m �,+n�Ǜ5#�v#kk������dQhy@3�N��Z�ӛ�NI�53���p�R�P����t�M�x����m&⇴��
=K�O��Z�详���#Q�;΃�V0�^��cZ���͍f�V��Cy���n��<>�(%rn�>�l��M�o'�GlL��s��BD���?�
�Oۗ�3[��4��vЇ*�*>���wτ��@�{�7OC�]��F�����%*��A�kdHx����bUJl�r�}}��'IŅ���i���A/���%S��n�v�$1^����3{ړT��e̊׌�����5�cJ\g��"�A��@�������ʦPAĮ#Z�H�I����rۂ��N��`�5�Z���\�K�ʹ�]��u3���%�	�e.�e1�n/��2���X�?�?�I�C�6*-	���Ƹ u���,N�9���NJ���7ܣp�j �������4�ˮ̗�{StYɏ�7�f�˭!Pk��������I��Z��#�xlM�!s��t}���tg�GW�
�|��0*l�M��H����E3�yq=1K��'Q>Wq��D�$v�vs���V�X �^�SN/a�O�_~2oչ�R�J9�6=�x�GI�]M�D�%���Ij�	��C����[�Mh�!�'�z��^e��>�}��fZ֔��X����(�gk���3n�����~>b�,2�\Me���#�c���8�^�AOI�0���u 8��:�����ձ�è����	�0�Ł�=[������=��NTR�tCmf�FA��v�6���{������t��\cHx*ުX���B����s���m��{yw���RJ������(�Q��ZnӜ����V�a��՝��^�<Z>	B�>�H�x���ֺ�AbT���'��ǯ6|~CSg�ϥ��6:Ѳ
mvIfT��y��N�B9D���=j#���Q�ovޢ_��Ξ�����w��+�~gN�Ĳ���>m�&����ܐ-������������/�;����`��"���N�����q� �rZ�
2��C�c���*���HE,C���%m$�|�]��2g�����YN�9[�y�*)u᭖��R���>fk�����r��%T��-����<4��P�K�ߪ����'RԤ�>�W��x$c��}��Y㖆q�ix5WD����$I ��5�����@�����(Nt����Rtp0���,��u«�D��x��x�dL7����W�룶Jy<}"kޚ
�^z}�:�&�']Bp{�!]����b��Ŏ�A'C�D������g`�C%QH!+� 5����$AL�� �t뱇���0J+��4α�酥��0��߃\m�8��  ����4%QC�C��b7`D0�$��g�^��1
�T���o�n{��/��U��o"A�K
��{��2��r�K{E�-��xx/3�"����ݨ�[M�p���\�h���������(s�N�::j��"2f���-9�m U������lfǚ��DR��_�k���
��"�ՋX/�o(�5Ңi�f6��E�c�aȒt����S1��l:~�����7�TC�ж@u�g�2�n6�����Ώ4{p�]Gm�b�6���JW�4�h���_���z�L�
`fu��^��M�q�p������	������)�u����������|D���ь.�4	����~
��&{3n��Q��k�3��7��0�u��kK�aIZ"�=�D��;��ױ��7�^D��ʒ�(��(���Ѫ@�����O��s�<x��9�&��#�i���D ���7�Px��4�D!����Ơh��4����B�? ���yqi��|��M�y���BEe��7�L�	����Y��a26�L��ba��4�P���V����!�2����{��ޘ�kz��H} f�ʴ�]W���RC���w��c�vd�������B� �|�>�U�9����%ʻ���ǯ>F��L��/���c�)����{�:"�z|Qe}]�"xW3M2�K ��J����e��(�R�b�jU�An�L�Fآ\.j��Ԗ�_���e����ɡ�-�B��@�����zf i���+nF���h�Y��.t����N�T���Y�2[�'�iL�5dW=$'$;*��]"����fv��F����9�����՝os����U��x"hh@�^!�Հ�5��\s�}Ff����p/��;*�DuzVУ�:=�0�w[�p�|7����f?Fŭ�Ơ��JJ	���	��{��/�����ҩ�}�O���>UX�S%e�z`���Kf�
�#�8�;Зos��_M�� �O�N�жd�c�O�������G�"B6G��v��=�дE:���ߛs���vJ\��U�́����(hݣ��qn���q��l�#��KL��9�����S�*"�J�'�����ǧJ�x1��dK��>9en��YZ��_?�L��y�����؅�������1n {���Y�`X��:H���������YTf\P��|�|4ςˎ������[U�Q��H0ٮS���+[�:�ZȽl�h�Zr�����o�d�҅����ƀ ,
��w�'����߾��E.��5+�X ��l
=%_X�0����p�z�YM��w#A��;�e�8\�;�	���������(܅�O���UF��>�˨<U_#��ȟ�Fb�בx�z0�ye�|3XFi�j��hС�f��^u'g���F`S����=NUvk�܅���aFojB-r���=���#��O���m�J}�t�'z�8��1�AN�u�B�p>��B|w��q{_�uٕ��rR�%�<�Ĳ˹P2ߢU�S@u�p
�o&\QQ3�?��(��p6�Xm|��M~���N���\���t��G/��ץ�R�?@]`�A���`�uie�t̰�Bꯐ�0>�C8ߝdS�#ґò��m���]�y}���iX���k7�C�tb.?�.����8���1�#W�c���bu3�!�]������8���4 �:�7h�7T�BUZ�.S�/��� �w��l¦��6��BH��NY��N �{���F��-��'�{��?�9#��p���9uP�yb�Q�"���J�va�z�%�dG���Sw���(�%BЭ7K����{�N�.�)z�m#�#�@�m��t�3�K����h+/����LGN$U�Fv�]l͝j\�#�J�ј�.�@$��:�c(,"���K��q�Há�@�_8{W �pGc-��e�������e��amSM5�G
�͍�oQ�����0��0��.����r��o�9�k��O��CX��n�K}��.�2���i�3��ɟI�.G�|�gC��o|49=ƌ3�Ãb�rU ���p�[k��t-�ɞ#ߔ�����?���K���S�أ|Ak���O�h0r��5U�kI�i�B�(�gs,�S�� ����9���Z��}����R�3;�g��;e��H��4����=�sk��4ٷEv�Lc�L�����1�����P1sJC��sk��y�u���W����(G���>�D>�o���!OI:�)
/��5A|u��n%c���"��RN�G/�5���YI�K�yZ�m<�k~H�Ƣ�����{8?/u�m��]�f[k��^{�)Ep�e�����ax��wռP�\ظ~�~BRs�v��ݬ��}�@�'��M\`��)A9&%>���G�R����y����M�[A��Š-��r��zR�������e.��G�����5(�d+9F�>�8��2� ��q��}�ے|�m`<ąAdCJ��*= 6A�����ڼ���
�! r��PNB�RZn>����T\��^�\��,�@ݔ���ȗ��e�~��0J��(Sz|Ι�nu��1k��X�_v�x�`�;�kk��[�G��YA.���6�ry2��=<B�[=����*Ґ���s�ڊf��8��?'�9
0YM@�8� �a�*�����Y�΀��g=������TQ� � ��,7�z
g19+<W	piu��p%�n~'�kvƕS�g�Cp� �z^�OJ��j���DU��Z��b��t`e�}��)>�
u��S{I�-_XVr��c�A��&b�d�	�c8�����V�89Uq����w��q�e1��Ա�^{,<�h� ��C�Шz��,T<s���yx�\A:"])�j&Db񥽴F^*e�}� �C���i�}�M`�bXJ-\DMH-!������8�h�l�� Y�е�z�n���
������[�+��G�y񜜖��;���nj}�r��X ���ןx�O��F��_�W[�,�l�������W�u��,<h�H���|�>�R��������r��&��}Q�L�yR8��m!�4��f���j���9<�R����,7穭(Ҭ�T�G\�O��>̥Gj�0�zM��&�%5
{������飂����Cf1���3E.�	 �"��_�K!��V��[�U R�G���p���1c�{�n�B��YM<$0�.�B�p����k�� ��o�� ���I�Ƿ9�[�RS'��^<(;EShdy�ɂ��^(iݗQ��R]���3�O����`X����A>aVj"��d;�D^���'�$�Ϯ��k�o(O7oN���l'4*K:2�]�	?�7����[%Nf�hzײ
;V����x3���Ј����,�T�a�� W�|��>�3�3���柝C+�1_�`󵾶Զ��3�=r

ߐ�Kzhu�H���b=m�][ӾQ.D�Ƨ��,�$�A��6�,�e1z��?��ǁ�X��q�B�����E��BY�yj�H��۔���I^�ڝvd�&���p���	IL|l�ލ��tx�`�\|�
/n%aX�����+ޮ������-Q����x�%	�f,ߔ5�s롊�a�vT�ێkP�7�╢�qӹ��)�)�����Oe�x~=�Ź��Ŀ6�&ԅ_��_�f2x.X��L����MbRV�=?i��+�,�]���9c"�tE^*~����2ƌ'0��q�P[��4���6�uvnF秳_;��9䇒Đ��BkM�c?�¢���?�Ÿ�x2p,)�C w̐��"cI��mBq�!��*�)�#�����~��4E���v�>�u��ph��̲Tqy��i8����I�p�.�(p�t}�H�V����PSq ����~/�$�W�����ɠ*��ϦG�i�5G�j2���zcX����1����ldf���݀$�=�_��;*(�pZ��s�ߴ��󇧚4��ofu�M��wj��UNeg�d���vU#�I~Vd8WL8�����Ƚ��Tg��V�Ŧ�E��*~2�vt�0����T����=�+�#T�w���sFX�PIw���	����4�:��L��������*q�4u�2�Ǳ��#C�T�b�/I6щX�����m���v���X���I�1����Q='��{���E����-�A]�F=��t	��W��Ɗ��_w�&��>m��<P��Y&�Y ���ʶ>�ME9*��� ���"6�'e+Җ3��_	�����GfI+�tc@��<�I9�~X��k:,��F�\��_�1e�����a��+�AS�`'v�[.k��6��W3��u9����	.A��U�ld&�=�P��0�bz�"z�c���ύ��oPbaiC �M�����#�����_q��Ҭ~��U�7���I�YMi��X�J�Ş4eh.q�sUޖx.�#{2�Ƥ(]�OQ3D�`��dN���_�D�#$����~C�d����:m�u(,����Y�Zi�Q^��5�{���Fx��J�E��屉b�%!ƈ�3�\�=�l�#RIsVѪ��R�FL��o�#ak�_j�ɹ7Z,�D���H���wqf���?
���^���F����zNC����o�w.ʠ�	`�=�)R9r�f߷Kp�l8���^�b���o��*� J��c���^�ZG�$ ��x���K�>�͞�aRS��?], �=y���i�PC�J~��tp�� �3��I׸��~�LA�˃9�M9W"��͏#���-M���@'�1�������5:'#O�a��ܳY������k�[�D�)v~�3�n��轣�@{���$�4S��#w������A�:��Kq������A���F���@R��ǑW3;��m����

k�E���̅��^�gc���h@\��4P<��Vr)Vp�.����y7����Q�Bρ���Q�K����nol=1�ۂh��W��З/��n���b�&���� ��Mm�0�m�������״���\�dBM���3q��SL�?���jU�k+uj��S�aQG�t�V�(j�&�oN�d�y�ٰ./���R���i�� 䢴��%U��y��e�ޡ9�.�;l��+�.ɝn5P��j�>!�@.���Ay3�<]r��z>
�t-��r�H�f"wC_<~���*q�lL���t	` ��ܞ����C>I����~���h���e��#[��%�(gd[7�df`[{f7�1?�e J1s�Y���N�����%�.D0���;�[,(s�*����һ}�Hҟ�qU�zG�3Ռ�_Ɠ�+κ`7 [��#fF�=�H��PR���GpGQx�;$�=�ǥ�M��H��ێ�ř�{����7:P��7]
�aǃ��{�<?��^3�aE3�W�kw/�����e� ��g�qB/�[+0�u@W�|��dj�&y���QG�&�@Y�q�K���˰��|�-߮
4Fk7|?p��U�P�Z���9�ʦ&]�8���s�>�C����x�ҝ��ȵZ}_�Pe��$K�9���];8bnw�L�q|�o���'�����w ���dh�?	�.F/	y���6OY%e��$N���G�\� 1�z���k��XW�n<L�,����c�@v݇�Bnq�/<�>�<�����6%bE���~��
�w��џү�X.x-VS�U�DRY�f���3F�?��^,�5�趋�N�/�V��	�4�����^��vxR����@��K�K
���H$�{�a�+z�n�f�d��R����?ߧ2T�v�	za��X��?���K��8�x��xO���w6��	R�h��������/ul�7�cx.� ��7�V���'�'@�I�Ŗ�/�����Rvnx�0�1`R�I�>	ؠ�#O���9��#7)�N��ꃓ������m�y��?�1�G�·Ņ���]����ROT�z��T��<"E�z͛�K\e�ek�t�@���6s]z�2E���ĦNYP��z�����BK���+ɻt8�� T=�m_������/��x�F�lՁ����7#F�������EA�X �>���84��3���Xm�B)Sno�������K�%�G�a��N3��(�
�$�K�:��x4�E�����&0KR��B��5�fj�qC<�Ў�&uf���q\�F	W�@x����#�rj$j��[&�gty�Ȑ�<��ʼ��������I-�����ʇT��ke��%+4^�d�64.Sa��;V��Y����ٓ�o���t)X' ��
I�����欘@m%���P�� Iˍz�i{���Gs*zC�4|��Y�NQ9���x������V{�ȅ��Fݫj&�����P�������H们pm����҂/�9"����f�� ��%j�'Q��x��/ɤ��*�uz�.��u#��T��w��h�T����"�("z�=oW���־-J!o�RY�R�xvc_q�r���՗z��Z��M�B�%;>�Ep��dq�����QX%��`�&��y�<s-io�4mT���b��YQ�i3����GY�c�kS��,<x#34�O-{G�]>l��%e��,�2vX�.�����Lo�vns"�[5V�������y.2vq����� ���6����5��P������fq���<���1LQ��V2&����!,����5q��g�ռQvMy���s薌����YZ�����ƌ�����B�y�A���I��	�>��=p��B�e�b��Н�:�1x�0c4g+�
�� L�Q���h�q�u�J���D���Kۡ:�"� Z�͜ڼ4G�!��ZA�&�R���Q�����1�Ӳ�y�2���N|f�-�\��z^%��x�Ѵ�%��Y^%#����ʌ�'�m|����PNh�M��q������4蘕n`[QIg�(,�ތBM�΁v� ��K.`�Jrɻ,̘i�ɶ�R���ڂr���Ȁ�]�8�7�.S�ϻ~a����dM��bn�Kx
�~c�����D��~��}����,�?�@CL�CA�W�];oO�S�(��@^z�F�� ���fxM�uWG&�v�"���L�Y�,/�>�������6�; K���5A,ZT�\�dyy������I6����53`����)(~g��B�
g�{[����d���a�t��xy(Χv���j(Js:o�[�)�HE�����k@����h0�ŭSC!i~��+��zPj4FR�/P����k6_ L��b`�/��t#]��6����疱�l��z��<ov�@r����/kZ�C�D6m�_0M�X����`�h�l�����p�%!{����w���qK�w�A��%��A��%M���.cO4qj�+��Xܭ$�.·�G��}3Reqh.]�G���-���4���]��@L��X�Q�UwO0tQ4�;��G\4����^p=%B�ԕ[��~�b��Ip����m������h%m+ښ�͋�(��u+��[���)cwh���H���m��A�n}$"����bD��}#66�I�r6�ܿk��k�iK�^�hN%H^a!['��[ޞW[�ߺ����z���<���f���V����o\{d�b����e	tO�MK5��2�a����qg�)��J��F����7Ο��]�ڿ�$��t`C;���>��\��8�@��ĳ�F謲"ςڦ_ՠ�e�t�T0͂�}R�~�C0�Ug�`����/��a2���N��>Xj��p�K7��Zz�jC��h���;�����1���"C$��l��0<�4�����rR�Պ��[�Do�G%��}�N&��mL���ӳ�Av�Os@fMRI�8��*+|��guâ� {ު�`��\�a��)��E`}e�.�����-�7��Ն�K4W[N%ڡH{M�ċ@6�p%�B<#N���P���Gu�!3퉺 � ���El͌R�欸�Z��ƕїE*7�uk�7�jA/�1�kmSR����8cL�?̃��F��+4�F����}������v7��+��=O�.t��1���+Ң�ɺN�GfժE�5��DQU
�y�T�"lrr�J#@���Mç�|�<,�%/9� 6(���{��K���p���$��wΫ�I�	V�M�!�U��L���F�2�m�.�bc�Y�*n
a�4<�n�׿�i��H��k��l,R�,P\��G��If`�4ʕ�fӠ�|�'��@mj\������*᳥[muI�,w=�<���V;�:<ud:�|�GQĕ�ҷ~�I�n�f����E�kKҸ=���7R�+qfrQ:ps�V���f�PUE1n�]*��Q��o*�C�2I}�B�d�^�I�ˤZ6΀;�}�^����&~ȑ=M�����QJ�"�_3�[�l����)ɐ�)j�GA�홨�t<c.!�m=Jn>*�"������̟]�ET'�M�3��y:6v�Z�c��7�&;'ў+�^�<.a�O$`�0�ze� ��q_Ч����b�cH�S�Jt�{_�V�:(&8-��G,m���#-����C�S���5O$�F�H嵪e�F'��p��t�ϊI�uy,�y�@��p~(N�נMx�ܛӀ����n�wum��MIbJy��$TJX	���y˰�A ��	�	�Y�\��%��֮��2���h(t��=�����I����;�!�c<��|�����$��>���(�]&�E��8�	�����w�L;��ê��j}��oǬB7s� ܯ�A���|5�3����$88�n.ɰS-����^ �������?�3��4�X��d2٨�c7���Կ���IQ4���!�:pJ�w0��ѹj��x��п�j�C��f4�rKN�ځ����+F�Z.�S�M���"Dn/��J-��:\�{�^4S3�F5����;h�W9o���6�`�pݛ�q�*��8�6s����2���/�d �e����xNz\�.��-�<g��u���ű��]�3�י������+��~���8�57�JL�M�U���ᲃ;��':A`��� B=���u:�&�VD[h��⅋F��Y����H�ڗ$�[��j� 	Wp�5�E���!,M��ܪ�\��������8�o��)�6���d�8o�I"���@a�ǆ�<���;���Y-Њ��{�;��J�L�C��Ztj =Wɽ ��{$jL=!�WA_�e������ �m�$t,v�)LOm�� j|HN����Ϻ�5xZs�v�����O;�W.�͒����Er�h8uH���jB>����`+E�w*�p�ܗ�ZL��|�4�n5��ݱ{���#�Tv��Ʈ�u����#nd�9{����
�l�i��80i�>�;�5E"��(8���?�L��OUV��U�5����`�;C�R�G7��*b��~�,7�q=g�����N����ł����V&-�@�5�
��o�=�gxl��\���hg�1|�W�O��GȆWǦ)2ho=t��y���G��U�w~�Q��K3q 6�m|s���љz�g����>��#Å:B <�� ���[?��o:T<dP��2�-Wk������wG���6�j�?NH�2{����}���ʗ���+(��?��出}���c�L�@o�4��jN�N't�=��<
�r�zA�`�8~�6�A��/��+�E�T������6�v^(+?<ŏ�pϴ�4�ӏ�eJ@�p���<<�,�ˣ�;���q.��XY��U�磦&��Y���M;X=1&�K����p+�F�`��|97���N�A�8]��C��^tW��\>�4�Y}Ծ"@�,CDbR/��wԾ��b�1�)z�,��"h�J�JNB�Y��W�Q\��Cm��o8K3���|v+�K�.���ۧ1	�m�v2�[�r5�rC}ͳ�	f=�$=�0x���gR��!�ת�a��.y}]�r���2��r���/d,g6��u�K�'8���:ejzZ�6d3�%�<�ed��]��ZBPD�<8���!5i�صf����1���Ksj�+U�%8��(�g�)6)�/Iy5������&`PYyK�ap<52��4�Q�;y��� �@�Aߋ�+����5�`��6�#�Wԙ���=D�r��q�-�CNa	��_�j��W��BYX�
]��������=tV!�t��+��׆�M^Qq]Z=孃���o��g��(�۹�W~��K o҈����L���4�3��� �!��Ҫ�j�NJ��9�퐋(���M�JS���*��x��6�S՗�+�#��v�	?.�E���p��'�1͈9Ħ_08�=��,٫�7�j�n�[��x�@iGI^���y=�+.��!�`\�b4]�Пߥ��=�vJ�?�{)d�R�b�Q$��r��]�Sa����XH[�?J���C�Z���}�1GN�p���d_�v�j��m�3�|�`��x���[�V�����5nQ��=�����:\8�G�*���q��n������^:�O%NTMT�Ł�=�7�Q��o��C��8�0�={���a�q����8�W���L� P���C�&�u�S!��DD0
"�.�A�[0m����_����L�ro^�2ƾ�[&5���7�9*��n��Cd�3Kt��Om#��Grq�4%=�[?ѪN��b�ZΙ$ǳD��A����N���7�T7�_a��م?��5`���sr$��0�#�<�Bt�>`ec�����f���z�l_�L�_1�����.�^K�v֝�9�(�+�������L�� Qaj��NM2�b�}V�y%R�x�\�JB,�Y�SJj^Pȵ�f�KklX��I(��X�Z��� ��)!��	z5S'0xn;cp�\Qd���� ���D��Hy�|��-܂��L��l����P]^d�#�F�o�qLJ�(�Y��aB��}^��nSC�Յ�GS�ݺ}H�>'h�/�Z��V�ɚ���n�t������
:]�6Q���`�rO�ˋ�J�����`�O�Q�_>�J�`��b`l��8���>�6SW�V?��0t���8�8 $<	�W+e�Ʌn	�`7���Y����G�m�{�7b"t��D��[n7�?(�m%��TW�Q�-m.,s�'<�Οǫq������Ƀ�U�!�JD�e�k����X�
�����"0�����m���j��������Fݎ�`����8��vJ\7H)I?o8����������Y�����Bm�љV��. ���א�^��֯ق���ڕL���d�/i�"Ν�J���à�vhA�@ש9�˫P;(eH���枂��S�6��*9|�w�o�Y�� ��\�R���M	�\��n �-��ɍ��"�#(z�k9 �c1�	�(�R�_#�G5-.�A�:p2��F�� ���񜍒<�v͚q�P���i��kj��G�r�Ǜ���:6�8�!
�}��CG�����Kܘ�'�:{�,��J�N��a��w�-�R���F�O}��n��9�I�C��ϱn�K%1_�ɽ�n�c4��+��~��e�����2҄��+�4���x�7�$��y�`Q\�w-�Q�m��v���i�x�%������ꕼ�����T+�s�+4Sj�P>~�ސ�������v��� ���
(��������>� �?=�۵���%��ƛl�)����GjR ��t�d��E�+6���W�I����ryp-�<��;�b����d3�#]���W�l����� �]t˼�V�j���J ��\�T�������|�hX#�q�4�6H#1N�x�H��HoW��j�,N�2�X�R��*�7��=  Z�.�MN����V�˖���^Q��>�S��.�P��<�:ԍ��kGhfڍyszL��$��ҡ&���TC������kT�1|��p����)��Qc���U\�?����-��4�Dq��\!�d])�K�C�fƳ,�O1���[�U�(��xª���ӄ<z<`��&8�%�R�e_jA��H�8�G�b�����y�otj��u�gE���7���j�z�u`X���.�D|��\��!p�s�˰�� �O�>Ƣo&N0�������[JF��A��|`�/Nƥ$��P�"$}3@�U6���W� �b؎�֐���(���^>�ժ�Ǫ�3���y�:q��Xs�a�c�/x&Gf3E���B�ӅYZ�e�d����4�<������Wp�@BC,A���oӘ���FY�Jb�4xfu>��B0�����7����c_�I��Ϛ�m}%
�<�������> �i�'|k"p�ϑ��_��=�D'�nq��2Rŀ'NRHy�Ȋf�>z�d�c�D���~��غe�������,��ZM��u2�hr��z��=�a$.���t��B.�}�զ��;��yPL��=����t�-�
�����ar/�Eò"���OZ1L?���\Q���w�*�?)c$�{� U��s[v�A���1x��O��ިI����$������q�c֎�?���D��#덁�a.��tW��R������4C��"����96�&���ʺrU*�a��/��C�viJ<d�+dl�{W�o{��G������lS��H�@�"M���/w���I�[�αSx���m��$k{`��ƲOv�������
Z@�QY�a�:j��}&�[htp����)_d�#G]t��>7���4���8p!�W�� �b���Wǋ��ͽ���8]NԷ����c�'�2۴��!�Syv~gB��fô���'����SW���peg� q�MA9u5H���G�Pb5~־�G��H|�۫�N?���Y�[��,h�d9 2Nذ�Etwo���A{�Z���Ɇ���B�U�������gavPM��|�P���W�u�٘g����ּp�Ɓ�Ɇ��m͡	�]����~�I�/2���C�ϔ��Z��}��4��Xh菏W�����j܃�2��|���8�1�)Ȫ�(Q��1	^ 93�kЪyq�-K����i�#F���^�H�f������j�R6�&ִ�'ׅU���+��K.LH���k)�k��_xH��.uIoI�=?�8" *9+���y*�O,��*��T�p� ֮��gh�U�Z>{z�ߦF]��Y{��W��(��Sh[�y�����OV��9}�e������)�зqY��q����#=�`��h�j�V!B�p-a/�x��/שٌ�����ڸ��jt�TyD�+�6e,�:$&�楍2�q-7�.O�d�U{~�_K��o6w,�B;�;
���F�}p[�C\�L/�c�Pń���zQ�6��J��+ԛ�8kc�6�ӷd�j2�lӎ�L`�}!���^�L��}>v�,Lѿ�W� �Sv�G�IW< R���Mȭ1�����,��� H�F�h-�9M��8��L���ŷmT(�T�K�g�p��,V[�
�[�5(qB��rF�����`�a߬;�̺�L�������'���Q+Ϫ!� ��AJ��F�!F��&0dU?=
��S�/��G��M΁��Ŧ	Z�F5��nq֟`�o��������˕������,��@|/�۲�7u���})�{`����޷x��@Hߑ�"q?N}%F��=�Uy���:�R��=���v��qX�@����2 %��;�t���G4lo��~�d�C�2v����PfEq�7�u���*�V�� 8?~W�t.��dԦ�E-�� �y�HeOYt�����]�LxC�.������T��hi�M�ut��4hU�]pl�ŏ�.<ݧ%?OG�YB��QaX�)h�
m��=.�%/����!���p��a0K���^��A�A�[ L���Q�}Af����8���ڗ9�B]U�(F`�P��N�=�9�6�t�a h���5�(�(���#ཟB���HGo@;Z`�)���o~[�.�Y�T��'t������J��i�i�/��,/d�Hc+�_��<��MY��.�jz��A���z����ؤ�w)GI(�c�k#Q$�Ma�������YT@����g�H%0G6~{�V��-09�	}K��K�gQu�E/K_�8?d	<>� ���&W0X��r��2iR�a*�@�$YS奡D�rWG�1�}�C���l'�������l�}�O�ǖ�Q��}N�.�Bi���Z�z������]�k��m^��$ a|�x0���cB���'�3Rw�ygy�>g;\�.T+|&�B��x?1=w�`F���ĊH�q3��VYI���Գ�k���Cd�� ���E�:������8�xk>���FR)��0И�'r��?��B	4�`lq��| A��ҷO֐"�52���~^�:������پ=`XN�-�#�쥠����@J���m
�\Ix���1�o�ܴ�ú��C=�4�\1J*�0�I/ްz�B���gM�	o���2
dȇZ��U�4]��N�3������<�b�ɐ�pYc��ol%Q<A���
J�^x����1����#tA.�;��T��I�R��)�f<�.�8Aev4�T�<��ݠ=��T�d[d�+�ס��%K�����������֏~�bG�j���.}��,Q&��3dd�aUv��~�C{b���dx5[��l��T��w����_XG��|����m��J-m%hY�ܭ��C^��T�Da�J�荻B����V�D�0�Jbj��g�E�!��{(�a�oP�TB�����o��G-�s^�:#t�Ѣ�^�k�� -s��W$Zk̗^i��]}��xQ�Wưq��i��U5�>�ך��W$��.�_;��G�	��j"DzZ��@������0�Q
YWL�o3��D���K��\�����>�o�]��̰���c���/��kL���]�#��0��󜷶-�j.#�((�$33��{�ڸ@���L4��b2B�%8u�j"ž� �]q\�9J�i�O�`|V\%}4��~�6vG�K[?��h���~���|��Ӕ�+�
ť��$}�dE�������^����t�������ēv��h��/����4q �]��u�Tib����dǻ((GC����I?Ö��dRM�SI�Q�_���X���I�*XP���r��LPe�L���<�[[�r�5�0�&������G���?�;������w������"����c|��,n$Ӗws`�̻�/�Jgv�1��QxK5q9y��v���q��Vf��Aqڈ���A�J�d�L�⮵���4t��ِg���r�����t*�9���Z�i�]��~������1�25��qQ����pL�C��ų��U0#һ훮����I}�� �\�E�-��lR�T�s�8'��@�̽���R�2�W�ѥ�:���+�/�Kڤ�^w�!�E&E��Z�z�E�rX�{X%�b7M%�;�M�5|
�'�G�z��Q&$�C�W�n��vG�(�֤f��e� ޽��ҩ# ��A$٦V���<N�*l"��#��~Ȉw��rDߟ��}/��^K�3�Z9���R��c���gz ��'������CQD�}����d���i.�:pu$͈��e����^��,��zn6\T�,��lYB�g܉�����Ҽ��àT��_GY�rV/���Hv:`�9��@���ɿZ�m����5~��:��j_����cx�AZ\sK~`"���S$�8�W�<߇V�[�m��Ek4G���E�|<d�]z�f�M��6�v;�.SI9}X-p�1�Ampl�VoL��gf���x� �k���t�k]�v��/]�I��{�V��	�9�w����eJ�,JR��,\��>�i1ӑ�c҉m�\du��=Q��B��wH��VW�k�j$Y�:�d��˴Ӕ�9)�?���=8xH�Dc~���r�'���ʀ}Cν�4[_!��ȃpB��+�E�'��/�r����b<c6��.��O.���r�SLt)GQ���H&QL13����d�p��p2崼�K�HVq�^��&����w�&~�_��Ay��{2]Jm�iJ��(��SVIy���U�Js�3�A\�������yg��ڝp��Z>�t����VJ�5,��I�#8}9a���4U��}�nF��Qi��A\2��5"̛����i�JQϡNkb\M9X���P^2D�g� ��6S�!�/頡�	�8���bh��Qxz�0e�9��s���G�sYݷ�
�z�=�߈��g�`:|��e���u�|��i��3i?N!�R���w���(�d��\��`/p{:5�ݯx��+������^���ǩ�A��.>[���]����]w��s�Vn}����g7��� �+Cؘ�$�|�֚�"�9���q:i�H�~�v���ZP���«~¡Ũٮ��q|��Yi���Cb�u-�q"�����i��"�����ױ:�T����:ZV:f�C��Ղ�.X��sNo�Br��+j�(*4�2h��]�G�or=�������<{��q�Œ1G��3	��s�%��F�%g���1��4G���G��	wN:�l2�t%�c��*�I��2�D��[����i�;.Ik
 ���g
`��!'q�&�k��!�&{�� _�q5�gz'|=��Ü���~��[����!�}�%
?�)�yEA-�a/���\u�E��k���6m�[�͖nt��LuѬ��o޴�u���6^^D��g��Y�i�k�n(�S,�w
_^�j���v���8wja��$o�d��cps��K�W{ٻg��R�ļu-�L��qx�5?�J4ee!ku8�4�k��dXQ��d{�N�T�l���ǝ;m빠3j63V�����^�v�v�"\�.�ߜGN���R�F���K�
�U�/�?"�H��a��ş���1D8�?~C���Fx��p��O-zp��U��L#���'�N�ɘ���O"����7(��4���~�/�7�x�� �b��m�����m����ֱ���y�#8'�v/%����~�@ם��x�Ґ+@����[T��_g��V�:��2�*�6勸F�r�g]��O��׫d�
�1��|���q�d�o�)���"����=5r%h$�e���;�9K���ݤ�I��}Ahk��X3�_����r�(&\Yr棇����ls?�g��b�5�ΚZf�ǜ)n����(̕�eF`Jo�f���th�x���p<-���<��C��a8��B���ڇA3q}pJ�L�_,�eL��LNO�d�� �h�L����>���m���;wh�{����\L��%�p�qB��J��z)ߠ�<u�6�TK�5g��9;G@���0Ӧ�����q��"}z<"C��w=&-�̔KM����[�i�`���d�dd������,��o"p|�V����e��U�˥07��KGoI�V�q	�ے� d�7U���[椒\J���ɜ��:�0.�\��}���ۺ�Ȩ<��M,h��Y�w�^�y�.������w��.w�29f�Pp\�S�0Y��}e~Uד���ı�fKw�����][4-��5������ኗTF�z���]4����l�#0R�ۄ̊$.���$��!zh�gn��D���v�-�O��Rw�p3�;/�q�-��Ùoi�g7C�����YYs# WJƄ@��{�N�U�JJ㾘u�(�4�k��1��  ڄ�G�:/@�+_�H1��c4P��I��J���KӔ���O���r� 6��Pw�<yBm�Ք	�P���E����#5Pn��_�n�k�20��`���/3Q��)�ˮ!x�Vs��@����	j��p��P��~Ē�2�w���W��ᘠI���mS0@���8���8b�2S�%���W��GX
�=��/��"����j�&�g+�� �����5>��A�O������ �����v��Q��Ѱ�����0P%���}��P#xs�zW��׫�zu*}��Z�ݥ۫C��D�c����m�ɧի���܃�2�\*�8k�ƳL��Ժ�GD�������K��D��#�L���<�8yk>�~`��Wy�
x~g�g�����-���fM�)xLy�G����_��ƛ�x�����9��&���\I�������\pb�ҴE5w3x�d����~\�-�'���'Q�|���[)���������A�Q�%?KQ�^���z��*v=��́,��?q c67��0��I��9F-zZk�*�Y{Π�LS9-x�^1�nH�]�b
�ad6Ri-%wq_���<���=RuP�&�s|�����P���]=�H��kh��<d{��2/�v�%q6��1s<˲/B����)g-��Y�i·�޲u��\z0e!0;�A�^8((�U���	G���7\]tp���џ���"��
�V�FK� x����Xg���D3D)�DR�m����b��x�:*�;f�s+\�i1�� #�nù��U�P9�'AQ���+��Vʯ.#�(֠M�q|�p�x2'���(�H���,c�Z�
%T������������R&��9����v�l�KK}�'N	I��v�G�mj��}	r��V���Al���Hrس��[��l����y��,(����n�	9qv�0P����c����ƥiไ������mǈN���J�bbG
��� �&3;ky|%��.��OJ�̯N]" �����4ܠU�G�.� ��� G��V��`OS����SwW7N��$1�S��:��Rܚd��M���ⵓ��� ��������|���j���3�V����
<v�4ҠX�y�'����Ca�w��xPb�z�Se	D�ʀx�б����c�+U��c�k�����-K2��cΚ���|Ef�	������M-��&�Z���`8�M�$�(��k����E��﷒�r�<�l����!�kCc5�&���2OU��ƺŰ�8��Q�Lo(1��u�yx�o����/f}/�|'����۳����S�	����u7�+YS*b��^�3 	8|D��I��9\h��_JW΅[���p\��ڻ���}�����V�4�{�7m��Rèfe+�P�UҲy�o�L��~Ŏd�T���=J�y�����(6���H���kE��X|��(�>LN��,d�g�J�/��\kXV���)��p�]:[{��V������?Jkwl�+)�)�U��]���˔��oƱ�X���+����=�}lRe�e��KQ��N����[����q�����-�γit�����N�7r��\1c���O=��ϖ(��y١Y�J~��^e���L	
�k��ח9�a�lUA�/��x>$�#�q���mU��;O�}!�9-tT�N0X�a�$|�����CL�D�J"�:��C�Q�5�.T"�1�OR%�<N���H��P� =�/����2q0�'�Z5X��9)f�t]��d�H$[���U�UX�����PY��T-<���Q@����$h)��0[G�k~Y�����U�*��do½�2"Y꾄r���g���st�U��� X�6|Ac�����,��5E�Ock�|�%���T(�WD�9'�ib oKj�y?﹦p&����1V��/��H�,�O��g��N�Ը��MjFxU��;R���`�XL6��se[]$��8�i�3mY=�S�k0�-;�X�t�f��PXj���_k�s�T�`X8�s�7k�%V��oa��D��Us$�*
���3�SP��1#���<��Lf�J����r��Ԯ���a\@ 8�P=3�b�ڧ�X�&�:�Y�E"��w!�(�oҤ2&��{�_������HUԼ;C�b??�,����	�K��!�	Y?��c�h��?�����h*���%�%�.�a��cO�s,�ieO;��c���5�[���V�]��R���m,�i��%s{�s�3x�&�Hu_6�2g�Jxs�UX7������Mr�&�⫁�}LJz>�#��2M��x_wwM(�����c�zȔ)�� Ƭ��,�0������ʂ��f4D���Z�����<O�k���������� �L[��D��PN���Do�N�B�nkq
/��V	ߨ635%1ʤ�c����YV���j]N�n�T��.Luס��xe���r^0>��GL����gSu�֐7�mm_��8o�� ��v(����\������
���vKj�� �'�]���%�z��:���d����V��O[�k�BA�����'Q�M����+����r���je|��BE��l����U"	�D_�£�CO�L��wy���G�]�*�4Q�߅\��1
<nb��JEԥ?�����^gxg+�
�'�b{���p�&�'N k��O���x_��~�j#l	���5O{�t���	 a�ʽӲ��������A2�̿��5���&��R��1}[\�̛2�DMY�N�ߵb�0�j?:1C�q�Y;�tBP��1�Ikw�5�/W%�)��W{��tC�JU[6>��9l�L:w�Y_ ����>�\��o�\Ch�Zv��]�b^���"6*�]��Q�0�5{.�^�G	}߿o!��H���4�lA#D���E�#���v�]^9uMR��TѺ�ڳ�	ny����:��7.��u��s�{.��M���ң��A��Mb��<@D%yr�X���;+뜜$��!o7��@6!�H�N_gcF�4`�;��R՞�h�z�ۙ9Y��^;������9��Y%�Fdvs����kb��UьEg�6��H�1�K*9xTI5�=�k��-�A5r�5��
�$���������n���6\�'�x#a����@>s7b���ʧs�ь\~#)(�����@��idHcwgh.�������-���[�b�iP"�h������܅Ӊ;*���a�w৒X ��P�V7��^���仍�r���5P9��ն+#��Vʢ�T�����3Ķ�pS̈��O%�}C��kȂ�N6��}r�aD*�ҵ̓�%lT�'�[��)����-���Ց>Y�b��[��ҥړU�AO���f{��ٹ��#�x��y��P��LB�p-������i�.a�l[��/��O���D�d��E[l��y��) 2�o��+���I])�c��SVY>v�Fg��C5�:H�y6GHt�����ɲ��uOE,y޷#��JT���;!�.�L���
&��h��	�m�����Sn�{�e�������|�K	.b�T7�+[҈�ǎC9�E#|�=Ɖ3�%���.L;P��6��3��K0�p�ɩ�
��8 ��q���=�ۺ'Uf���W�3Nrf�Ȗ�|��M n����a��v��o�%�ӲQ7%7���	���g� ��jVM[G���O�&���]���#��������/��&t���X�)���/����5Y�&�ўf�S�q��s?m%��ҿ.���<,�1���Hudr�H?���J �Fr����^�p,�Q�z����-��8�v�&��U�;Ԥr��=*qfUw��7iOl�u�y[���K��_���h�[���[ƼYc�W�W�a����Ǟ]�(�@��&X@c������y�~f��(Q}d���[�Qݟ�e�Tt
�1V>b��a����k ����!\�Qܤ�!"#���|����7g�d�"��+-,��f�+���-"PI?{�?�flB��v|:�]�;�:;��fj+\l	�P�S
c"
6����0�lRtg�%t'F�����;�$YB��r /��q��=$#�G=�S6����"��Վ~�
tb��
�Ǧ��L<V$�#�t ��-M���e�]E|g�!m�c�sGL^�f1;ƍv�&�otU_���'�z^e? �Ճ`��J}�k黈oN��8�S�������U�ty�I���������KV�e���I�\+��L��@��A��d��ˡ���g!'*��oU��Q�R����nKiúZT�s/�y�B���;�$&�����Q�7�y����;�}���"0��sW���E�DA�� e�{1����j�9�/~�,Ტ��|Wb,�Њh��,+I^R��,�|~H�r���	��6L%`q�_>M]87K�h�((#M�M8�o~�b������]r�����)�8�\f,��B���"��w������)\����~N'�ދ�
���S6+���h�^�Z���2��V�ވ޻Vi�RȞ>#���ǂ��U��S4��d��Df�����Tca��[>�ޞ�(���ʡ��H�r��~e��3�E�=Uw���t#a�!�d09�V��
L�����_8֣�Z�����h���j�*��x��A�!�!�k�]���0��2Q���s�Պ��~ ������f+f:��>���׭N	 ^b���+�DԵܢ�$�DR0�(��tDM4[��Ui�E5�Ѕ�#wJO�X�!�vti��qH]����iJ�9x�l"�U]=��/<#1ɷ�Q9=�<�/����SL<k/�q��A�t����r	�<�"��.���3ho��[���:Q���U�3[�5>M]>؋�$�����TS��jE�I�ǣ���e�$a�
�V:��j�g����w���R˷�����r��X�q5/z�-�J�f�����ʢ0�	��9�"�3��ePV��+i��M�7�X2A�e6�?�±ޥ`�GhC���U���6�����K S��"�=f�	#�-/a�o�0�ks��mӈhr�����G'�rs���8V��\������{{hI���* n�դ�ic�+���o�\W>�=��m吇1�ok[2�E����x��Q
~ű����@iFu-?c��l��Q�(� ��-J�@����x�$�%D�}�Z�]��S�v&�S���*g��G�i��]�X��o�&��pG�!�o�XZ@���gX��a@�O�}NI2�%!*�}�#�2~�;M~�n�#�rE�F�d��;�맷���Y:�/\_��g`G{�v�QD�~��!���,��N�����k�QdkLx��dĠ�� �W �愕d_��Ʈl����M��hn���bv2���pJ@�i��<	0�Z��Z��~����e��L���f��|JnTC����;}�J!� �v�6�S����_���n��&h�B��߈��c��DVA��IGl9��o�)q8��M��p8�*��Fzm�9��ᤢ̖2����,�՜�qu+r�.TԐ$�T~a�����8�?�z5�͛�K�s91�jK(
h�m&�-Jk�C��h>ۈ���o��ĩe���i�@SGTT�f*%��L,���Ŵ���@L�h�hU�}�P;L<�-�kç�u�.О����?[�N��!��T�|A)@u�S�r��X�zT��5ӏ��(OiY��'.��o���8��a	�l����E�HZ2�� %ԩv������c5�����؞��s��8/�:�͍d�C�%i|�G�Hd����ȥi���=޿�0<Ku�F�)��8YWs	$h�7h6�иSP�ɑ�*׭�Q�-l[����[�+|��ajS�JF��Z�+��
�w�J�h��a���b|Fo���t�M�3���($~N�B|�h�E;"����H��oxT�s�_�}�)��AK|p��i�`���ۖM��:J:-�:0q��� ���L�)y�ڞ��Nf>�\�����"��.b=�\d/{��W��P0�~+-H#z��ƅ0�qN�k��5�b��c��S�ӷI�?�\�i�Z��h-Y�jR�߮�Ϫ3ӽ�d`z����K`_�~���%W�R���"�Y#�4��di� #0ň��,6�Ѱ)o��q���@G?��{��;�b*D��=��!����@�8�-ܶ�	eI�)��k�!�q�˕���an?1�M��S0�B��#��U����3[q�ȯ2�����l�/�t����}zr �THǀQ�$tr�l�^j��k���x[�K~�+��#��|E��y}�[v��cFp��t���̑M�S�n:ҋڟr'l
��>F���D��P��e$���-N(leS<m�Ȁ���ũ#a���.B-��G�%RX�Bb��!��n񯊲�/��`pl~�J�\�C��T��V���ݣws���¿ ����Q�5���c��F���X�v�bb[i�	F��%G|M}���a4i�+$�؂�HC���6�ȍ�f���)vF�GB���̲E��eƢˇ�q���B�C�bd6�,99�9SS�aJ"w��{��d�ytT}��|�HϨٻ���d)���w#`�b�����Q����x ��R3 ��C(�4+�����ﲌs�~Gt6Q!�j'���bNH����`A����w8t��}��ҿ}@/�~E��a�~�u`��J����	���
jD,�I.'O�7��B�Kq@�s�9�����҇P����	��IJ��F�5���¹t������J;���B��)�\�r;��/8y~s��H��M�:���r�A�.
�k�4z�3ƔT%`�ij<pͯ_h��P���$�ކ�.�q�A���ϰ�s�=c7�I��s`�:���|��kN>�ǌ���v%�`�����c�(.>�����!�M����~��w��O� ~��,��7�F�����b�s�FrM�U#Lm�î{��xm_X춝�\߸���Ў]�����Oe![�/��g�&>9�h�z��)��L�T˻��qK�~�g�U���b���!�>��X������')�^�+JbfNS��F�AN}�jۏ؊a���=�0tz�p�a1j��B�c'�Z��GU������T�(c�Ϯ�_!��3�1���DC7,�����[�]�gm"#{:�p@D����6�ޖ��ڒD3]UvCLWȄ��  g(�[�;(�e���mq�P��x'��S�(���HlC9���a]����鄦�F����L���+7�-�ۼ�؈Dj�a6� ��b��"������\�Bĵ%�yԳۭ�^i���`TTL�#pe*O֓ѥ����BQ)���^�,L#�J�����	(�>�� w�A�U��U�/QSD���9y�Z ���\�M���wg��c<	(��T�(E��:� �#���)� U��k��(�v۝����Q�ڡz>Q�{�B��c:Cծ��A�"^7�B�c��(~���y;)����3��� �t~��$ʑCZ�3I���.�u�M�%u:d44�+�	��BO.]�CUP%��Y���_���1�;�A7��	���Ѧ�}����9�@���VF�}�mEB=�.�$b�mS���~+f�����_(�7B�o����~aBxn�/���-B��k��d��Xe��;����1� �?��S�L��@��u~0�f�1�O�Mn0�����
[���f��3"#�|w��������)R�o��SZ\y&�R^��A�\��smϬ4#fC��]h�x���30~a�;YPq0u/�8��g�$X�(�3�_������)u) צ��5�4��ݝh+���LDt�"{����3����R��	]�b'�{��hq��{� �;�I�YH��ǣ�װʆc>�C�2��sWj8PjK���-�z�!�r�x����H{�� ���1 =���P��ʾ�.u΃ �c�m�w�*�Di���A�A�R�_-���H�+9k�e�	����ֵ�2�=��;ia�r��w�O�$`���bC�0� :�5d�qt�)����t��%��!�;�ә{S��c�/��e!۫>�3�U���sw]a~>`��!����[1���q�nw�7=bD�eW������,�&�[��&v��^��7��"�f"�X��r�b�x =F7`�Y(�������+�V���B(ͨ<��oE�,�������B�Ֆ1��Aʷ�} dMЯ�h�P/O+$�fl����#�A�]cv���&,���=�%��oUo�@������ɝ���ķ���닫&lۛ����5\����1��CM��C�6WQ\�buJk����漚��h ;S���3W;>����)�����%V�s�40��%�1,K����D��[�oc��r
*z��% ԶU���E�i�ۼ��;�szlA7���_	IxD�_��Jsyt �����ŮMqTAjV����]<�h��y�|�W����W gI�8)�Nr([�Cx�?��[������F����̦9�&e�(\� {M���hf���$2:�.�JF7 ���Q��66�c1�X���G�i�@�� /v�>G� 6`z��������Y�|�7܇�{�}��B��8#ؔf��x���wɨ;��G�9����|�i���*�Q��H��]ř���Maag�S��� �S�t���9�u��}�$:4��q�^�_���d�S" I����6��uԻ���Us�v�gNa�r9��T"��>u�p`�!�5���`�����-nʆ��ze/$O���~��L6�h�ѩ 'H(����3��8�`8��
��WO��Gٳǩ���\���Y�,y�ީ[p���=�_V+8T2�9��<m���,}�,;��'G�x?��&�dA���?���!AuU��2�0*��+%<�~p~T7hb"\'N�I�kqP�G	��0�����Y�e��u.j�������
M�-�yg٢-H ���
�	,��L-t.S�4�}��g�;���>� կ�>℔���\�e�6���ո�tWD�pA5W�]��! �{U������Hj�� :��%�������B@T��+l��.�����|1�骵�c@#TZ��ڇ_`o Y�:���»���oY��J{��exQ#@��Bny�O:��-L����{�	L�i� �*[��	��S�9f|㜽�{��QT|3�V&ՠc���������$�z�a �|DN�n֊���|�P�����Ĥ!�)���a�oS�W �ǅ�aH�S��������1C�}�<�)m��%�z6鼋mi'�y�i>�w�Ck�u ;w�m��ȏv[�q��˗���h���ή� �3Ȍ������cN�l����o��9%^��ȍ�}���$���;�Z���M��rÐV�5�[
["�������X��lJ%�9u`,�ly���TʄW�Xw]D1Rߞ�HOjjj:E�Tq�����$�a�>��O���m�eȋt�n_���"��i�;�{�/���0����DT�a��kAs��dU�.�G�Z�P�*�6o���~��|k/g�|�g�����;�w�#3x��P;��L����vK��~�,-³qT;�=h�&�(m��Jm�)Ʋ����l�NةB�xt�4i�����L,.�N�V�4�	�I�n����쌹��aNx	�1;n��M1s��F�/��uf<�=@5z@EB�A_b�<�2�gU3k���ǲ�����	�I�� x��m;�CC�I������`�=?R☂-	aDX��]�1�}�YBn�~�m�!��h� �l�ձ~ZC`Z�:�hir#͉���Se��!R�DE���Ս������4�ۈ�[ ��/b\�NO�߆���� �[Q�W����~�r��x(©��IC�V�`�fs,pG�l{�1Ra4��4���Ax�Bcx3/& ���J9Nt8�dO^�� ܏�FPl��ʩ��d�+u!�m{g�������k�Ⅼ[��m�*��\P�V�J���*^3ș��_6�|�E�<?�9��L�2�?��5�Q*:�g	��͜��_�q%��1�s
��i�)�����P[�X��f�*g���  �E�B��
u�jjx�	�Dtf�zs�m�H�ZL�`���,�'��)J S�q����ۈj��Ti��M��H��^ЊO(�>�w<ꄋ/�S�"��pW�so�7�U5i�a7����N�5�,�&�g�Q���~��_h�U2���;<��8�s�wQ�w+b:H�ef�F�\TC�QX��\~��`̶�����A}��Ŵ�.�p:ǅReJ�UT�t�j _�O�l��j~F��c~n%��>B��`���+�RX�=��Y�zf�qI+�A��]xQ�3�xr��2�W���j9���Z\������Wv���/k�$���`}&rT>��+mO���M�-u��t��<���?��Q�O��_v睯=n����%|ǈÜU��W��.b)���y`��\������D�\c!7~�yXY��A]*��^=�9K�2��f ����G�͋!���"D6��
�d. /;��>W��.��_{0�P]����u�`%��jvJ-��U��}��<q!���r"Wq��3�*m��em�ë�w�7�l��1��#�Ey?/Гד*u��b1�/Ч`)�C���=�	ῧ��b��Tdl�<̥ &ùnz���.o�����[�1��u+���$��m+),ȉ�1[�9i]i���y�/y���%Rf����8�e�gn�u��G��`�d�"�~�AF�x�L᭞8v,T���s�\��rE����n%2��3D^3��$g^����������N������
�Ky�&G��Ip'�Pxd�7D�t+����x<�[����Ic1�*\𝵋[�況@�?�N���7��t�  �kU�C|���\le��g��4݋_}?c2ZVl�0�C:�ƑN���bCs�4��9�w��I�����ƚ969�D#����"���E?�H;�#/��6��F��9�֢fW[�Сܳ:����1�WeJ8{H�ao�2�ťt�4p{� �9\4E�٥�ԋ���z�P_�(�J5q�2�L	�O��.��n:����5�`�'+���'DG=��V��9g�P5]��D&�@N˘h\Z%�b9�k�}f5U�ݏ��i�����3S0_�G<ͮ���/�kQ�U��|�
w����W�JQ�y��8����j*��r�)F�9{%F�d�m}��GqV�1	�rG�O�S�J�..a'����}�v���L���h�裎B��4.�2
��\-%bmB/ו��Xt����b�n��>���w�~���)��}q�,�Ԍ`U�Nq�E��d1�%�6%@��\���\y�IGb��P�܌����0nZlM��m3�Q��D��Ç�ъ�8f�a�?+�Y��`�*��R�}����fFc����zT��$v�Ñ��&�T;{���ő��QoO��6��H�ލq/gg�5
bS��<c�+���j���Gth-`eęwbװ^ؿV�%	9���?���?�/��M�6�k�r���/O����q�	�j�(�v<��a�Z��QfQW���\'Ɲ������>|v�N�"ISd�5D�|"����*��@:�%l7����@^����|�H�^{����nC�4��JD�ѵ��٪����;)�b�Ԟ�g+}AW�1�{�m�b��nO��L�=A�9�h�,4u�oַ�����_����]Rx����jc����������H��[��6�{3\�����E�S�����~� �f�<09@y�~�ō⠠oD���5�Q���Jp[��2�@ᝐ�N,����tQF�DB�d!����*��K>��a� �~�>�,�����Qݶ��`O�8#Z),�z�t��b��P�X{��(�OJ�g{�&�;E=�z�"4�� ��{(b�����k��f<�ipʋ�@�W{���µ?L��{�Rѕ鸾უ�ǵ��r���KҤ�|st/�qn���X�ez�zaBK_�כ|�C�D��'��7j`�q�ꭃEu[ɖp��}3��,V�j�^��2�(�v�8OX�="W��_3J;J:ϳ;���Թ�Eޜ�J4(u9��a_�9]�C�y��a��,�Ί������/�A�g�c���4l�^ ֏~i�O��!�!��2J�N�r��C2������)2�X`�Ɩ��u\jWk$��ۼ���1�/5�$A���?x���B�&w0z��E�pK�9��}�I��n�����	!D�xe����93,_��!U�-��2ᄇǰPx� ���~���88H���;T¨�&,y��IvɐbY���?�-�l�)E��;_�]I��.�����j�� SeJg�$� �N���ێ�[@2�+4��ƨ~�d3���R�:��ZBT ��;��7#�q�l�s�L��JB��έ��ӑT˚�����Hȥ�Q�^�!�C���V���.ҁ
��>��Dv���ڔ��~
K���R��7>����|���;������;�$�S��9�c5�w�h��yl����`����#�x[�	2��rU��-7]�%���
::�.��'U���B�f�ɇ���Ro�M3a����r�r�(�ݞ�~�5�m���/#����Ub��cB�ǻ�u&k�!_\�z��w9x�@��V�d��&)R�
���^ R�%��Ov��B��H&��v؈�������?^�������^(8i��#Y~�8Eq���<�!��m�T{ʑ&:O`^��M�gqܗa����ʅJe�kn����޷G��fȔ�	�@t�\lGy�w�C� ��U��./\�)�'G?PQ��'���Y��Dތx�Ͽi�%n�?�gȶ�|\2�D��>3�왠�܆K�kK-/��hńȆ��ņ��nG��D��@��1��f�e}�2f���/#R�=[��i3ŭj�9��,>Gp��ݢ�I?ֿhY@� K4�)o͝�!-^+����Wȿ��5�߳|:j��<*�p����E0ǰ�Y,'챚Yi���0�*x�u`rVLlٟ�re��ژ5��������}�R04~��ҷ�;�<Aՠ�gd��
�x��h4x�Dv�dn��i*	J���|D�oW|�ps�C�����9�:J4���Z���b�e�p�w��f
��(Q5�8�S���'yޡǭ�Η�����q$�=�'��'uw���!-�b�ـp�J�����Gf�J�������@�;Z=ě��H s�l�=�}4I"(js�,���UJ�!�9�$Uw�1�4G�1#��c�'�N�C��I�7P�1E̓��X�=��ϛSёG�>�eh����kl;���r� ��}�	7qm�G�ޙoa����D+���u~j7�p�6�?�l;�����NN�)�W��ј$z��/+��Poo�e��眊�b(	ѱ\4ؑx��g᳞
�UՀ��:,
��`)�#�ؘ�i�&��(��ݾ��Q��/\����u��V��d�P�v~F�(�m�Q�ׁ���׹�h^:�*�W����O;B��Г\�2��&�"�J����3Gy6���C��_,�ʙ	4Zlb<�tG�R�*��1�>N��zC��@�O�F�>�~�ɄL�{^���o��/��	J51���k?�
K19�tm[Y̦S��I!Q�E��5�H-6�o"S`�]
���ϱ���i�M�lb�r���%7fY�����I���G�	�~e'BE��f���W���@�βDjqs(�Ey@&.{����X����>�)E�y��.�՝��h?s�*!*L�hY�68��ͩ�SNkZ
�Юx����:�bg0������}sL��)���'�h��:O�M����x�_@4�Ⱥ6H��r�Y�G�^ݣfg7~�O�uM��]��!��$���Y&x����^�:Fz���)�]4;�F$ʉ�e(�%�ܨ��d��ln
OP[�c[v�������u5��.�uj��K�a��	������`D��Ĺr���'a>p^��B��VH��;���m��Ã���6vg5�n�K�t*���؜���VF��>X�gO��+���
�bUӁ�(�]5���ή��t+����.��=DvI���68g�yl�Z��&� �/3+|?9r���������!�=�(�f��8Cs�%���XaV��P�cD[�کt�����Т���k��I� 3�ʻ)l��Aa[�������-�';����Y��/�(��γ���6��w���%I%;�]uY��=���6��T�f��L���+Ѱơ����c�����2m�7���Z��њ#@f�9m������$��[;�r �5@x�i��{%�͕����nubo3���6�����A������_{L,�2�o+Zf%VG*�B�r��3k! �ja�0s�V8� �y�5�����E�
/�}�:�O�Pw��/5�S@��Ql���i�r�m9��:d	֥GM���7�@ � a���Da�]�fn�����?18o�Qb��G���D�pS�y��w��YB5�jř+D.�Q�(�	[GK(;���"�}Gާ]�9��;���E1���6'
(�pT��,�s(]ó	��2.�ӳ=�w)�+�,�)P{��?�B�0��g��m�'8v~�K6�r����uO����^��L�􅕮�UH����MR��r��7K���TT�\��X��[��&E���f�Ǜ19	у�.U*
����1��<@~���'���%�T$_��׽�+��aRS������������iN��[���H8@̔�XV�Y_� �!
(�m�e��Y��ڕm�˄_C��=̩������|���\ia�v�2��̳x����b�e��?��Q�� hv�m�e2R˔sR�y�S:4CT�Ș�lԡgN�s��ZP>_���e��|�+�tGȇ�����h�'A�!�f�%؁��*��WMn�I?�����3C�����|����.�ǧ�����z>��`\LC �6^�'��h?��yM�W�A��k�9���~9��uz4���L�E0��`�@�W`���P�&��ƹ��h������$,�8�ܦ�<;IUi�����{ �*���K8[2�C�x��y3��s�Y@y����T�g��ʱX��1�f��@�����G���E
�	*�(s��Z��u8�p�6�!��̪P������c�BDB��c�?�y5r*�^Uw�S��ׄ�w
�a3���Kdi�d&B(�Y/!v�_�	Zh^�o�Y�l��� ����gud��
�G+#�יn��cs��Q�S!�@����ٛc/�76vV���+�I��@($)dR��9�{#�K�'���i�Iu��g�}5�z�:�q�1Yv�=�(\�"��]��^qd����&a�z�M�냺�Y�Um��6B0�jÀ�
r �����w����8�"��kLj��ʙ�'?l��i�*�l4��-����u�{,��������v�>�P��^]?�)�� 8��ȬO�9�)��ִ
$J?�`7��\e���j��G��X�6u��?�?߀t�����p�6�lcȍ�W�;���D
�T��N�c�G����a_��a��
X�iףH�؜$�d�<�A����4I1�dVQ�KI;Ӝ+��lT�����۟N�UΤ1���OP���'�b�� M Z��f�Q�x3C�43e���v���;2(yW7U�E8��q����l2g����"Ar?����(�%�Mݾ�-|΍�%���.�X�C�?JG��_f}�u3k�AF�y'���i*�(�B8_�Ī6�NJ��E7<R�ߔ����Ҽ*Nb�3�?�(�x姶-;{��L��j�Ne�Q3nP'4'��K�E�*�{sW/��q=�����i��#��9 ���C�}����֥��ޓ������Pw�Ռ�����O'�#�
�@~��qJ��(y�cc����;��o��5}��R��@�O&(���LWã���/D��
���fO������)P��m�"��ǥh���ͯ)9�F^S����ot�F	�+cio���S��;�s6�R����8�]`�<zn��ENU,Yx:�\�J��B�m�%�N�m��9�ZqnN��I��]?^���P2�=���EA��Z���Y=��{>��b�4��>��!�C����z�ii�i���7D�up}0�!}I���;-+��]
/]���>Iޅ�%*�둛uM�2u~&�Bn���U
���<0O�Q߈���?�,z0*�	F4��n�dhU�ͯ��~�$��P��ha�ϱ�f(��1��^iaWPT*׼������[��B8Ҟ�'�L��3�|F+���~�����"'U���d��5w��3����\[/f��C8N��
��Ӄ�����M���ʹ&�X�mk�m��bH��c֮<�6FČ�?� W�_��P�_�7?C�GF�38�./^�ƾ�N���z���sBD�䖴�Td`��g�G�C�5'�t�L����t�W�?ڈQ���^�6u0�1J�tSx�x¨6�]]YW�������/%�N-��?=ogc-JHx�bRS2��BTO�8+���%Վ68c�#���+���U�Ѝ�$��L�Q:��U�:�<�x��F~�K�=`m��70̽�$=��_<�>��^���!@�t/%T\q�-F$�z���O ��GT�#3����Ϟ��G����#���	 ^�=�輨Զ�����َ�i����7`���a����U>���Q���n�x�������0{f�A�ۓX��VZ����$�e�+�]X����8������Z>�f�¨U��J��H��Z#��E$Yd��<)��Y���|b�PMw��k:��NQ1��%&w.�@��}�1M��=u��U����W8j�wkS����\O~V�qo�	o����P,t��<w�A�5��,d�V:V��b54���_Ꮧٰ��d�d0�9U���Oh��C�X���#���OV܄��to�XJ�x��#����O�=$jQ�-��NB,��PD�Ԟ����D2�����.�fa�w��bQE#]��1�~v�{jpd�!h֜&ĥì"� :<�mC:��O������|%�c���;&l$I�S5E?R���5�۶�5��H�r�E���Yx�J�^�VV�X=?10�L��5�~���V�f����l����V�Lk��Kl	 ���R�FL����gx��Ć�R���s�=#���?�r�kFQ �2���0��Өz|�s���FIR�X��G������(���M�p2Ď�v�a\n�9�51�%Ҧ~WL����b6��=V��ť�e���Ɩ�2j���I[S���
��R�e������~Kf�m2�p�[����Јd�������u��m ����$�s��N���ms���S,l���4>(kb�S-\b�֠"L�pP��x���r�~��<-~��c����-Hߓ?_{ȷ��;�����9�����J�Uæ;��E5���'�e���v��Zy>��`�@�.�,a���xd.���e�|k�^~���k9訯�V$�m�P���UHzt#ī���e4�:w�Jg�����u[����}�Y/�g����$�nMwv����(�
�9����U��۽2G�R]Ce�[�����r��wS�%��)i�3�#�1-:g�#�&��%��g<ȭ�� H�y�4����3]W��&��M�j��:���Q���-ʟ�.�R�z[�H9nK���x�(���]/s�ٞ��a�|�$b
=�=�9��7K �C0!��G���6�
�H�y�<�z�<x�Q��Q�ۀx�"�Z�	��KWK_\~K��2�[�=>���7E:e�����AÊ��iGk�4f�vp����]pFFi	�:�k'��?�ި �<[��xgj����m8�ݵ^�w�Y���t�P�4��.�=���)g�rwt*ȕݶot�&�|�Eڝ@��(��������r�·��_H�/��zG�*E�����Ts��%�Zd��e�~�+G<��)Τu-��d��>!���AO�?S�:Ia2a��/����`�!9� ��o�,9��7K>R�=Y$'�-�@!!=�ˇ�o����~m���_���7���dɞN��<�++��;|�{Cc_>��/.y�޹��XERd��$疯���& ��{�?�E<W�c���T���5��<β�q�a%�\"̝�C��0[�����Y�:��wv|��� �on����ze�j�Z�^&�M>)�v���o<�ib��^��n���L'�e��mP��[�"$:N̵�i[�zH�rgd��5C@n�uq�*5�h�3@��No�F}Dy��%_{����F,��I���Z��si�����r�ݨ��EN��I��v6*� �����r��v��㷺�����\��s#nO��]��d�σ</�A��@�`�����bz����}3�䣾f��C�?y��=��aj���5�=r#�CB��*#���Z��#/Q�Lib�!-~4�W'��I���]!�����XOV{�M��-5�W��C� .2L��h�Hd\�������Z߈��CK�B�)�8�+��?F��(X�H�Y��:V�/Z�Ցn�"��AUF����f�[5�:+`�1J;luZ-� �ꕯI�Vm�o@��C!�ԙ��g��' і�u��m���jY'0���!�ll��B�j
��-O��]��{��M�D�p��g5�:e��ΛTI�&c�Ħ���'E�l��ќƍ:�%ȑp��Ʌ"�`�e���^!e�'3{7�rڗs����q�ZMe �����¾I���p�x-]|��Q���õp�-��.����x��)���.�M�<��j�hiT��t�X�n�W�%fW��������˳F�9��Ӄ9��3�f*�$�Dw�c@�ޖ�nݟ���k~U)�:fb��Ѩ�<t�C\rƮ�P<�H�_+QYzi&���0���� b`�&\S�ft7���PԘ�q7� �X΁q�n@�kT���8�"�3=(��/8EA�>���l���W���֭ܮz�Y{�g����_��M��m׬��=N��,/}	��6�t���1��U�%��g��JzS�5`���< <B|��.���������}}g��u�I�1�j?��	<�,��l��K���i��vF��Y
.�����U�|'�i��1[Ww���te�1\N�m��,)C2/�jJL� 4��%��� C��M�ޭ���}Ny�M̈́Rg� ��l�I{{5D���p�LuLr�b��緿"�B_I�����	V�5(���s���B�
�o�,�|p��5W�����t4�coe�� .ڑ��iK>�9��n0,�\�m5=������6W��/��I�z��͵E�@� �\�KH<WK�ɶ�O�>�aw Z�p���q�"m���\�Ss����B7�r��	��s�b^�-��46&Kа������U(G_����|�N\u�j�_.v9��g�����z���h�SJ�R���;%�z��Ғ�Ư�
j��қ Ns&�J�ӣ��F�i���o���E���$�d�����#&�	��Ǖ�H���_� ���+Z4�?�꛲��#�,z-]�C�(�1��6F�E�\��⠺�,�{h�v�6���y1���Yeg��ϩp�?����@�_3F"����|~!�烢�xI@9��,y�P:B�EqÞ#>��)�8~�O���:XR0^�I�o;�2Ћ�Щ`6��z�*�������z3��yUSa5�c!v���M��5�sOT;�D���)���;�u��Ⲵ�<��u�R���4�|X���Rc��/�qf�����|��@�k�@I�u�r�ٴ��!������w%x���"zL}b�g-�5-��2i as�V\7�|J�(|��ڰ��Q^��B��w���㦜��Bm�
H���ˈ��{��z�E6Y�JD�%E�����H*6� �ETs��l��A�z5H�&���(H0I�=-�L$����^>��W3DnC�����
LN�Ԝ��]��G�'���ˏ���Q���ݰ�wa�!LcٷY��˱م>abÉ�]]&7�""�E&Z�1d�2��F�-5���[S�g5,�X�U}}5��6��Ӽ-T�̈ 9_�r�x_/"*�-���SO�i��y-h4w�ł�RX] �x�YJ����eYG��7���د�z�o�_���&~g�*��9����{B�
���ty�Ci@���/mBq^��&�ޥ���]0�p訜���~gkp��47$#�w�	�*�.7Q��Y���M� 	�м���9^�
�Q5.�5j�^w>���8*$.�O�-O�L<Z�ƚ�J��d��r=���Ӕ��E�z`�\rkn6��3y�e���[�#ON���E���3c�4���(���:?v��q�	U�܍ �0D���֥���saE2�qQ|�
��	��y�*����%���*K�>���L����bl��j
�&�2?K�#�	�4�eSUCi��V����~~��W�ܓ��P�^���xi�nH�|�K����� m�/��_�o�=t�Yl���n��V�T�Db����
�C�3N�K~J�����i�!'�r(~��z�g��|W�����hA��1��z���1D���7]���$����&�e8tN�$�����Cz�o�s��-��'-���)ڲ��v��B�x�+��bo�b�6[OX�j�|�Y��K������Z,g��Ȥ��W���ODEn�M]v���
�L(��Z�|���Z������ޑ����p��eJ�TD
��N_��"(���<�4��k i��I��1w�?w��ږ�qM����|^=�^{?%V�g_'g�l�k�yF%��j��OU
�_ �J���gF�gV�m锠�Y��t����l��(���?o���M��m��@�qRn�������]t��μ�6���\}Jho�R�|�p����W~<4���$�M&۲�����v����
��t�5�����)��=���c�_�s_��oG�%b2����5Z�QWx��֎��^_ �dk�Jׂ�%0��S��Qex��j5�Y�HBB�퍌��[SJJh�6��|�r���I�;���G	�H��QFH��}�Z&+%�-�xPV�u�((�^p��7���Z�Pǚ4�|b�q��y�PS�;���Aq���։��j�=7w��j�JuOH�5��H�������F��^	�%;��>�`,1L�S�0{97}�(��]L���p`�}Ub?L՘��>W�?!N�a�R?P%��rS5vS����Ϲd�~�*%8�\ٽ"A�,N�3��J�B,�܆�5uC�KƲ� ���1��.3��*�2�y������i#�ܙ���H;F��y�R��!^�3�C��Kk�w��@���UZ�Ez�����ҟ~�*�LG�T 0
e������m�[����R�V$�#��(Q6E���T%�f��H�T��>��p"����(;�)�����^���:R�?:F���F���v���d�L؞#��ł�QV�"���uR�{��`�2��Y��)F���m4<���@�T��� `�e`z�Hd���'�ff�"jMݎ&��i�Ɩ/���F�)�k��"��#��v4(t�����~'������x/������J�����w̏��;4q���vH�N.Q��܎��O"{�$1|��ɚ�#^��$�1�Bғ�ט���yu�),*�����o�3�������;����6���jvPT]�i�8F7j^�*�l
�����f�6z(���i�ܫ�!���wʸ���o])2Y����P�KZ��������/B�ONi�|� �ܠ*������<�L�q)���w	`��V
����7{��"1��^���	�Bw��U�ǈш����
��N.Ĥ>�"�d�T^fN���-c�U7-Q,H:W�b���\α)���~鉶92����|��U}3AԱ-�j�	����j�_iC�}d�D�;z�о;ഞ��7�	���nɧ�T�Bu^���Tua5�g6H�+>!ȁ�Py>���� �4fhJ�S� @�������:������.�w��1��w� ��M4�ݒA���ТD����@����*Yv>ix�L���7f�{}�-V"���H
�|~�g��*B9as4q�qva�"��5(`�Q%��^z�C��(�����o�JaMb�M�}�)J������+����7��u3���cZ'QXoDʹ[E����@��_e��?;)�^���������aQ6p }w�/@*v���OI\�#iƘ,�H��(�j��%�C��sE������p�R_Q�Kǖ3�P�y��깚�N�G�Z���Rn=w����4��m���":a�Ҥ���U�����C�M뷏��f���u��A�Z甴�����'��T��%%i��tӦ��!�ĵ<@�W�d���*�+d�F_U��ûm�	M���'� ��0���ie�Ds�?+t>�i�2U��9L����}#�g).�`�νU*b�OM�4O� <�Y��F`<���o�O��s�b��VF������׏#V�n���t�"D����Hu'�����2:���}�w�0C6�����d�!��ϖ�~w��q���֝OB�%?��L3/������of�I�m������!P�H�y�Jhz��C���m���س*?wz1?����|]�a'�u�7�M
��N�8+�>./�HN_FB���0��B����q��_��u��|�Z�m�[r���c�29��2Κ�Wp�)=����O8�7�����wNwK���7��$P&=���k;t�/N*V�M��򣻌C!j. �Lv�h>�iY�?3�)���z�H������c�(.�Ǒ���R�?��ee���0�Y9O��w��N��ʡ�1�T�M��O��J�0����x��̀�0Y�s.��9.jp��/����z\�)�	 ��s jЂ�K<\A|�\u�q,Ǫ��<ju�<�7zѼf�d�s0�c�α���ꨧ?��ʣi�?�;[�dê��V�*�,0z&V �w��>��}؃�&�����-O��x��(��+�6*)H#O@ڥxX��Z��WB�.p~���K*��ǭ���/�X���|��KI���;<��Щ�ߔ�T�7��:={Q�3C3g���3���砒��F��\x�F�ձ�����s�f+�cdv�S=ZL��I4���P��� b'RB�LU�rFw�p̓f�F�&R�U�͸�E2�Il�0y1p�N1N;�}u΢��Dn-�0<���=2C^iE��BF͍��P�<!\�b(��Q*m���	�
��f���DnD"��X����..�{� \�ٚ�B�T*��1����ۺ�Q��["th��W��*�T�(�/tb,�&ydH��O���s�@rC������m7Y�M�n-��d�6q��2�*�?A;�sW 9����?�#��~���ͩ�˂��+�����߯�Q��h<'�d�:}>,ܦ�r���2Sz�|�2��B1l�I
���4���e������8�߉��ÿ���A��VT����>��i�SEq~99�4$o�ϓYвl�4��K�Y9��% ^6n�$	��H�[�+%�J��m5(�<D�P��?-m��Z��zo�fa�h#)�!�ْ�!�pqp`2��g���U�j��T�յ
�E̈R�j��e3m��j菓��&�H�MA���A0�Jx��պ��~�=6�s���ށ����Y4�臼³��?p�/��r5F�lbI^ u)jc�9�驭&�#�:��s �q'��i�躎��4�3s�g�{0;�GV��f�ؙ
к�6�#���Ղ	��bG�n�j�
���QXꚾl�8W-T@"���u��7<�!�D�|��YI!(OM0�{�;�,��/�1����;��ԏe�*��e�]��=��!���'˩2L��9Gh�2���V�ǡYf��e������л��G>�*H��f��%m5Nd������^�ȴbt��פ�%4�2�|���~��� ���+J�'�qVn���a������|�)��bϋR�	����9�����
����ɕ�#�)�8��{UWtF�,�U��M_m	����!:�������7�޶�/�V�h�
�^A:x� �Xx�iom8Ƒ��5�f��v�}�7x��k��(�h�R����aAj娸���,��}�-ӷ�K�LQ��R�y�+���~޶<�v�˕�#{�&\��2=�A��A��������Ew�y����Ir)B�[$bI�����l���ڒ�=�m�Um
��_����U�i5l3c�_�ܝ;�Z!�ܣ3��o��ɿv�'n�:���}(�cv�p�SF�A3���c����S��<j+�oI�V=�3P\]�&�w�&�o|U,�&�Am:�S鋏�	*Pe��N�ؤz �x!A��毨d��{�]I;�+�MO�����,�!m�!Uu�g��7���{/FY3zR <���~1�xEɊ�bR�O���k���"�	�H����qjO�\����|�g� ��A��s��t"��)a�p+��
\R�ѳ�Ţ�WE�&z	Qp�ߏL�cH�q�F���jr�����q:��k�r:�-k���,���5l�\�C���"#Dde�\�PjRᰘJ8�"���z{[��|���������.%�.�J��/��u�ǌ��!�z�@J��O��qȿd��4z:-� �[�:�A�v�:s#���\5t�!K�bt}o)
-sc��=����zMEBj��\��R�ɤ�͠���l�2�j&���K>��C=�g��;�fBϼ��?�(���DS{wt��BƱ���CkY�~�o'��|�iC����!��7���Y�����4�ԑ\H�{RC:�	�|.���*���5�����'����֬�������<H��vj��- ��riiE�\��,'6�'`�s�̶��w��$t�#�� t�
T��M��גa��Z���s�}�`�I:�:�簖S�I8�z����0�>�dL��d��D��_A��[ ��VP���_ͲY"���f�u�VD��݂�a�iF�z�Э�#%�׆�eY`8��c&;�I�KӶX#��Xe�}�o�*��S��wqY�N.	�ͤ~ާ¦M�	�g��2�(�W��9�����*�+Ն瑰�9�a��K�N�� Մ��e�%L����O����j<E�n6����T|��5ă��<PU����>����\��yH7$?��R�٦lZ��N��[�sI�SX�N�:p5!�N*�|of��U�����Rs�<p�{̴U�)Y��7Xݺ4ik�c\(W���s���]�6U7�Ȇ)a�Ĥ"vߋ�ų!�U� I4�e�nE@F�j��»⫄������e\��"��56k~抍	X����-�"i���W&�f���a1�r���x��&�>xp>���5��GN2LwB��s��?�����?(�+�lܿU\���m<�)w�cP��:����d����
yY������L��OBC1,N�A5(W{Y}%nʧH<H�$���^2"}���.�Wn�) �&������C���5�t�Q;/�y#T���d
s[8) G��>)�% '��#7����^i6X�;�_u1�k�w�{+��3K��D��+���G�����G�)vpa��ƕ���S����NE��l�ܼ7x:�+��f�(j�¢���B�UΆ��0;Z�	)#ZWq���r���ʠ���i����g�.B؎���;I��:���f���?°'�d0�:x׌��K�i&s�J�`a��2��9q����}"3�w"��0}�����v���SAD�3X�X��d������y p�R汞���xT�5�e9p���l��ử���E���������X���d��*L���AP�YX���C#Vł�ҋΚz���w���0~��N:�p7�ytt�}M��M�?	jb�
��kh9�)�NH��I/��t�ɬӑ��3~�ԝgNw!%;�$7q	:���-Q25�`�]%�qp܊Bψ\�4� ���RCO9,����ϯ��ߪ|���:�]1�����g��ɢa(���I����㯦{� �^t����|���B�@m�}�R1!�I��x�}�~F� p{���D�������Jv�r���p����uvT߉��m���QC]:�w��!=�C���S�=P����j5l&csE���/�^���l�6Y#x�&��B(Y�Qkb���Pc�e��!���%k[O���q��A�}ݤ)�n�=\bi��p��*p��>5�8�.O��PZ~Y�4��F!�U��jV�8�?@�!�c�BX*ODŨP��2j�5h�!e��ðɊ��P�.E^��X�)��Q&�K���+Ĩ
����-$xj*��/�7��/���ǚ|�mN�QH�`ֻF�[�3��`Sm�.����T���-���E{�P J7�k����
��_ǖ�v����m*B�k�!5y:+P�G盚J��:��k"b��-�>�����1����m���גּ}�_"����^�[����#Q"w6�׈��1�8��ϰ&�[�]M�ɛ,e�U�V1&��c��w�p>�����^	�ǽ�r7qh��g5|�>�m��)�ǃ�\��GgY��6b�5Kk5]��CN2�3���H_�=ए�ͪ"r'��Ku���ʀp�Z�_�cwz���h	�
� }S�<
쟒G�~��^{��qmtR���T�z����"z�n7�7��Β֌��x�����i��W���Q`�a~���N#�PG�?����I�[-=�����DR(��OU��	Ho���huF0:"Q*2�D��7��� ���[�h8Ahi�|%|M�D�5�qD��`�6B�����$���i�E@N��[ۢ�Z):��e�˴�V?�����h�.�E�L�h<hQ��|V�x/�y��
pj��j�d���gK�����,�Ϫ��4Ws�9���D����4Ѝ�ho9���N��0�kk�c��*�U�9� �c�N3Ps/U}�fEocB���J"3f-��ٓ�R�i?�Ǽ��&�ph�hgk*߀ڝ��K���02�A�FW��@�}ퟖ�k"�Wˉ�AΝStF��Ob�ZrKF�7�<a�"`��Ed�f�!J�����9>�2�]�KS��:^�$4f�+K(XS���i�p�(��#o��u�(ŻX�a��Y�챖úAc#�5�kSZ���ea1d���*#υ�hg�YO�#��P��#`L�2b{8���Z瞧�i�M�4,��f���݊ڏSp�	dX��;lG0��|¸�v�&�]�F�I�9t+��Ҹc�:�]Pk���N˛�=���]�SaPP66�CL~5���Ͻ��)M����J[D
KrPVt=���^0.(�Qߐ�Rw�O��-�ۊ�)Z����h>�SM�iP�)��<k�!�ݹ���jk]W�Rv�f{/�����
��P�w,T�\V�?��������K�`c̐��Þgy��BɼL]���ţ�����fE���w�e�(�
��Gm�i�xT��^������x�T�F�|�}��M
4x�����yI%h븣�1��7)OH�Ԓ!i�,Eo�B��}���p�ʹ�/�9�Ĕ�ɇQ�;����؇"��xF��ܲ�E��TzR��u;�,Q-��L.Ha]�j{	|K�K�E\��˱�ȌO�oeb�ݤ^o�s��ge4{Z14�3,��� /� wM���e��N�e�u«��ٺ���i����䎎�ۛ,�*g�3��r�!M���mf��Qֹ�h�7m����ɲ��hG_ϓ����4��"��T��K-���0ӭ�����N�_�K΄B ��rĝq��]b�����.7��г���2J,��-�ʖ@R8p�R��W3.L��I+��v���w8q�ו#m�sh���x�s�M2E�U��Mw�z��	���1�x���'�DI���C�����e�=��=fH���l+Fo�Ȩ�"�`z�Gg}�|˺�N��$�:�S����Ùz���;�C��e�+�޽���>����2��3�ۯ�a����o�?A��&����!M�<���ז������qF��W٦�~eAE�<PcD3a�Y>�F��/|��#(ފ��{.6|B&,�������iK�����������3������D���BLG��1^� f���4l�T�u5]*^z�M�>��H#�

r%p��� ���2e����urD'������ˋ�_��[!lfI���Vh��?p{���3�a��#0�z�I� �����m���0Z/|rȊ��R	��b�0A��ސ妧͖�N&����T�t�gQ��R���e���zrdW����jY���v#����/��o�-q�qʪ;),�ᔇ�9���ͼtL��׌S+s�Е0�Ř���w�X~	����%Goozxƣ�����s��L��`��-���Y��n[����i[�B<u!��Zj�#!!�l������5�v�?q���`[]l9T���"ut<Sw5m����s���]�-�'��'�3'�Ы�+�AE��E���59G��λ,��s1@ ]=oa����k�b�p�g�<��E�S	�7��b�<���)������|���,�M����Y�z�������\G]�A��\�a��w ��YW�p��d}��>����>�� �ަ�@�)	0R��d�淀�ﳎ|a���m+�S����>�b ~8���͋ߓ.<�U�M��5>��VV�.Z�]a��qչlU7���!�MDO�
�9���|*����֊��	��!�����.�x9_Kon�(F�W ������>W悖qMmٲ�赠���KQ��t��SI�]�f��_ �<8�8H��Ϛ���5�[>N��%s�m�*�>��>=��n>~���=��[^��2Fu�`ņ�W�b�ך��.3��T�.K���ͨ�q�]�PP�	�p��%��(W�L;h�i��&�?�hK�
���1��BW/��0NQf<���o�l���ߠWLۘ����Ԥ�1���|�v7�N�8��[R�D3!۪���?Ɋ����VQW�qi;�=	�E��LT�*y.x�y�T����B�D:�\��W�>D��%�$�DUզ0ܭ�/	��7��6.�甌�{pV*DEo�R�����a�9vF-�F�/z%>����J� ��r����5P��w��c��MCw=:z4&!L'Fej�K�q(����5�x_�Cŧ���uQ)�/7�ࢅ�Dԩ��" ya���?�%#C"�Rbw�n���op�������LgYmn��R�Q#&>+��g���,��ؤ�"u.E![z�q���Y�-�鎼�����[B����Pg
�8Ӹ�%bVr�Qtx��o���BN�H�986,]��4B����w�5	{�wJ�?wLV2檐x��H�F��*ES�*�/ʝ@�'�d��6~1�T���S��!�䈣�lE����D��~sI�&3NH�E� �dD�}(.E���D�9�[6k%-ɱD%�w]�3�P?��}�h��}�%�9�3�v��2�8� ���o6��T�q����q�n��?���՟na�R0�����)��0�x��������'9�b�SI��S=�����V��'~ ���Z,�L��v�1�����W�Ԭ^�p���18�^�Q9%·l��1���֜�@ZE�q^�-��w���~�+�;����<RűM� �^PD.�A�A�J*��&\�w��
Hkb�[s���W�6Q( �i�7�*�V�oѻ7� �$��s�1��d�Z=�б�ɮ�3>N�Y�3O����k���!^��E��
&i�f�t��0I�]�F� �դ[frSI�HמK�7����
og�ݞe�f�g��e����0�q ���h7w�߹�)��"�n���8���ƅ�ˈ�mt7�n�y�F�\0�����gk���0�˄�+���ȶB��Ȋ�{y�]C0}~m��J�T���Pz��B��`ʡH�۴��aҨ��J�.������d?�^���}�V%X!)��O�L��=��cB*LR��E��l���y�4~R�	��j���6���|G[���&[��.�F�8o�>X7��f�`N��}D���3?����B�cKb�d\,&�9XaMk����� �;Z��� ��J�-O�j�aF0��R1�d�Z�����b?��Yw]T@7���h�9��G3�����vt�����$��<w"-�=��?2�7uT�����g`������i��Y��<�:�i�s0clSm?�\�_i�"�^ѯ�����2��O�yߡᶍ���H��e���n)�S��j�
1b_��as�� �����\�0�ݏxu�ǭ��F��@c��H����������柬�`�)�P�DMn���
�z�W2F���];��y�!�5��fًʠ�0�ۯP�I�š��t��!Hҿ5� �,)��OA]er�Zcl�0��Ʌf-��䫔B���S�7>D�~㻝����MUot�"7�:ï�X��5X6�Z�#/�)~Y�Ih�����c���9���<� �!�q�l�T����u����*O��� ��((�B��^��ki*���b�[�`o92q62�X&xzUOd&Yh ��b淓�<�I�9b���	��<[�3�d� wJ?_o�(����2�Z��Dw�I���JCvP[�F%�J�ӆQ\ڄǪXb1�\{y�p�FUp�<h��ֵ�S����F���j�������*�F���rқ+�]A~_`\'F�0*��  .�ҍ�6R�
�yC�bFt�n�����yAjR>��!�U͙���C �|���}���eX&
��x��5X摅e���b�XkY�VV���)�{�e���e>ޙ+w����Gr�y/��������$�ُ��|��%$fL|O��lչE���~[l��$YDu:u�^m|���6L��%a����`�]��@�o{o?:�����t���jH�$9���R9���ԡ7����u ����'�;�c􁋞�ݰ��֖�i���X11�:�����b�n�[7׾Od���3��E�)&Ww�J���0�|Z����\v�J��aܛ����p�Ϸ!�Y?y]��z���<���4�8�,Jn(��+%j[�&��8���
�^f9���r3�C�
�КC��wDz���`ϛ��I�*}�6㏗C��xD�����Zr�T�u�B@�O��"�"4K�<B��s9�K@��#q�`�6�V;<�T�FcRɄ���'�b�ţ]�Q�Ud��S�U�a�@-|�<�f9�N2�t�G2D�P<[��nN��~�Z�P�Ͼ(c�:��lY��l�a3��dX?�P�:�
>���Y��\�Fl�[�)3-��h崧���]�����c����Q�ʓU�\7��2gY�5�P���0���XTΩ��+�����5X6����0f���-���'ziB�Nλ�P�K�&� �����~��{����r��p1��D4��,5�Y�.�C��0��#��7*,Q���w�+����{`�p����OOk�s��F�<�������=B�m�m�)VAs^sY8�X�H"�^�Oq���b+c)��7z
�Ј���2��h�N>��&�gl�w
z��K����� H�o" pc�g��D��a�Զ ������S�� �}�	��6��F�_�	:�=�6 ��}��>�#bT
�`��2�H�XN�i�t��tغ�D�+��D4E�n�;���i�4��6Hwr*+��v���TM{۱#��kǤq��a{��iq֊�0EM��8����C����%�Kf���[%0_�'��'����g7!p�i��@C7IIf��6湚��}g��n:��V��^ŕKJʔH�`9���_��k�6�D�d���l�c���s��S��^�8NWK��ǂ��(zـ�ޢ+��(��߭_�x�~��?��ݼf�<�3q�{�<�K��}+�󙸕���m\1�� S�C<�v!"���E�b���|h�K���{��� ���X@��B���e����3vo��L#�A�V'D�ͩ~�3Q�=[v��Mu�;������+�ɳ����1�Zl
��cA�ﲷ�\&G`]0�6��b%x��/��4=?r<J�1>���l�����HZ�Ѳ::M�*3.������t��N�d$T|�վ�0Ƃ���S3��Z�|k���(<ߛ��B��L���M�d��$���m�pb�`Z{A�BG��"�vu��aO��ÖZ� <�uNǥ�QQ�
6@P存���P/��y��t]*>\$��wMnˏ!#��	�)G��;�ܪ�*Ĺ�>�%�t#D&�m�w����XG
�0�K��R�[p�
��rI�a/&6:<F%?be���t0�:���1Nu���9�^͒ڟ������F�E��I���,��S�eO������G��P���{O�G��H��,
�O"�d��9�	:`�N����֒��8�I�3�@�
��݇�������?��Iv�����v��(�5c���(����O��-�!(�A U:��+@������LE*Y�YF���gaXo�=�K�B�I�"!+n"#�޿ꑱ-5YʶUL$wUset����1�t�xVg�J��"(�</h�VZ��%�	t"x�xw��?o�}.-o&_�qӼI~j�C��X�����#� �����?��C�c���A�Ll+f�`\�����^X6�L��F-�V�#�:4[�'�:�K�.�6���Y�@>>3��j���6m>�﷏��xb�O='|�����q}&m�˹|�A廬��8K�eu��W��rV|� �0�0��d
A�bu
�Pj0�y	z�v:�5���M��!L�9~�Gt�Ŗͤ�?�*��-!R��G���igT�r9�b�"Is_S�V��
���v��;c�P��LO�:���ǉ�2�b�Y-&롼[��I�(�ݗa�ol���_yN�`���i���x*`#�S����S��xWS��˱������u��9{��q�S�s&�o�*��H��Ǡ[��,*$Lw�s<q�q����N@ �o���k�^��*\~ԛ�7
]�#��M9(I�F�·5�=7����[�:e��hQ�M;�0w��lZ�b#�G��Y�ej���fឌ��Ri�'�&��;B�m�	3� !�#V�I�7��y"��;���$t���6�;J���`��]q�"���9��
ئ���
�D#TE,����m���tT6U�r��I�.SS���ik�&.����ҿ"G<����f
,��+�����r��w8l���B�Wws \�|N^_)�؈F�<S?����'bB�2�h�E�mr�G���GH�+�!/�z4'�W/�7���o�,'i�K�>�d�x0�s{�C���f#��o��}�o��i�wVvW�D�C�8)�%F=7#c�H<�<�,J�3Y��Co!�|f;�94ŋm0\��2Q�i�H{A#s�<��c�ڒ~��\�d�s���RL)��xu�cȻ��$�?7��Ni��묒�~���3�U*�GG�Ǩ�����h�(�Գ���t�8.�%r��O�	Q�������+�����@i����Ө0]>l���;�3�p����+(/�C�т���1��'ʜ}�T�������L�D?���
�vJ<8�lȚr���D�ɢM�U�ꙶ/���%�\gZ�Qh<a�S���`��˸�U* AٕS�����v*~�?[�a�w�^�z�C�1<�e��1�t��T��^�A6�����ր�x��kg}������a\H.b֚3��oZtd��5Qv�<.8�����mP���nw�;��:#S���!M&�w�]��|p���䘤G�K����[B�_����f����ivj��d��=��,,������)Vͻ�����@��;S�ς����)�|��v�'�a\�,��ѫ��&���!ˮ�����{���S��j�%Bd�m47̨������?-�D��,Xz�|O�\lCVĄ5�<�7�p������P�F#���XԄGJwh�N�o�	��Ղ�lB'�xqS�\N�p�=�A8}�J�1@��	��=�|��iJ��US͸��}�C��jl2���;@�{����Bgʙ��������DO�F�vi�n�[����~4������a�	��:О��ɿ�x �i=E�mb���jE��h=a�;ٟ22Q?){+ �L�)�@����l���)�"E?��3?&�|���/�n���q�f���_�w��-A�܎��o1&&|�ꙕ����|�χN��=���QE�q����)�-���V/5G�*�Q����z���/+��Bz[���/o�p�.z��ն��A��ǌ�H]MC��n���#��м�*�-�<	E�ENf�K����W��������^�O�
�bڗ��X^q�z���x[��� ��ӌ&�wU#���e���6���^������i���6!����k~N����K�e���Բ9�	��������q3-���q}������B�����sprJ\G��!
-t�.�P%�Т�|�Z��xw�-��q�d�M��vB�@��g�)z�HD��Dj[�8a-�CQ-��!$���*�BJۤ4�Ɖ�4� T�eN�9#@v$�<]�~�#��Eu
�>��d�7���l*T��H�h��V�n���1���3ԍ�)s̰�@1�1��V^|��ڻbJ*�䨆�q-����G�i�>�bX�3�{RSitDk�{ݢ�H+�^s]s6~��L)`�VQw�:���:�_Pq.XY�aG���f4��Q�<�zFvӎ�V�Jn#yG��n����=��j�D��ǗJ0,mt�Q�d�vin�Y�A���WM�)��I��3�j�U�c���v� w}�G���RHXy㋎7.�k�ԥ���71F�f�
2Mgs�y��_����^%��[�|yH�'|Gڤ��<��ʭ�%�6���ƾ"�4�H�����-A�%0�P4l�q�(�=�o����F4Ǹb��[]ӊ�%҂����?��� Mع�
����Wt �5o5`D٥Ӿ�L��^�N�Yp=��> �x����_�X>�]\�X9��B[9/��[��U�; 7��q��hİ�{8o,j@�#�'�4�9P�@�zY����5
j[e1�K�<�}�waY��ڜo�0��A�;p0�@�YEK�-��+1�'lBU���}#��5kd`���W|F̬�P!.�����m~�J���R�x�y��t.^}i��r�Qf�E�&�bkR�ݾR'N&�U�I��I���Ao��-�G;B[�s�	|;�Ip����bx�f�D����]�UT�?���Y��8-���#�mɠH���<�7 ���9#�H��+8S_	�1�L@��,��.N~�6�o ��%3�/��_+Z��2��)Q|�X[��tǅ-��u���ju>�)�lļ;dwح�f�N�����t��P���x�j��X��-^�Y�:�~	P����`#�6~�]�3�qV�d_	�9fd�/�� {�F��,�:VP�QFvQv.�Q\�Yo�U��"��k�U�8���(��:��F��<1*�J���>=��S
���[<R����!7��{"���u��V|�x�Џ!���̽�T�+�$�8�r��1��ٚ��_�lE�V>��3�qo�w� (���K{� B��ȹ����(l���,'�:�_<�K]�II��q b'b���DA@oj�� ���m��%d)|Z^mA����&�*&((|~����	�(D�S�QO=���=����Uoˡx��z8B���pt81��B�mC7jq�Mޡ�,����}�ʯ��bnΔsLt`���Ě�.Kή�Y�8��\�������z��*|o%����E�+ő0ώ��V�H:B�aS>���nz��bq-[��s��ŗ������7��*��7���eT�T��n>��Iǰ�!��/z{�����MW��y�e�0��E'�M09i�� T9��ܞpOQ+6��?ʞ�߲�P��J�T��X�*�0 !�!�z1����̢��_3$	A���6��ʢ�SD�~�#�m�
�� ���[���Q��<�Iw� {;q�DX��Ǉ+`i��{�8���A��qA���[T�`�����3O�O����r�x��{N���������E���anA
�ꅽ��-�L\X�2���X?(�]&�HC��[���#��R���ʻy;�$:X��D�S@�
+"���;�3A���5+B%��5i��F}�����(�:�vA�ar�B�F�?�B�M�����b����j(�"���L�45�S� 
��G�i�5�cNn�xRF\9�������tV����H]�?w�v?��zMC���������n�d��M�bs��z
���[zqo �GV[hk�l8!e��H�94���l��I��W	����U%K��?پ�9��`���/^&���V�\z���=t5'�o`����3>�#Z����E�ϊV<�(P
�������er��6(y��*��Z�T �p�<�*}��}�u�K��6E��`h����%vbA�
�e��p!"K�����O��Q��!�wY����P�o�{o�.������U{�6� ��}�����蹊!�?�S�{xO�3�L�B�۰�z�/w��m���Ib F�]���KU�n֍���oo�U��q�0m��`F|Wj��� {C(R��Ay��SH�CZ�[�Kqf��Ʃ4W��m�Q�bI|�{c�CX��q��<(����(�ͥ�٭&IEc�#'ʣL���_c
+Axiw������W�^�@��~^���(�g�ni&��k���_�pW�hĦ��G��N���-	���v���/@R�z�uӠ��Jp���UٙlY�)p3��tϗ���$ �+��0at�;�\$G��r'��1�rH�	�^�,��$v7wp
�n�&�0�Y{�@�]��р�"X�I���d�>����C�ӛ]�ggl�v���d�a���������������m�
c@b2����D��O��5��B�җ�m�l��s�Q$Fg8Qgǋ�R�wvS�$V?M�[�Z�Nj�3���^&^1#Ty74��ePZN�)bQ����r��̻��)˴����ժ.]����ɯԻ�P�32����)��(O�M�;Ёx$}��c��W�\hB�P�IH�_l����q�u�^AnLu��96I�Me��쓇���'�皍ǣ]�$�`
#�c�|�>W�n_oa�<�4�e� y�cV{B6�����a?XG�[�j��{��NG�i��9@� g�1�V�{<���I׺NJ����a� L���C�xw��.�4��v @Z	ܝ���G��~T5��5���߉� g�n�^\����S-#zz���я-��T�b~"� � �k�� ����о�!+�e6c>,m��gI����4�����K|)�M;����b�N��G���Ƈ`r�5v��`�֔��:>j^�,ӻFUC��oH�}Ts�s�զkSA��#�9��m*�S���.��.��]��"�0[+��]|Vw��9ݦ�]���>#Z��%��B�" Up7o�(cr�~�	�
����NJ���h�H}ĉB���y:��%d�=�Pv'>9��B̹�
 � [=7�/}�xv��z)�r�\3|Z����	�?��0}U�m���M<�h���-J�K�:�����>�f3a����,�'�9P%`��C�&'9 ��X&��,�?�m�6"�Y/G��*� ���ax����}$��;�mE����g�g:�*�j�+Q�]Z��b�^W#���{��!�
۸]���]�s�3gE���p;���&9)�b�}+(^���5U�a��Y-�J�,�^�_���x<�2{�%�����\���0��b]�1�D\Lݽ����+����������@�Bӳd�:ⴛ!�P�i�Z�� Z�4�����H�u�'�/8J�2	@(ϬS���!��ծ�oZ�~�D5�w��1%�B�����v��t�j�ly&"�Viqj��?Ί1v�f�����CݳT <꣖�K���nX��۳��p���X·��h<b����&ϒ4���,����+��y�����YD��F"� ,פ�8[	I&��%�l�nD�ے�=���^�Z��ꥧ_Cn����� �U�0���YrzW}\�I[>�Z�tGz�W���'=�w�:Bv����2��i0!�WJ�v����}���!�'�����,��~�� �Z\ ��K���;섚������i;��JH�"0���2��\��-w�#��Z����A����2��T�Jƙ���� �:�?W<��k%`�N�s�m;����܃��b'I�$��ݔ�[��PoS�@SJ���(�����7���'��gm��PX��fitb%;��Ӳ`s���3ȁ��:
pB���������4�SB�Z����l�)��sh���| ����x�J�]����V�3�ǿq"W�����#�HU�,�Z��p��b)���e�D��M4.��GU>����!Kn����1[U=ٹa�)e0�dǛƃӋYo��``�yGl�����А�zň�����Vc��:���˪��@�K�*8�D�j���%1��c��\�_z��2��H`����c�HXj�����e��\�fhRG~5'G��n��L�������!�6��'�u����6���.��L oX
����bP��S
�P���)�<����7 �o�޻~��k�8y���R㏨QC��4L�s��08�x46�0��'&�~�*�X��:�6`�!,�'��|��G�\е����'��KE�҃�(�>C����6���
�WW�UTUnM򳥏 V@�? mu
�k�|^yw�R�pIx�xEMk�s��أ���u,�z����Ñ(�[샔ӂ\G$-5j#sNq�ʚ�,.:��v8��a9�'�v[���* [PI-Ԟ%p`�~'�%`I�*N9:ɷ(��
���������
GlU�[��&W�J�y��=����yw9��� ��3����dQ�Q�+xg�Jn+�W�D�ǹs:�Jy��G�<�����,�y2 �,Ӷ�k������w��m =�kn�/KkM)�1����t�f�i�����C"~$�ݪ=N`S���r��-��FL��Jf7����~ѱ7E�^� g��YM�
V٣x����vO?mO9D��U9iO�<��ebm"PI&A{S"���+��UV�t�N>�o0�B�wQs����C2�}�`��j	�|���8Z4�H�)��⼺D
��~/���Z6�D5U�;"���f��Vud����6�d����}p���Y ���p�=�y`|IkA��"m�`ί�]S����;#Z��=���^���h�/]`����-�^Ln���&���=.�~ť�K�2�Q�C�;�+�q��z��8c��nKPX��-�&����
׻���`�-0:��paV�|)��<@$�1)
Ye�a�����WLvᘫ��cP��R�1a�g��O�-Ov�s+��m�̜�{/�]Z� k.m��c�xۖw�W!ns�����&8��py�eu���@2'ˢ�f�X����c�/S��1�{�����B���/��U���D[n\x�=�E�9�{�ΈS�P�;��b�P?��~Е9�N��r dfЄ"5����t�+����O 7�j����l�>�
&�,Z���[���zk���t�є(cCĽZ1�o�(���_B]ً.����7��h�|rY�f�̷�����l.aε|4��UL�%sF��("�s��ݙ�z3�΀<��]��b&��W��ҵm͑��#�q�g��H��	�D����g�c�*��{�.��~��o�)a���7��=���7�۟͓v�	��1c95L�(���`�r�1d
U<쐟���������3�Tֶ�}�{���S�V�@�� ,�M�ߊ�
��k�u�x������ ��ů���|��C�y�Vp;�nNv	���j�a��ӨEʱ`�lȫʡ�z�6z^�':��,�b��e��ވX ��/(g�Dg%�6b �s,�S�5�1�8M�gz&A3��d�
�:;�#���~���i8�7�V�r���9��}̉`�8l�6��:K�M:�5�T��[ïx*���H�He;Hy���|.���J�p%��~�)���� �Z���B;?��J�~�>�}�i��d��)Y��]nc����#ڙ�
��%b�n�ʝ6��|�ĳw
�D�X�! ���P�gmY��7��-Y-�7y��~��p]�b%��o�Mb�8ןQ��ϗ�G�=1�:�c=�O�ث����F,�O�衔*��To���n��%f��~��^g�O^�|,�^l<�v���m����(��7�gfQ �e�'��4���ֽv��|V�J���G��QX��*�M��o�`�e�37�*;bֹ�H.�M]n	��	��9]��S+�q�D�{��.�f�s�ߦ�}���֨A��X�ɷk^�>O�p1/���,�,�U8��|��0q9�w�1�'�y��~����*�MkV��^�k����-03�D���6�T�_�+Qr�Å;*]V��w-2Er�H���{ܦ�S����e3/����`7Y��f0��;QV����W�����.����'�w�VOܑ&�!�q=wʟzJ��g��[F3y�����?�F�C�/Y�o���J>�y�*���W��ɔ^hܹsO��¾� ��8��V��]��-�|N�O��ș�t션��t��;4�H�ߜ�:wl4����.&�����gH^ @��d-7�S0��Y�h�_`٣N>a�vA*N�q�Jq��dN �=�,Ⴟ�MWMq�v�u�P�M�~���G"P�r���4zͦ������ʛ�ɏ�����ܔm���1;��9]^�U���ݡ��{������y�V�_���QX�˟�]�'�P��y�&�(d�Q�S��F7�ґ���\;��@������NWV}�X�N��/��
ܰ�!�,T^Qio�N�jUZYX<.w���VT�G��(�M��+�q�?!M��_�� ն.�����Z�d %��+����֯�s����>�w[�`dg��Z?$D��y��T)������3 /�M�"�q��VC@����oʱ%���ζ��Q�`���-3�T3nzu��1Q_6���D��$K1���j�G��Lo�o������ӝTȿ=,X�g�f��u�gA7�;�qZ쓬�����o�Y�ROU�ڒE����t.��|тt��1��oX���m��y�z-DS7�%�!}�0�����GqH��_���K.}�q��?-�B��Уuo����>bv����R���ˀ�B�����#�(g;�I݅=C�9��.�p�/=r)��TW��$[�&�5Kz/�&(�Y���T*�����T3��`���J̼1ߔ:��!���G�p�#}����4�\H�[���T����y��يM�MYr5�� ���I׬2VL�j��;��xTW$C��Ve�l��z�,3�8�:am|v�➢q���P��}�ٺ�]�`޽5�r,	��`�{���aI.�����@�#�=��D�]��m�&��7�� ��[C5x����т������V��;E��|�@��t�� � ��[4��pQn �4��D���d��L��e�����c��>X>5�U���	��w�r���[�A��;��e�|!S�(�O�MwR�n�h�j���V��?��L�d9��a�eO���eʷ%�'�[i���':y_i�eY �=#���Ԃ�L+2;��~EkH���[�
�F�9�g4�Z,^qY��i�4P�.�Q_z��ھ|�1�Q��!��6h�[�I[��XSj�НA�'�ũD�r����M9pɝ��#�
�\ԧ@SNѣ�i��ƿ����>>�C�Gn��"& g��t�ˣ
?�����q�BG|�ܕ���,�&uX��&��
_N����r�/'eU�EL�C�M��H�q�6�ѷ���B�.����%FjL�6cO+$�>Hi&�z���s��ٸ�~#�r���2�]��_�x�>P���9������k���ZMXWY��&yPx?P��M?���5���!���A��+���^?�Q	^c:�r	L���Ɵ��Qx?��c
C� ;LY&�
�4G�hy>l:��N{ZR�XC��_b��	v��Ǭ9�Z��v�9^�o�6�G����_g�keb���M��n�k�H.�{��~�?ϝ��3��D����1����.�I�}�5������d�������G��tw�pYw/z�\�y/Dx�4��0ᶫ��H�:�W�	V/���gl�f}�_�U��ǔ�T�;�iߐ{(E�ld7:�����_��B܁��� ��^���ó�l=|�����C�TP��ki�<���Ӧ˱�P�Y�#`�k	�G��6V�ɐ�-�.� *eV�x��D�3�G�z�^r���LT%�Q�g��RR įq7�˶V++qҺJf�wL-���D4`�ÜGrg��[a��`���^+}�O|g�5�أ��m�h7���Ky.���G5 ����𐅏}����z0�����K�+=�/w E�U���>Ӷ'#�����+ �(f�CI���oD��Gb*R�̕�:���Cx@p]y;h~Q^"f7�]��I��w�6N� &Sp���S��z��wEn�ź�M�Պ�������l���ڶ�=�ԛrZo����L^¡+���[�[���͙/�r ���8В6�JQ��s��BB�7�ƾ��{H�6�)�K�Ec0���T}0T��mԃ�R?r}K/OnE����U�ͦ1��x�y��C�xGF)�ٕ�}��R2�?�+��y�8�a��	!#���!���%bS0��FB��(ؤ}ɄTˠБd`O�M��B�
W75i�D��kk�wR�H_�Hu+�<v����(��%\&R����x�5�U�\��icN*�z6�p���a�XE߆�������5���@��v�(��ź� }LjC��!"¸j�:��Vx�r5W���w��
%��X1�!  B��������Q��W�u;o�2��^�(���^ò s�Q[� ���|^,ۄ���$���� �]O�c��}ϰ��Օdt���SYd<񨐴�k�ɿ�|r�"��~�\)vuu�k�cZ�H�S�����0�gD]��A4�@����b���slQ�A<�@����8������.�+V0v�kh�� b�j,a�'�'Nr#6-�X"v�>"��kBN�6�H��=���F]��>����m�C����4�~�aD�b�����k>��y��%~D̮�OU"�J��	X����~`W(<-6^���1�Cz3a]��ϫ*�������5
C4�(�>�7�Y�[�MRi9uKv.3�7����"D�������{��?[�g-����>9(.��SĔ��+��#��@t��$6a��=k������,��RU���i��}�Am��[��M��B�&�ӎ���.�@��s��e�b,/�w/k #��AA}�C��Ң`���`�����1��p�
nF��!�y{��\Z3�H�+���N��K����N�(�j�4Dȸ�7��^�	�TiQ�S���!��?�Q.΂MM�G~��L�x"�1t�<�!Y�/���|�Cf�����xPRI��z�X�d����Იz�1v��w����J�������� ����K�E�s/*�;��Y�X������4�Z�4�v�#��`rC8��#�5��H�H����o��mQ��ð�χe�`��sov����nM��B���'�"��k&L�y�t�%L(n!��1̦KE�^Z�Lq�)���f)��`�P�w�h6���f\�.��0xwQ������|����`^����
��<����Y����}~]��k��L)(�=�?8d�!����{D��i������5�O�%F1b?ܪ����ӱ���6K��j:�c��s�_U����:���9Xj��RF%�[E+�91���т���X.A�Xҭ��#%��y�����˽�Wﻑ�UF��sJ�N��py�}\9D���<���92I}��0 ��<����[�Ѓ��������dW���D�C���|��<���BU~l0���� C���Q���6�ݭel�ݛu��ږ8+[�@uC@)%Nĉ\:��R�8)ה2ty��V	���6��Y���4��Beg��N_�����]��s��f�{Ҵ�̶+��dO�n2���a>�Q=2���6n��G�h���
>b-��mB�3���2*3"���R���h�Y\�󎰝������)���k�m�Ĺn�Hl� (����L9�������AeT�J�C��W�9�Ѱg(�Z_%���h���Wڸ%�.�����N�uhѦ.F$�����"��{�/�k];��~�����9"M� �0<Ԁ�2��nQ�t}�{�bO*�8np	M�#��"�m���E����3��1��`/2��)n�{Q�!���DFek��I��w�z�>��ˈ>���u����Z�x����bR�6��ڢve�)/����bV�ү���}&R�S�d'0fR$5q�yn�s�m�=$�
K,.�er�Tiw妎���í�2Bp_\�A�A�rT��VU��b���	}	pt>�$x\��#VBm�zȫ���6\�|p���TJ�����6��q�c��O��w�<ExRb`!�����	O�7���3��S�[C��5ej֠R5�%�~�ik+�����8�����>K�-Ċ��dԑ$kZx=T��q�u�F������PA4B,w�y?�áS쬙��L���U���!��ƕ�[��Q���J*\䌿$���� �N��;=�So��wFi�����Dv�%��������6�V���9"N^���- �ʶ��Wo-��i�.�v��ٳ�\6x�$:$<�y�eJ����{j}����̯ۘ�0m�D�o�sN���y�l�4�¢vo5!4�Q������*p?�F��:q��FuZ���O-�aT�Xޜ�ZO�I�ʔÈ�2c�Ff*�ͭ��/��3�*Ö����@ƼaZ�'�'�G�D�xn
kY��Cυ;+"�!���jѾ�VJ�B�t����(��6$/X������̙���S��q^ ��p/�.2}Ö	�D�Y*gt|�(�}�D���C��eϢ��lm�^$q�����Ȕ�G)L@^ћp�c-�@D� �V�}�g ��Q[� ��"�r.�����BqW�����H����_l��V�غ��0l��/�ߚ�� x�\��@\�v���� �`��'����T�pZnb��>:�s"m��c�z��+%a`3)��j�����s�=�"�ϣ#��۟x`#_8�f�H��:ꓱ
�x��~(
�H� b�]rd��_{��HU~ĺ�5��������ق��T�DהDQ�雑��/Ch�Lc�C�Ŋo��9C_Z�Z���IT��7.��dM�YƑu`
�J�#��͕?�5�^��olvս�('���K��|�)dT6%A�%�4F��D�f��f�		p��&({�"�����g��|����"(�wn`�rf�w`A�54��H�'��q,U6?k�\��n���<J# -�����B�u�^=�Ԭ������
��+9�[7�#������D�+�l�ycK�]H�̡.i̷.FC��˛�X9��T2f���|��j�]o=0�L�1"��5�C�s�� ?�a��PP��'��7�5~5��t�8Z)S�}˗ݎ�,�Z?��~D-����83�e-
`!������L�P��҇k��f`t?[:�L"��PF���bҗ���{j��}��Y�-����Wn�&^�ǟWJ�4g�7�����fZs�)9S��
�?5e�@��J��J-��A4nQ}>��L�0���1&�F�r���M�)��D>f�u< ��x�=��ȴ��&:�i�⩇�y���������(�(І3%t[����]�
Џ߯����'c���W�v�=*M�q���x��!����W5M5cK~��ɧ�=�{"m�����Z��l�j9�F~w�B��^E	C@� ��aȶ5�;�_�%�\��Ut��ǠІ�ی-8{ە,(&@�	A��d˵�+��~���D$8QR}�FG�fԿ�5��/�e�C]s���w�ŧ1oM��6y�~�ed��dW�۪ܮ��[*K�~�-�n!�c����T0�Z��5�zl�]I7�B��,=�+ZI NE��T+��YvD9s�Mە�� !&��O1nW��ɐdBq*�#-�0i9H�U�#�1Vi#�^����_�|y���!w��l֭��CT؀ۑN6e�겅�bGI��8�,f���.���ˠ�pI���1(�{���fl��;�/���c�a<GB>�l9pL�ґ�u�gT��b�M6	bku����l���{��6=�!K�*�_��p�J����#�tv����($oED&Ȱ���u�H4Ȝ32.n�Q�5ÿ�.JLp"�9��\[Vux&`��� ��K����1,�e'�x�\Y�Z�'�x�"��3s�r�'���N/�K�R��b�}��m�b4���s������R'�4�d��,UX�^��X�1wU�꒾�a��]���桐�!�@�p2pu�m�|jN_�BN�i��F��'�r�Bt��I�;��}����^��0���5[�37��C��U���#1~��H�";0�ٔ� a��I��k:2m��J�'��x�lG����ϑ0._��$B�`��'p�^-	�q�V�I<��5kԱ��Y��m�T��:��I\�����F8JL�aH[K�� ��=4��2���|f����aP�Sn�d����P/n�VV�d|��� ���ʤ�D���i@���ں���񯄹�ᙤ�y����{�u$�+���ɂ�ܽ�����訴�1<�l�i�̗���ju�H5����$� �(l�ߦ�՜���S)K�`�\f5�/<��y����&%�}��~��7x��k�N��	�=�P�I���1ѡK��Jܹ�ƅi��0Y;$�ZL��Y�' 1.f���3�q�_U�;/S���v���vm�~r��)u���H���j�4���Q����\l�w�@&�~P�g-���N�ό�<�`��Z����{K�%St�Gݾ��mu���� J��7���� ǔ2���"�����y)H���j��b�?T�(5��dAF��ًW_u��DE��=ӡ�(�~�@�'�o�N���6����Cwj{èSB��e��Xl0����5"�K#�+~���G�B�~q���ɀw;r: G�i�b��$wSt��o��WN*��q` f��B@8<2����3��:����R���e�Vy�d�������,������͊\#�͝������=Hg7(u+�-�l��t��zaHw�c�̇�)�i���%�K慆&�]PL��`�`R�'sv��}�|:U��ِ*�0%�+�+e�m�!`���me�=B��D��r
t�;��������7� o���I�ޞh-�S(B
ƺB�z6�,�f`�s�m�EK�n2�0b�s|mY�Uye���(/����4��r��l��^���:�>�z���|�v���aSgU%:sa}��޳�9&�F̗yy�[��]�PC���z4��z�k��02�*#�b{K�^��µF]��|r��FV4��X�����i�&��*�O���+80�A�~G3JJE��\��Mƛ��M��RC�xm��� 	��\aeJ|���������)�I
�h���ih�
�|&�Z[�����<f��H0���.GQl��|o�ҙ��շW�9g�-)eZA��2�/q:o�c���-��Y,�ͺ�V�i���!�-��}E�@�ȹ3I��~����b
��b�y��7hKz��'�+g9��Un�[�4Y�\a3��H-�!�e�~?�ՂcB�[�֬ss"�1*[	�7]ے�?����F�ź�ț�ڴ}*��Z�/c���,�!<�XqJd�@�M�^�Ђ�	�F��G
�F���s�XށC�a�%=�)��A�L�5���Q;D/:]����L�Fx:�]��)w�r6o���/Њ�)�#��v�T�����oCc��?����S�p�0�^k�G�ɓ�oZ����g�Ъ�m~�q�F�|��%��N�PJ.%v���0��i)�&�S/p��eՌ�#�ߑ����d�P���Y-J�VAj���;jW��L9�C�v?��'�ػ�C�Ԍ/I�����|�<,ccf��ǣ�I<`DCF����$^��%�g�6Aa���)*�f(��hӃ2j�NfW>\��=�*HOM�Ji���di6[Yt	l*M��p���/��Y�	�(��	`�s!}D�Y#�/���0>�,M�r	�Z`Rhf�5��0|����������&��@�����} �-5fc|~eGJ]��p�=@Vpɞw����Z���#�%\�E`���ã�']���&�OOk��vW���H��.f��-&ŉ5��m/��ihϋ��!A`��&�T�<V���
|gC��X�8�;��	XnH�#�E�D,�~���
ƇeY�rlq�[<
���y�T~����Q�@�W;����5Y�i��\Ä��^��~�N�����H��7M�2d]A��D�ڭ�*z|/
j����jB|��J�pz�D�m����NC�P�6��Ň��������^�n\R:Uq��(�=��6�	��� ��)v���pa>��¶o��+����QfA��G5/��3N�?�&���������,s�KK�������v�;8y�/��=atG��2�l�Ͳ���܊=�������š��g�m��Ur���}� Mք7#=E�R@j8�r����#
�qCR�`���7(����e����(��%H2S_"�߽��o��8Tr��|��q�!����7.>�Md���sh� ��/x,<����~}�����<�T�
?tyY;��_�G���#��]�&���iIV@4;hG�{��D��U	����9i	-p��
�4Kag�����i�����RU�L��s�j�i�U\��,�\I3�J��h��ϋ�	���$%ۊ���9Щ>p��6y�����/ ��O�v��䈯M 0�����)��h��On���I>	� �!�������(�H7�-^&~��bvC�%ꍵ�����~l�06�i�
p&*�>�����$�Z�"�_��_�K����e�08��
dNP�$��?�2����p8*Pѷ8��]_Kw`��M#Xwo5N�����6�gy����X�2_,�G#Чj4_���iA�+u�2���vY����g=8�g���L^�����Xf@��c��B0���]�k�k;�5��&[��z���RdԟH@M�#����F��w$�w����e��s�+2�.�c>����b����4�]ya!�rCZ�Z	7V�5��-gd���W$?+��p���zzNX7f�78�ltFC��ZJޘ�]�<Hnb���F�<:��CrIO_UHU�@_S!C�O�B��������It���\#?�t���(c���.M{�8�eح��Ve��R��W�Ƿgi����H�~��L�dLf�^��wv��n�m����k�ã��R��4�+��erjK��+]f~|��-hi���#vV�ՙX�R��V���a߬�"q��ɻ��?�6Sw'{Yc��*�2�W�J������Eͫ����K�74�����<��O�bP�v8�"Ì�B�@:���DX�m�Ah`(����1�z�hB�>��+n*[^P1�����!|�VqF���N��L�4����2�cTJ���-LV��S|�67i��e �<��#���*h����`�J*L��uP�}�@4�46�Y�:�G��AV�x�tkΌ[:��b�:	Lw��xE��A)/�5-�"���޴���9�	;�������M�I����"�n��)�A�&͝����n
EU0fe��ޤH��]īO-sQ� ����0�F��]��[h��t���#krHlߪ�@�+�ȞtԄd��3wX,	+��zI� ���=��t�>��;���� ���&�ܟ�\!�Q<�ɷ�=:��C 5���u|�/�"O�O�J�4Oç~E���N~E�G��̼��%��~^�$��%�;�PrY.�_��]pfB�zS�G���Bo�`x�����^��X��7i[M@P��!?�j��YU���0V�;�)�x��S��}���n���sM���quA��41ʵ҇�m9���k��f�g7��q��Z�SFC>��)<J��N�����$г��k�ˆ�@�Ε��۶_-FS�h�Iԍ�ۮM; �����M�+���q�Ȱ���>�V�����r�n���)�w�XD�/`E!�)�?��tJ�[՜���#�Y�'�3��?�zs���O�s��Y�/�k����s�V��i�7˴���MOB�𭮒\$y�EW�\no�n_��& -�,���n��dK�� ��,�����E�g3� ��S_e�䔺�cʵHH��#����m�@�uF�|��Rn��K����~j�%h#���L�8s�₷�i����h���u�$�d��H��N��^/%�S�4�H��|d���2����PIĎ��&� �폷�3�������Mqn��3�dE��Y^�z}�F��wcl�}I&c�L�鰰�F�a'u��2�k�&����
3c���|���ȋ���Ki�׎�d@�y�h���#n�w%I��/Jf&k�����酮wF��ә-#
�ZL�Sז�M���V���d8m9�M�\��P���| ͵��%��&C��K��>�\�q>�W3m�f��B�7L?c�X�����@S�%�/�~B_���<�B%X����l	���Dei�BMS�2�}q�ز�7��p@�)���%�m����YH��/ޤ���g������%p=�&����|߱�:�m;R��٠_��KJ(85~;��*p��M��Jx�~�����!�uo>S���M'���:eG�.���q�8����Jh��Z����<���\a�۸+��y��]fעfh��*�یڑ3�Fg�<���<�J���?�7*���'����Ex�C�5p�O�-S�'ݝ�T}������c�.�.GQ5�:���o(��9���������
87��H�\��~�}+�he���/��Th�J�tD��. 3��{T�w��)9��h���]/s$GCBW��d��Az�):�{el5�j��C�Ka����m�+�̒��x-M�P���+5�Y�*)C:�p��U�3m�
���.��
���)
�g��,6wrC�i�A��.R0�{����H7�z��N�����{�)���c+�"��R��(@���U6��x�SV��;��w�ׄ�%˼��]\1��A��H�A�H�L;�CH���*>a��_e��$4g1��ĥ���6y��t,: