��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jåا{�\�u�?߷�dn@6�zf��r������; mt�M}Fq��(4C��-�+����ɕ{�q�>
�����*B�1�۟)���͘��À��g��W)<���IGcu$�k`��Z�< e�k�	�����x�Ĉ�د���q�Q���p?Z�jآ����e	J#J�������RNK��ƥN���1�k�f���C�, ��jû
FV�ny����*� �B��_�E i}�M�u�sO��\�9;�ͻ5M��mϠ>�%cP#Z�)U��.��Ds�5�e�8C�bm�b���;)۪UN�����z����RB@(~�A�#Jy�h|k�5.��8�������n&o��_Pߤ`�E��2�Y	��Imp�r��Q�*#�7�W�1Þg���)H�Ǚ6��F|v�I��%jğo垌|֗9�d��g�cP�p(�T�F_����9�"Ţ��<���;S_n@$2<5M��R�H2tF[�Q;�D�8bf#8�	=��[����]yw��pГ&G���-R��t�;A=�����X�f�����du(�BH�r��e��_S��ƽ��"CЪ����_�~ �y;�*'.���5�g�P�ؕ;XD�M�*��z�!��6�#~��[k�e:�pK�r�ff��{CpLB��Z �HuQ�`wDt� mK������&_��Q�L8zg�aԂO�v[�����bU��1����G��_i@�Dj�Y���ƙ)��LU�k����Y�@�^��fQݬ�M�W��;>܇�# ��0�D�a)�P�8�~�[���.�q�"�'���/=i�oq��ځ���?�]�,<"h'��H��~��Y�\ޭ�9��� ԩ,���}LDn�k�~�Aȣ��L:8SYǗe���p��v#ȫ:?$�8��\y'h�.}r5�8���Anq��	�}�d��>F��q�UyW.�^m�����V	Q 7�s�a��o[RH+��ß�(D=@�gC���y\�8�16VđU39t<<P�x~3�0P�Js��ť;��k�4�H�%�Ǉ:�Eؙ:I�]p_�:�����o���Ԡ��M���n-kW�{K6�L��o�1��K���Q!Ģ�B�m���S�͈-���0���?@��c���
�r��y�b���XeR���^�pS�6*�w���F/���aä|<-�x�R���vLF�ᬭy?��ʋ<Y��ȳ�j9M��e1�S�.�|`��[V9����1����t��H��RQ�6Lj�9�E�v�"$�7��,y�V-�b$<q0� �1����ҟ����c;����h O�r>�)�ѥ\�<�k���� �M��<#��B���W�����+o5d�s�LVͻ��~����s�d&zL�B�&��2�9q���q�&�G�T�K%����������O�ϱ΍�+[Ҝ�2
!5����&���[C솳���6��@�:�b���mqď"�=�b$ѫ�䓦|�+��X���Ɩ�֢;�{���w~K^�f>��>�@�4����x� p[7����"Hր?%�-Z�m��]�Zڎ8(�S��GnF˕/j�13�qy `bx�v����]}k����S�P�$q�
���29H����,A쾸bg.cX�����d�{
��>��d+]<�ײ.�e��1���������m���q�׾B��Cwz��0�i�Ie�Ʋ~�3���u/������T��,��Æ'z�i֕�_S&�KH���t����Gzv&���<�^>'W�Ǻ�(�R��~���3�ʹɭ)�9�y���3����?�o���Wܽ�!xB��7��4,�I��0z���!��P��JM����6���l񢏝)@t��#Ծ���:K����� �*/��4����3���0x0Af*�p�G�t��h��,�aI���z���>551�ૹ:a�Rj�0���'Y9|Ϊl����Z��yg�v�6B��UakwQLP��T	#ܻ:+��*��l�@]����#(��@�U!� ����p��Fe$��߅�Q:�Ė�yH&-�z3'u�(� �}!�{���g��!��Q� ��@[�S����zm�~�U��b9"���4\��M�b�����z��h��NA|��u���g����nQ�k�-3��|���9��q�FÊ?!&D��;����l�)��Č6��\!+L�.�L��}۲?]|��޿��>x��LУc�`����֯�l}\��br��(��bxo�l�wj^eÂ�t�,z&���U��'�L��SFw8�_���)MJ?D�ī�(;�w�_H��s�MU��o�+|#��w�k��l�,"W��v��{1X���/���"��	/����~P��e�w9_O���v	���Xy1�C�0�}�#�
3!�2��{�ҙ�b	�S�/&TCy�ِ��,F1�fz°�;J�b�tmȾh�7�tR��Y��/eƃ����t��{��^H���i*	��=�������]NQL_6��J+�� (X�)3'����8���!��(%�kݥZ�uN��x�Mqu��x�F�nbfAW�Ž:���<N�{�=1Y�<$w�4��]�^��Xmd�]�]��I�g��K�}�[d��x���L�O���n"��{����l��hV��8O�t�\���"L?qxE?db�]��݊��'b��Ƙ�ty�m?��*��p�^��#栳�:�輸f�vqz}�����	�'�]��f�yk9�{4�0B�2�9�t�����55(�.4�T��w|�����F�B(�`��eQ<f�!ݺ9x���Rm��Q��p��Z�[��4\�dI����wڷ��[�����(/Έ0���G��0r�Z�����Ţ��_����'�*^4Y+�qѓ\c.��1Y~����I��K@�G�gxa��>pu4��`�Z������@2i�7�Sr9�#_�f��О�QN��^����*J	��EG�)���q@����L:�靺�x;�Qඨ2��=35������ު�xz}{�v+S�Ѣ� o^O�&��PF�~bQ�n����<(�q8�$������NU�h����7�]�	�C�t���:�2����}B��}OUnž��A���-��A�A����t���vMl�\�$�>:a�X[Ҋ�M>l׸����KZ�|�P�͹f�?��<��c*U�H�-�ԃ���02 c��mO��P_��ZUH�CV���g�"��.���XGڿH�bran��?b�4x]�ǒ� z'�+qTl�g�uH���� &���/�ZX�{O��ǭ)B����32w7���Pa�w|Z���]�`��D�+�Ğ�o��9���J}�
�9~�}Ԥ�r|g�����A;�`)>I�-cBG�z�d~9������G_�*\ �GB���-`�����������֊�I��NR��~!�rKH�
�D�{Ro&�;;G��	��<.L`��1��?�IX'�k#����?�(�R��mS�Dq�3�N�y�<-���)��y���׶H�Օ.;��ҿ���˔=���>�ǚf},�B��J�A��Q`2�C�ɜ��'�;��ƙ�g�0������`��x����آ#(�ko�������S��&���4ٙ>`}	/;]am�mЩ�_��B�<:��>�,'q5�:��.�@?���ΟSL2Uj��ăJZ��2��d,X�Cπ�`�Z�*>~��}��҇�U}�(As��t����!��(�i�L(�\|������/w$Z����El��i ���t��h\�J(+�M���TH���+]�������c�*�i�G5�(��6��b�����ED���_�rj�>~F<��!9�6<�����o�~�N���b&x�h'꺗��B�p	#���nU7�hK�Ф�q[��"�� Ϡ�������X�Rb��;��C��+B��Ġ +�h�&.��Z�����&x��;��FN��nλ�!,��`���k/$�z�g����ǛW�9��]�ҕ���۷��\R6�y����v�"��x�<���������8��C��*�\���w�h�{l�Ft\y2O�i�A�������sZh�1ژV$�\��K*[2��,���/��V��[�	:����
̜�x����p���
���I��m��P�dr��?��p�!N��7�B�F5G/���������\����2�K�_V�^������{�^�}��#��/[L�ީ�
����[0� b�NT�ш�#�֠�ܬ�~|����Ul�� )��58���K�d9kLP�/b�'�Ŭfylг 5�eO���44�܋����CX�yz��� %Jܖ�Qu5���%���5�$}���q���m�����5G%��p͏O�U��Ņ�5�����8�̾���١R�\��;d-բ7C,+���+ε�<�:ʕ�*�*g)���m;�F�n0I'[ނb��#�GO���:��I�������\����x�CcS5!3�"�)��[e�5z��^�� �0�&B)0Nb�ɱ�B�VA�����f{�,��-�*$��U��h���)������0�z���?����4�v&���T�(R����6V��券��R�n��7Ly�`WںgH�׌y�����=x���� ;(�GXD6+��t
-�l��rK�q�}���."��(���|�A�y��P�������������6�P\!,�?����J4����|��{��M�ԑ��m�*��^*ʯ��@��Up�"T�:�� 7�FG��N 1Q�h��pS}��J�㧤��kg��U�������_�o�-,�'�ACi�ߝm����*��|�+)�%Ƚ/'��5�|�yc�:]��u�蝱0y���Zn(��D	��J�{�q���qt&�2�V�O�;�;�ԫy����8߃1��ދ_[����PP��W���2�����!8ǈ@c`ud�~`�����S�W��=���9����^��4bR��OBw!�I^�a¸CJ���<	0$�z�(�=(	A0����X�-�UnU��^�Z�0�{B�'UTŋ�T��}����-�y���e�a���\SV젭4!�b�.�$�Y�ըh��/\"+�c���Aw���<�������/����i���8#"�dY~����4�!ʖ�H�.�6�p��5�k#����������r
~���O:̘Rg�����N6U�xF� FM�k�?Ώ<2���mk�I���G�՛�n4 ������D��y�����$:���t��9@�0U��~;�XG�`�M�S�+�����
.�N\_��	�nq���+FW�Cj���}�L�Ry?>����7�ɵ�{�67]��J�}%O��md�|�C��L� �f��D�i'&}+��1���5aLa�	ki�9ނ����t����dGg�"*?�Z�
�"��=b��-PdDM�
u4KW�T���"��L?_{Oҡ�ꊡӆ�Y<��ʎޤ��⿂��-Ə.l:rA7	���6�e:R����X��W�E��&K�H���f�9o��ԚZ=��[˸��]�gLn�,��̀��#%4�8^xe�'w�����M?Ӳ��|�g&�ten1��(�u��+��F@@ew+�]��܋dj�y ���"�m!q|a��������ٸam��!#�k��+�MI�~�Y'k{-�|�ʫ�Q�}A-�ô���,�S�_�C�}'�{s� �5W���g�Ɏ�����KhNR%��n!����}�lrb3��K薞�%p�Z���J��#O}�~?��ʭ1����8Ԗ��'�?���{�."��eNy����D��Q���ɻ�����I�|T��W	���3��V����'j(�g!�3^�E�`��
]�E\T)p�g�'��Ks���ѽ6�E6������� �ItԨ;�.lԜ��/�9QG��+5B��R��2=.NZb��J��/R��#�%�c�~c�͙P�1���J�;6Ч�$�@��r�B`��L#�:�E���`����d����� ��A��9;�l�[b��5�)�d��q]���3�b�P�+�u��A*�1!�hm�`ϲ�}U����QX(�.����y��{�����8��g���ʒ���Y	se�.N�w����c��|fצQ���m�=�J�I��.�iZ��p�YM})�闍1�FZ��?A��z�=�[�l&�l	�E�aY-�3�����܏
k9�U�B�q	޲!���-j��}>���_!�ƚ;����1E�3�ރ,����0 �C3�����>KZ�ϓ����+�OD������W�Z�7��u�4�7wq�N�@ �~R�:u���􆻨~L:m~1yи����Xa1\&�.�\�l��j�;ʔ�E/|�*�W����r�}U�v��j��B��l���2ԏ�'3�����{b��c��X�: ���ZÛ!����װ�����OK�����.X��B [��K�$�\�dMU�
ϭTǌ�b������������a*�1�n�S����6$�ȧѮzHзBH�tI�0٠�:4a��ȏ�1S���q�RY�o�P�5���P�h�Nqp �A~P�ĳ���׷�D'R+������F�n�B������{׬>�{��Ja����ܱȊ����M�
�-Ȍu�+[�F׆ zw[HBc#z��p��M̿��G�b��mױ�Z)gj�G�9�hǵc�$#�]�u����^���3�����z���E4vR�c��Wj�Ip���V �O����b��_鯐���Wha���l�(*����W�$
M]]O�M0l�6�r��U�7�<Ig1!YE���WS�u�	�g�
)/� }Jn6MfR����L�@�᏶�vJu�M5�|�sJ�:8�j���� �[ZA��m��vw!�IW�:�4�s]��f�0��kD��Jq'KK����6�j��}zh&j�s�n�ZQ1� YJ��J2�CCVmX����~T��e����
dL`&d���>�����f:7n��d�ӓ�j$te�Rtc��A�A�K�I�V��_��{��  �[B1'꠶�^��ߝ9��l( ����
��n���`�h�p ��S��:]��ǫ�v�QQu��@���-9KI�I�i�&�C�
><�|k6_G�F�������>6+��o{n��Hט���{$$f�yN}�^g�W��4���W=������Z�d@���Q�c�O�d.�@�H��V��)��n)x
��V{/�nU��DDV���(���Ѭz��.t��L��\r=�nj�5���+R;�je�̧�5�	W%�\"�4_/�"���y3R��3�p@{r�bܳ�ўQ��h���w�G�b�Y+<a0vɡ�a�y&|`����b��N����op<L?��tԂ��:<k��8��-}�0OrH 
�))�_��y�˔@ҏ�������tWS�����i�gE\�V
��_�ЊA�Y�
�HP?�J+ѦQx�����7��	�|���Ǥ)
�F]��\/�׫��B�07�#{eȂ��.�{3�k���/JFO֜�8���$�	��DS���5P��K*�00%�У����7�2��3+�q�R���n���^��LWV��h=A^B4j	�j�����yT!Ք�K�KP�\��4n��C��"�v���'=8���+o��u�O:��&��R����򜈐Kkgx7ͨ&�c�Ե�Ԑ���o�"|�q|g����5�OE�ѻf����ʮ]�$1����8�o�ZO�W"9+�%W/\$r��ǟu7��H���>�h�5f`��V����8���j��@��*�������b�� �Gl���J��4�$A���\�Tx��c~˸�#br\��qE��D�DT�x�%q[�B@.z&|�#5�� �[��F�ҋ�}҅v���ï�F0~x����
!�+�A�&.&L�w�'cj��N7!:
Uff<����L��d��s�+}{��-2)�H���6T��4�`��+©�S}&ԙ��hny�Ǒ�b���N���8�,N�*S8�`{�N1�"�!�I���
P>�n>q����jl-Y�:�sJ�{Ġ�o'�Z�Մ�yt��ޛ>�u-�M|������?䯕}f�;�0���Q}B�`���H|Z�Y��6ꎇ��Z�9T_���?��X��S(�4������>
�96�W�ċ�V��N���B�QՑ.L�v���U$:��� ԅo�ժ�5�#5
ؙf����� �@	j+sBCn�nm�6�iՇHF͘dtE3~���5:�?j�@oN���Y�=swAS+�c=&��ݡ}�L{@p �������p�Ҕ������S���f��Ol��N�L\�G&D��}=�PH�wB(�ɀa��˂y
��M��#Z����Z;���T��6�PO������\���3Û�eF �ӷ�E{Y#���D�N4��Nk���x�v�s�C�5L�� l�U���%^G���j�9�w@��0M�t����P|Hf�-Q�J�Ӯ�ȷ��az�~F��+�d��+r/�e'L"xG|���w�(��7� Y�N�g�+�kx��$�J�ʴ0�.ʉ�����0�g:,������{RB�"��t�a��k��`�R1�0HՂ��b#,$���p��M~A��;�������Z�(L�{(.>sE�MmҾ��Xll����o܇Wa��/^��	����ST�R���Bk{���ӷ����F�Q�K�5n�����e���9�{Q:��.uȧIA��
>�ة�FD���1)Z�5�ֹ����$\//�_�EC"�B��{�ei�KJxXV뮇uNJ1t��A�KM;���_�6T��i��+3&掤�G͆2�+��aC�ꟽψp�!J�2 �l��R����i;>A�	���cNY\�̵osef����.���B9��u��R�X�UvØ�Y/	6k�a��7��ځh葌q�!VG��*�Yf�D�~?�{)Q�k�(��O��k��ia&��3R��H6VbQjc͢'�ބu��j�~��\�4#�n�Q�0Y�p�B8^��eE,��M[�2r����!���������XQ\����Բv'Ÿ���?��uqKwe(��edB7˥t �|�`LI��"�B	�K��
ݻj���Շ�Ψ�Cjr
Q�	��#h��+������&Yo�e�6{C[�Q��fr?W=��J��!��/R���E�sr\���0��KT��������7ݹh�'�`� �$:����t��M�]}c�J�4�iY���[�n
ʦǄ�eĠ�
/� �^�
��ij�B��m$�f�ں��_o�����Dt8�v׵�"b�:�3�n��m��Ɲ�r8sv$�������G(*:'�{��oe	�2?H�04��w�J�<�����\GR��*QI�v%�nfH�K�d��s�5�ݓS?ՌB�3ML�ig��P�7�@)m����8b8SC�,�4�� �=E�xը6b�h����'�,�� ��{�&&6�*�B��d'�X�ԃ=�e�8*X�)b�TAB�eٝ������UR�&ބ����]w�š��+�n���˵u���@�W�Ʈ ������u��-��)b� )�z�E@� �J��;��t���
��>�s.����&n~���F|`�]���2f��\> ��2�a��,ҋU�$F�T@���∳�W�5ڶ��z��K{pG<����`[I$�aT��=��������!7O,j���yrX�)�uL���Ox�zJ(���s��|��O�VU�'X���B�g�<Ɣv��I�z9���������0����\�^ϥ�4��u�UHU�kH�;�$�ۦK.�x�WA��+���9��=sx�R������Ɩ7��?�zj%E�ܪ:7Y�\���c��HSx�R����\��.�x�
�,!c��9��Wb�^���5���ɎP�\�0�]钚��L!O�	-ކ�i@�3���j��
,8K�
N���Ϛ&����晈m ��ݸT@3uh�����7������9���*BE##زˠ�Vp�8���_����2Y��L�	D�iԂ]�N7���ZF2�V�����@#�5[��](�qY��g�p]���k�v��c$��#|�#<�5k!��]�
T(���v�G~BT�y�M_@�I�!��I��v@E$�
��c�� Y81�S��C��L�˞��h��s�e$4�:f׍������է�.E�=ק�l�������qcJ�$��79#��K+�0]��F�,f{�~�{3p����;�q���Pn5�H1o$V!B���� ��M#Ӏ!��y3l������Z.p�	=��)���ӂ���PE;)e��3�f�3uw�ő�н1Xq�*�e�X��f�O0�]�Gִ#�x�6�v`��%����xlY3�,y�t��P; H��s