��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf��4Oᐢ��\����.��4M��A���8}��]�j�Z�I����7�KC�����#�~9���-+_�J��[�O����y�p����i�������+9"ƭ�ٲ5�����I�]|p�|�+o%z2�Dx!n"p:���T�O@�^���aoC��_7��ؙk�e��O<����T .eb��\F�C�R�_���ń�$�Ҵ);І=��8zPW���㮄�pm�P��eۻ5n��1���؊芖�u�6|��-A�� ,��픬E�C+/Վ�'�Nx���AON�V�!ڜ_��+�{��Z~@1��i��� X�a���g	D�?:�S����>�7�tvJ/� �HƮs�j+l�qi,K��ݢ;w���d��,y��0��	p��"UkZ?�ڎW�ąlAރ����J-�+���٨�<qC�����p-�o����k����p���?x��$�F��Y��<l9������J���E3MdI}	��M�,3��ZFi��JsDX���X�6q�������	�Ї�c
hs/�m�Br3}�o���3-.��_$�ܪC!fc�k��csL����y;Ag�A����1���8�O.6]��z郠ŏB�A�e�����tv����h�U9g�xJ�9��^�]1���Q��a�$b�kLā,��%����'�6'E�p����8�?Ƅ�ﰟ?�u�SV⋚Hɧ,�^�z�}|J�J�-�r�=�1��l)�f~3'tʫ�N]�13$�P���ΠxsC�e��F��!�^Oᒠ�$��q�a��oD�G�c�)j��o�5Ur���:l{|+b��T�{u�+�~H��2TU������B~esApa��;�g����v�2b�������u�@��JAu���G��|�m��t־+��%ʓ�����*sf�7a,�x��GS�9�����+�/��$���h�7�~$��Qx��a'3���H�.n��r��z����H����¡$��p�:1Μ�Ħ�>ۦ�XBye������0Z���)��tQ�=�����⡶��(V��8�6���uK�I3}9<�sN~�,F��Mc�C��.�ǿҽ%V#4ͪ�
]���_���W��̧�i��4]��u<T���;s=�蹽e��j'[���d���@�C��x�Z���o���\M�`Ȫg=��)N,!��w������9���<t��Ǘ��^����]{Qx�6/�H�g� O���8 f@�E�N۬�R�W�t��4 �q>�v��5,EIf7�)L�z���-��X!�p��H��s�Ȃ���ċ���0oSs���߬<($v�kU����˹�$�ʢJ�O8���R4|@��]�?�1i&}aZ��Xf���=�΢p��bEM[���h5s��ӌT�dV�o"��bB7q�4K��]��������=�v;�U���#�Zʱ	fBkA"�,)&��Y�'�/�B�6������.,��m&��Z��L#g�"�pe���U[D[F�a�
���\��c�$�z�Ͽx���f�D 
Ũ�^@�$�g�����g��c�k���/]A���� It$*��(i����ȣHY���[�Ӣ���6M�.O���
8��`������{�%_b��X�����tb��@A0���g�n^���x�����0�7
<�h��q� �X/q}�E��d���W�Nx�$���:
[d�3��@$CQO�\�Z��o4i���"���@|`�� 5!��'
���R�9`������)������Y��y��ʇ��C��QJc���)�w#̀���H$$_?zi�uQ��)�A����<��w���&��q�}�c����1��ڒ1TڻE`� �h2�=9z�upp�T�A�/��/�J�_W�R&�s�{�.�r��+x6Acp�'�RV�B��p�Āu��"�N|�h��P�*7ya�� l/]�n��rz�:�g�9�1�iй��Q�I��� p�,T�����?+��QI��2����w��ԋ��b�P�7[�Τ�q]6�p���8d&�2�� �s�	}�Z��7���'�T���Q��dh��jb�&��w8�gP҄�����tC�h�^\
&�{1s[;3ah���C�����Y�՚
k�&iE��8�V��gּ�;t����~��L��R�D~�j��X���&�4�!I����(&���I�0�ɶbe���x0�i&^a;$|RG[��W<���i_�7���r,���`�jE�3��:7�A��LؽE�K�\��o�j��(�b���`N��������/�U׽'TU��c�2�/���0��Xl��ieN��~U����sh����~��E�-��_�*�;`E�H`:�>7p����A�B �ʣtE��5/T�x�W��{�w8tώ4�~Ic4E��f}�^|7����lg����zdZ4F��2&r�d��<M^tOx�
����c�@����~������M>#�f���6Z�l`+@Dq>ATD��� ��Y��@���M��ϮP���L9�7��ȥ�Qۺ�z�d�R��.�j姙`_��ğx��'��5�y���^�ð���-��Z���Fo	�H$y�COŉX�d�ZL��e��"�^YL�^�>z}#ʣ���
m��e��6ᴒ�&�g��J�3V�&ج=�����C�b�C����!e0}K�g��e��E�b��$G�����F�J����T����C�z�}�I[�ܚ��l��*vRiM�b	Rl�h����$�̿Ņ�w3�)���q��F��8�kݦ0���@x�� "Gc��d}ac�/k	���9|Sw�*A�گ�]�C�i?|�p�#���I׏�ey�p8�M�m�~T��c�Бd7"�8���(pQ�Vp�d;� �Ͱѧ��(ǽT���[Y�)]��B������]�6
�2��؟t���u��*���j�s�4�Z[!V�q����;��s��X���=T��9�_^q&�T��vF=��_ أ^�D�7%�����D�/��^]��_��ja׺�K�OE�eE�hk�����<�E+�1	2����p�5��HVW X�Gf�4|+��dZ�/�I�Y^4��.^	��6�k_��PTMU�&mg�-O%���i�s�c�86��{��1���#p ������f8W9��j��I7���=m��R}��2o(r����n�u[&Soy�S�K	�\	hm&8"��Z)4>�G��Az	��yඒa�����F�]g�Aw������;�V���Rd'����YU�ZO��O~R��7�̎ɪx���$��1j�D���S#`w�(�ű�X���Tz����@�.�s�w��I�6)�b�@&���#��C��8�Rǟ�YL�Mʧ�]��*�yc.���<�cQ��O�p �G�5�]�v!u4PT��M܉�no�,M�o�L�!#�>��\�$%���ԕ�����d�搽�5�Mԍ�ls� �a��mV.����:K�ԹT�g7(�r�0)�\n��sE<���M�ןv��<���Q)I!���`F��#�z��׼t���#�O��1x�{T�l?,d��nS����쇮o-�/�9n�qL"=�i��G�g���iʋli��I�U�b���	��MPTպWH�;�;P=�8���;	p�y��mTE��,��]M��I�N���\�<�A���ʦ��M{�����߾<V�lԿNS8����v�&d���o�}�;�8�WYM\�Τ>A�A��-�8=D���G�@��K��?�����Z�56t65�9L�7t 0I{y�`nC� :�Y=\�|���9�H�:##os̕z���R&��7Q���<lR6����c� ������T���*��\��i�d=��j�"ą�K�`ebô�N�F�����w;�0CV����F�u��,�]���: lx
S>Ŭ�o/�5��'@�0����2}�BX�
��1>���-w5�̞Vl�K�V�o� ]�Dw�6A��/B�W��K������	,p���(^P&�1޵ `�n��&S��H��< y�^۱�S���c\[2�9P�Nw'����y�9_g�(r�p�}u��XG�B�w��B;���_oo�kv'�M�N�'kQ51ۉ�����NmGd�*I������Mj��n2_�'���򂿔;�1!�]�v��晀�A:җ�:�i����jnt���tݘ2gweʒ��GcH�1����llO�z�<�R@��He�J�c�L��S��<�1���~:�M����|��f�G.]����d���Y���<^9��'����|�\�c Ln��\ZY�y����#ӎ�1�tYkH�@ 9��NɌWt���E�#E�g�f/@����X�� �iN$7?���UZ�2U����,Ǉ���]����b��x����QB���$��>�.���޼3D$5[DO�xI����db��[;�Ҁ�͔l�� �pa��>s�%d���[V���� l
�W�[���sH��CG���I��^��¿��Y�{��Wֵ�ٛ��A��ێt�j;n�Y��O��c6*BWH��u���/�[��י�W���B�a��~=����,�Dk�u����W3X:uM����3󫬡�k:	e���ͷDq�w�m�ZIY�ĺ��E)V�^���~�)�2�����#��|�F��9ɊO�rY m5R'��.���$u��߿��߀ܲaR�\���0>��������riZ�J-"cp齀��xY v�2{-�mp�MfD�^$���8�Q�*Sx*0ey����B_Ed��Ѧ_)�.p���y���R�ϝH�����Gfl����	_|�oǴa×��չ��ŷA������<���B��\1�u�7��O�q��͠�b�c%D��x@�_qe�% 
��}<x]S3�=���E"�M��X�T(х}�O��$���ܗ�yr͋ף��Д��ձ��Z�0+f�KI@��,NlGY�u|5�c1Κ���@Q:Ao�b3m�2�,Qk��b<�j�g��S��C�
��
-&O�L�h�Z��_����	�}�v��h@	Mj��{�:� .����%F�!�G�u[��i͙KN��xLC�CǍ[C��cn�+e��%3��{��u�NP֧k���]ȿ5o��|��s1����k˫ϊ˅�"��e�}i q0&+y��0"��|u�-/��֌F�(C�#�?uΚDĸB�=!�^����H\i����¶j���l8��H`�c���fT�'��Jn�>(Y�;�g�~k�G�=���W���W�����yF�U.��YD����X����ZZ���Ɖ�F4c1��}�U~� ��GVJ=Q<��_:�DqTU��omEBX[Z�1��+��Srވ��Ӭu��U]�����Y�	H�{d�VC�r��3t�7L3�� O�V�9O���TU���a8���j�ƨ'�X�"9J�hU�}��q>�r�Ɂ�)Z0� } ����cԋ���D/�i��,&�ǌy�#��X�gڿ/��1D��S#3���ET*�.�r������+yd�5-GA ��Ë;<l���7��������׫���77���������P� c��"��L��(��A����L�?��(�٬Cx'��_ 7~̘�a���� V4G�9/�����K�_��	?^�߃��Gc�F!H
g��K�at�� ��Z�R�����L��*���i�$�lS^��7NJ�T@�OD���LW+"�C���0�"i�b,��^��������D5+|rV�DR[�x�6i��p7�ol"�-��9�����^��>����H�x޳;�D�A���Tq��f�G��6
GT2��O ��dDf�����[\v+����	
�Z#
t���y5n4z����>��ϻD�RȅT�\�:�z�X�(h��(��������:�ю�s� d�a����Pk����IASL���$_�����c�BX7��#���|��6D��r4�;�"u��-�h}�lʩ���Ǘ�������l|�w����X0ʄ� ���&.��%����6��>@M�0m�,T�;8�����ɩ�ZP�k���%恳{k"Z&N�y��(�qx��;^.�F��J�Rq�g.�C�B�z$�@���%w�֌!�h��Z��Bc�{�c��_׷ϏT��_��?J�,YJ�({��J�z#7�NC�AuV/��S��N�W=��h�vb�*�7?)��*������w���#��_�7#��9^����=�)H�3)�B����V �R�Ƙ�)$+یN�`1.pCG�Bq�J~~��"`�j:��VWt�������iFZ�[�����'��"�`�[v�F�'�7O�m���m�����Xx�pŌ;��3H$U�_\� {�G�uZܔXg�HU��j,n�E�=�|��a����b�=�<ͺ��V��E� J�*diy��� ͇�8ٔ���.�W�p<����� ��_�Ѐ�q��C�ɋV�"�8�}��vU���0�3�˦��Q$�ͨ��ʈC���*�ڹ����\�? (�iWŐF��3�	�qu@�����:��d#�c����~��}�B�"�t����ZN�yP�%����[I�8�i��YM�$6JD���W��-��a>T=��F��,k�����чuL:�l�	x��{�-���
Q�VA� /w�'�Yl��=7�:�K�����9��S� 'ܕ���v<�"��o�}C���W�$mDg�Q��X��U��q�ϑm���)���0�1��r.�X�q�U&U�]�W4=��J�8�G�*�������H�H&���F�O��^�V)�h�U��>
��d���T�G4xB%m:�)�&�&%9`����I���ڀ}�!�n�i�� �h捲2��o��Q.�@!��n&�'��[�{0T	V�]͵y��̃����ńl�ka�Ai,���|F𮒾��������T�^��vׄU:~��~n9�ǝ�An�pF�����"���pF+�u��ޟЈ鱨x5Z�U]q�M	���DtL?����7}&h"����w�H���H
5x��8���pS3(ex��iF�[<wx�BN��\��L�����27�h���}���o�5�⽳]w'ۣ_ﶥ����٤��1�9v���W��X�K��0KT�����|���0��O�߻r��-cGJ�������V}�ӂA��hp�X�i��B�Wt��0�e�迸ccu+�������	Fg�Y���;�x��a.2,��I�?���-X�z\L�ͭM��~:,�x)�O i��p�\-�����|���e^���H�h��W���>�ꛤܤ��BCE��<�Z���+�W皰J���h� �Q��+�Д}�ԅ��F�OP(�z<$O����}�J-�!6-d(�,B����#�����#rG�>�+|�~��&��۵����8��򁻀�1-N~VƯG����{txM�����z�X��!<r���.�0o��ƗT�QhT�ϟ}�PHb�;:O��{�cw�� �����Jx��ڶr��&tZ��4کc3�>y��R����O�����곮����P��i$�ћ�-k��E�a�Ȃ��|D�U�?4F�̞C��r�bG�����R���&����Y8<E��	�\�X����O8T2}��-��y�u�^	s�R�o����/90W�� ���qx��*���u�r�]��x"�{P�BM$a�x�n����D�g�N"`w�⢎��l'	�]=j���$Szq�5�po�Mn���d�q|9R��êܱ��p�;8��V`�+�t�m�-ݪ�~	�tz4tn�	`N#\։R�l��/cj>e`�֨�H�g� �^������V�R�ğ�}[J��wa��p�621�?����V;q��<�듌����)�Z[= ���bz��"DD�o��R�V�4T����u8�<�?�:ǝ㞇W�����%K���ٜ��ԛM�T �����U~��m����-vb��~�,G�V�~���Xp�c�ۣ��u����Ӑ���j������EA�]�b����	�$�Y�� +g�8��ya[��V��%&r�D'�a������1rx���.\T}����:�|�����%	k��^P!�y�T5�+
O��'$�V���!3�&9�s��.pe/rjC$]�����BU�#�<%��w=��&�6��T��:6b��v��z��iA9�^��~n2�Qdq���H���,z��p!�9��/�ά"�*H�{������#�&�|�Ja&WM�Q�#�ms7����r�/*<��lS�q������"��9}SF��su�P�ѫ�eu��K�����59�Z`�R-?S��9���T��&$a	�����}���=<���(B�c�o��k#�I�Oqr���s�̐ms+S��v�ʝn*G���P+�y$?��2�L-.Xlr`Ka��L�����f�H�G2Ly6`j����F�r��wwf�h}�<�,}�oA�r�7��b�U(�ߗ�Zή��"���˽�L��Nj�2�V��'�[�Y.#B�!��k���g�%{9�m�L���Tk��J0�HN�uZS�,�}��~�-�Y-�:�=FBЍo��3�⁞Az3呌�X1��ZS��V�}�Zi=r����#�}-�M�J��Gj���k���Q��>��>�]�I	qsPt��;��Y�*��J!nZ4�� L�C�� m�vҲ>���s�138��E���N�:������MOu\���{�_#DW��;G�9����S� ��������D�j<Ut? ��Tmx��w�U)RN2�s%��G&�H�ks�3�|�u��� |��K>��e�W�K��.�`�ns	Υ>�,��M>�<��A�;@�tٍ³�8Y�7���4�*c|�r�#1C�@mDs<�Oc��{��J��
�/��Q�4��,tЅ$�|��a�a"���a���$2#f�eѢp(������[�B�`���L~XV��;�F�ve��Ƽ�8|/ND"�7z���x��zOQP�&YH���l�W�ϊe�˃��y�\Dvl�;�Vd��/��3��d�!�������۸]T>e��ڒ�F"b�ց��w���@�<6��o*��Flo9�I���=Pe���nc��]���B�wL͞�G�B�tU^�����y�*q�fQ�d%�W`�����FG�@����u+m3�|���oh����D]����}ܣ�����Ə����CZ�$c�ݼ{�PuǨW�U�����b���3Ⱦ���i{���u�	)�	�W��Ւ;!����rP$�q3@��lI�Hb*e�%��'=�z�`�fOLo�aϘ�!�6Ԋ�~N�:������k��yo-��}���e�����8g���=���U�'�U������O�[ �w�.e�4��\��)����C<�����I���� GL�����P�1��F���dqZ�\����Y��o<+�t��#���{�9ezO��`�t\#Ő�%%li�x�<��ۨe�%�Xp�=���a�t���l�g�*�2�6��=��1o."��֮�(	D����G���DX:��x�oyׂ`��#�|�a*���ʮ����m���ӦV.Յ,T��������e�\��]�4eӭ�`s��,`I��I������D�h�W���h��(��W0s���}'ewW+����tG���t:���V|�u��W��|������U���/�=s���?b[�)����ڢ�H���̥��W61SX壙��(��O[�e�"�^D{َ�6cƎ
�hp���0[񲿯�)�h���UE����s���pĹ������]|�D9s�$x�pfR*c+QF�e�C&�ƿ���X&I�� ��Y7v�A�ݼ�~K�)c����%��\����7�G���M��ը�I���Ӡx8��6�h�Cpy�L^��#]����s�l�qd�i �:U^V9c�,@��Ԥ 2aD
�a4%�S/)3ı'힃��w�V��~�\������?�qq qv���Ir5�����)^,̐u���};�e�үHf�c7��m��CW�KC��UR{����
�r�����l"�?	�_��9w;�TF�/�R#���[ܾ�?J��P�8���(�ͧ�$Pe�t� �q6�L+����w9�zKcB�����>�A?�jH��0b~ x����i�a������!���I���R���:Ųlc�}As����8�1Pݏ�ۏ��X6*Kj&l��&��p�y)P=3�����_+��]���E+g�gxt��.�:�����l�D'N1�JaƁ��"nH��VF&��0���>ok�@r����v�r��)*�`�-7�����+E�M�3_��׌\XF{4L0G���p�.�Η�bqb�etP�����sWMZ� �b9~��
���Sގ��h]�n����E<�f/�g��)!)BWz�����i-�N�$U����q�0l�?+����1V�M5��G���yy�D��[��\k�^u���%ʎvc��c#U�A��m���a��u�k	ov����ř�P�=�4>�_Zfh���Go��Ud^i���m�7���G�w���6����).���F":�BfeC�8�r�wJ6	�t&���J�5��
�c*��aF$������=��S~DbW�X��x7vj�_u��H�Z���Yb<�U�]u7�ˍϸ��Z���2QA�����O���~�	<��Y�+?�j�2�����.�����m����妩L�L�9L�=�]�E�R���s�D���d߫�K۸â��т|�]lO7egm�P'7�z\g&���+4���gqm�%��U��)����O��ӢW��Zt��+��7�{ v��r(`X�lb��W�BJP�j����i����01Zۯcs�+S�i�欿��� &k9?�/r2��v���Qb䮱=������v��Vki$�Si����̡���^�`�!#��|I�?Iw�C_C�^���uUF�C/Ig������o����a��)��y8��烞�^��9/�it�m��\��
�4!�v����N�9T�~���E��U�_����v��&r�(�\�o6��ni%7��J�����Z��B����Q=0k��$@��n����ƾy���7P.BWޱ�:C�5�)(���:Ž?����PR]G���U��F��f���Z76����I~��I�9j6s�Ǘ!�xwS�"�J{������`A��F�d�]?�����Z��[�"���tUى�G���v0'�<�1<	���鷇Q�0��ߩ�������}c�]�;`C�&�"R�m��R	�5����2~�������[C���U:9Kp숈��;�������W�a���Q�=�$7|9�$s���݃��J�,+�J8 �秧�ո�[����?g9�>Nl�Z�v������?�E9{��υ��Q,���Dey_|h�-�e�)�Hb��5�f	��'��X�'1����EN��Nf�2����d���5~�d���#�&Sm�l(�~���Ж��&�j��Wh8�wK�̋Ͼ/�Q��=u)R3�po����_AG�ڬ����fPQ�!uO%z�ѵ�Y��JЦ��X�f큕�Q$��Hܦ�!S�c.3}�Y�v�ߍ��]8E^zF,KmI�����x;O��a"���Q��
�����`�E��&�m1|ku�z�4l���x̷�8�4`�<<����mMg$_��6���f�(�G��\�o��b]O���C^18�R݆s��e�� =2�.[�[-�!*銦�����K�q�wJԹ� r8v�zU�Ck��z 0o�W������;�+]RčE�+��#G:.�X3*G���݆�tx�3�,�FW��+O{�.oP[C�:�ĺ�nCH��k���x%5�+�0��K���M�`��`�zJ�0��4� /
F?�m����f��"=ry܏��ֺ[:�ǽ��u��掗�DA�+ZT}��cA���?�����{	NK��Fn�kX	Z�F�V��`.�j*�
$9d{�I�1��*	�8ϾC�~��� �usC͔ґ�VZvb�Œ�7.�w����c/,��ȫ�-��/])@P�T�����O�$��{���=��/����Ԑ�/��G��o(�`�2\n�M��C �k"�<��A�d�� ���j"�A�3��p�0�(�<hY$����쬣��%3�-���s�9�o^�؃�<�N��H�oJ��-g���dY�Hvy3�A���R;@s6�f\�>{�T����*��	~�0z�T�>�ǹt�R]�iw[��v���eS\��a�Ǹ�ծ{���rs�Y�w���Wa����tC��9-7THWL6n�ٖ~��~�F�I?$V���i?v�/���c*������](����uRE�)�zlH#F���>��nX<�Ϥۦ�w1�T���]LE��7"��s��t2h�ŗ�AY�%�2ڦ�+-��[���D!�g���ޚ=���.��������~4��4�Ʋ�e� ��{���9^���'��u�jc��(�,� g��z���o�=�yƅK�Ԇ~�p���
��������\���ğonha�`
v�`i23��5(\���Vqo<ńT3��`�VI�5����kWU�C�7�����`����ˇhp�f;:��O���ܳ��7M.j�M�㫏���T�J�*I������y*��rYl��d^%��1�_�j��aO��)�cڛY�/��H'��er��A�L�,�t���['�>��^ĞC|�DE����A�: *ۗz�HU��j��7v�Cka����@�JA��pOv��Q��D��(z�� ��RH�4��Av�D�ۊ\��2��{� 7���@�-�#��aZ�e�Fo0ق��8
3��-�����X���2��+>��.A�n�U����ow�����*yܨ��3S['�#Z���3*(�V�����u�E���v^�S�߽,'����L�`=�g��{6����$DRG�g�`X"�Qq+R�i;�Jۧ�'�Ib�"mg �%U��tj/o������b���<8gZ����̑h�}�`� ~V� "h364E?�5�l��xM���v!+���R�G�����Xrh�sw���i�&iYJ�$.��џ��+_(��hy�Rlr������mK����`�D��s����WN=�)Uϒ��!<�hy�\6��g���A0����������*�j������� �Dq6^���HC�b?�Գ�m���1��ƨ���ET�����
�s'�aZ���mH��2Y�qaT��D�I)b�yC1�8�x�x���U�a� Tg0kT�_�3[(3'�����3q�3��?�B>�����L b�fe�*鵗Tk5�){�dɤ�$�8�(�9:n�i�J5-A1q����f�82���)��n�-�1�{��^��4���e@�l��S^����I�O�<Gt����m��?v�#�׿F-A� 5��c�b�wc@�x�=P�xe��HnZn�C���T�n�ꦼv�so�$�����L��/��ºӫc��G,zqRY�q�銲 ��X���|F"<��8�5O�~��U���d�� '��fY0���[&���Ϸ���I�T�������Shun+��q���3½�<��q-ǰ�����o_��@,ܼڱ�o���z:�t)s���D.���}co�mc0�6�y���qqgN�nz��K����u%+|5��ɐ���R��?���dE�a5�<A�P�i�b���x����!�M=���5��Y���gGaJA����^D����3]!h,�O�dxֶg�H��<$���5n�%��=�
*B����i�͝�v���r�t7��i_?QjUpB�I�d?�B���fʲ����lV5_�gW�gˊ�����F��ރ���K��"te�lp)��=�hƯ���qa�O�w�M���ؤ
,jg:=�+�G��٠���wdC!&~Z��Ϸݦ�.��{O��0�{�5�?f��@�.�-<�	nbQ�_'�!7S1����p�p�ǼCXދ��3P������cE����5$T�`��A	���TZ�#�*�0_@È�2XS��Й0	*�V8�:[6Z�>����[�Yo[yc�:v�Ǎ���݇'��o���`7of�̗��n�uS���`&��H��|�V���F��g�x)��2@��`�%ȭy���i��}gv��_c�ՠ�f>��|�E��¬ ������,PM,�3��1x+뉜���0�i��Ά���H�&�@k�9@r�׾HyO�b�W�R��)�3��
D^:�BFj�w3{ٿ��Ye���9Y���_���=���Yܷ`�YRG9F��'�R�6�rܐ@9�Y�'̕��V��V[��ʹ;~�Kg�n<�@(�Lr��I��6�1i4Hb�z=�$ph�?aIDf�;.�P�Ä�YmM��1R"�s"Hvʬ�?|���<�Ñ�{?�<�ڷ]�y�V�3w���UY�8�蓛��6%��RG���I(o���Mo¦��(^���VN�|���I��t}��_1�oC���E��zS�&�7FR�0��ؒ�b]��ܲC��H�]����L� w_3Ω.�
Gpߠ,,�j\Eb/r7�{v0�?D���՟��D ʎ���%�aj�z8ĦX��_M}�?A,�����%L�6�Pc>�'��C��$0V�s��Y����1h7��c��va�˨cН\X�G�4T�@�Y��}��
4z�l�<9$��� I����tn3�U���KТ�(;�$��x�0r�T�����q�< �[�7��qM��˾��������7���?�;�Sc�V��TU8��������U�� (�A�W��K�:����'bt�7���P[u�|K���5��\�g;ҋ��������ⷈ3}�o	�%5x�e1�!(G5ح��7xŬ�A�t�f��^r�dBӥ����m2q{��<��i��B�$vWY�#TY������'���#�Y��T��^���F�'�X6��}�B�s X�d�[�b��0�d�7d�;���-W%A1c*�j��2��RI���˙̋��9A�_:�Q�ܡз�Ee�{G�������(������a���Hon�(��x�PIWS$���C%��c\r�qъ���A!�W�U�B�n["3m��[�XtT{t�'fD/E��@0���rͣ�[*fw�	�A1}�5b.������l��� �����DU�k&/��q���r�f~1�09��pj�V��_����o-�Յ����e9�F��2b�mD��:����ŭS"����s��^r��(��:�WQ��UP�3Lh˿�M謾ڑ �W���5�|x���h�@b���U�ր4>�Az�d#r��jyچb�rz05L�
 u�U3j��	Z�R,Y���� Bjh1Oc��4z���)����h`r�M�����jȡ�lT	3aq�rM�y��c5���$�1��S�߾޽<��h����z0����U�c|��n���\]q|�O[4 2����zs�@p"�����4���.�B�tJ���"��E��ծ2��]���ll��k��w<�e�{o�:��]���qܝe��K\�W�S�$�,J�,Z�q�C^X,���h�$�{"<9����w��!����4n	~j��1>��>'Ts�w��չ��� W?��?Qңe�f�ڠ���y$�ų��L� ��A�򨶖!8�Yq;X�{����1,I��w��5ZڎǠz�܃Y�וI�S_Jw����-V��(vˌ5��+�ac���`y#I�U�s�f�E]SZ�����m�����H*�׳&�y�������T�C�kج͌V�����PzV|n��0�����d����%԰�:E�_�$�ԛ�����m�LN���Q�G^��sd	���t�zj�3pk����Ed�V�b����|<��< �M�`G��j`[9>���_�
�3|�ov��z�d���34�t6��=9�;@�p�bL ��Vh��������n��Y��ۿ�-��po���5-���i#Ī=�O�GT'�K�R�P��ᵧgtp���X�gf�?A鏺�:�b0zA�G.O���5�S%̋f�wp�B2GF*3�h3����������9��
#���/q؉�:��%��X��<�����KK��Q�Fiy�V���;[��N��&�� ��_Ͽ���v�y0(BBʙ�1�?4e_�0H=��1�����q�ka�|��l
��1�w������xSC�.���j�<ƕ¡|Oa�bo�r�j`\*�G������49����ho%jȯ��*Z���������(���禍�[����(���;���)�d��o����\�/fCi+�;FCi�4O�>���p����tE~�_2�B�אp�������4��HX������.�
YPH@�u��XE�oL[s�W�h���}���y>�敵�=������.E�\h�T��ݶm:�H�?@���,i����c�>��ڦOV9- M���0P��7w�oeb��,l���r�猿�����)8Z��ވ�q�������������������~2Q�3���-���s;2����d����2g,��<C��Z��'������i��A��r)� ��Jx*�T	��,���Ȗ�8�L��_ �mK�P�G7���ٗ�>IOM����}�;�Е��@���0I.	�����Y��3�+U�e��$=h�_���~���Cr*X5�P�k���%
��$	���c�JZ�X=�e�5���}$��f�[�e[��]e���4�ϥ<�Z���&��2��� +�d�lc'ߜ�g;�[�x\%�뫥�߀=�8r�%��y��~9��� ����� L(*y,9 �g�G��M���^�d�\���5 ʢ@�$���HQv��)$�0��7�g���1��v!g�\բ�r5d��LKuʡg�݅ꟼ���|�@�3^3������G
��O`/�u�r���g�n�;��z�j��,
�� Z��?��`�t�y�O�ŠO|cf��\�g