��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_����m�e"kxu�Uٲ"#oB2�-g�j��h�p� M T�(�P�+M��&�[���+ǚ��.n{Q�̅Z����&�;3j6dED=�Cl���ȸ����8�^+����K�\u��8���f�u�$$��LF���ꆶ��xV���*'7}�� <���.rQ	�+ed\���M�����$0	���|�v4�6X�Ṯ��݉�g���ܡ�j|87���}	fܧ8ƐUԣW��JB~���s����ia�5I�� ?xuV�D��rl�/����!���\u7�e����@¤� j�8� J�
��<��i�}�����L�g��c�!��7`4S#�1��pϏ��j|t�i�\��\��"�4/��)1_�=�Ul��n>��`���ge�|RX�3d�X�7)���z��j[/����b��?Xd.oL{��LI�d>��nٸ��4�d�Ƹ�x�d��="PG��
����� Eƙ���F�����z�2s�a?t�Z�k�������%����?@4���y���%�:�:Ԡ�Z"�%��h�7 �Qi�Ӧ�S2�'�ԥ�x��S�㉰KO
L����>���y�����H*��7h�~�6�Y����C���*♻=
�A�`:i�s��_g�����f@���}��ݧ u1���+z:<Sk=@͎a��p_,����&�y��^4�����[��m�
=�~��y���<�R��9���f��Ǥ��v<��K�)@#g1ow�mX~�=��PH��=�Lь�a�!�^�Gl����6S9z�o5
�F�~&�1`�����I�\k��i�7H�KD�(���K_�������v��PG�$G<��t��������4*���i����!�a�A��H72���w$o�Ig`�g�����g��j������pi��M~A�u5*�Yt
���ၪ��<Ǫ�$f3��i��U�pM�����	T�_b���1;��@L��JfI����rT��h���i�g�yAL��y�?��,�O謊�k��6����#�^�8n�;�[f��1#�3�̒,a&ĀOt��~}4���k�{�!�xx���ݣ������7�����ĸ�����?Qh��m��L���c>"�*�;Y�����m��.mV���6Te/�j��:����p�۩��{hY�i��N�?y�K�P9��x+G�T<"i�it��	��*��?�S���}���b��<��IO�О��P�#ʃNem4/G�R�|�����$���}G93�����9���3�&�p�rd���}Z����8(��D|kv_D��$R�մ/8���FN��+�֧2s$�i��Y>hB}W[��'I��jԂ鼦0d;��\��.�?��oGy�R*�Eu��Z�� /��d6����2Л�@�eN8&�v��J�]��Bj�������l�:�./,��T֚đ�}���B�����+zդ��H�[7}z�]�Z7��ߏ��"#/���}��<�����̙N�D�h��(e��eˎ�Wr>"nh�jM�'kl �Z��gwü�!���Y4���I|�~�mpG�b�_���#�S	&#��i�R����N(��:�N���b�~N)���6�����+Ջ������}�������m�h�wTl��W�z�<�%;h4����H\����f���2-������I����a�6�m�NN%�ϣR����I��>8����|�M��1!�w�h����}�1e �$�mu�!Ab��s�!q��
�t�M�R���(����ӗ	��
�Kd��!��|s7���>����pZ���z� �+!M��g�t)�҄4t���3['}z���=a�,Ǖ'N���.�	}ںR\{���K��j�޽�Q"�$Y{}5�ѓ+D�
/�<�Ь�G���q��R��o���� ��/�[;:����"��j�"[��c��31��_>w��4E��&�o���(Y��j%@Ֆϙ.>ߨ
	X�#��Pګ
�vߩpӐ"dp�C^"��6�� Ug}wZ,/���$1��(�Ќ����S��U��w����aC�G`�R���y�-��sE��Ky:�⨉;U.�#����<�	�U$���x���|��y���dk��x����),8?Ь�y'ʁ��Pk���-�+L���Zc�~>oԿ��Up
��xv\'��Brێd��