��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8SjfSު�U��w�|����H���4�&Si�C��-��T�L?yE��ֲ�l��z/�u����)�?�C:2��iK�QF�nj?�y��t�q����<+4̄D����;�0���������)�.M�pd��`)��,j[�����(/Ȯx��f�(M=��g�6�jTE��kyJ�ow�m�p��M�������'�C7[
��mB�G�oEh��FM���ԀM��9����0��,��y3�W�U�;A�8��T�#`W�v�'�H)hϩÔ{��R�2s�7Z
�a�gv���;)8[���+�9�gR^
�B���<n����Ta��_�AF��s ���8R�����$�Gȗ�N�k���ν���,z�R?�K�ҏ?�C�2�Y,g/fvZ^I	���|�0�C}Ya����9�J�8"B�u�L�֌qW�Pn!W��w^�2���)�UO�TAkln���_KnW�����H����=�Թ�|m`vM�\�Tݪ�@��GT�MX	'@LpE�<��t���cKy�+
���B�>D��-b��H+YFuo��<}����J�[�{��L�貣��ri12D��< �k%����m�;�,�	�"�+X>x�W>�Wۧ�Zѵ%�F���h݌�>�n�xSu�㬞�sc3��d���U�T ���P�,H��ԫ� Zb2DkW���ؔc0O5��`~����}|[xqwOXH:�"�:m�r��7�dY���m�H߿�:�ܿE��(�+8
�,%㖝�p8���F�@r/����J|�۹F�D���l���*B�;g/���2����w�b��P2L|X��^����k����-.�Tb�{gE�����i̋�᜴��J��שd�OA�c�0[�&���%r��B����/�ҥ�g�9'��nG�Y3����2���j��覵BD��d���Y��\s'�f�ռܔ.*ݦp�i1*�o%�|����X���e�/eB+�J�G!A����[kh->��n3aZ��J0��cQ����uN~�����!���~��D������	��G]��?�3�����&:�;��g���h<%9���jT������[О)rA|�eCķ��/3.@3ԡ�z�UJ�,]�����Z}����%���|H=e�0�Im��>{q��p&��������`�(����Nj�8��oY̌��	�^kmW�쇒����Z��)��n��L��teX,���A#`r|Ջ�Ȉ.�W���B~1�A�v0Es�Pָ�z��k?�5#�}^�ߑ���SÁP�}�^Y�E*��*���q�.�}��y	#iF��ٲ��6-ܟ�D��e�h��3?�]o���G.a|(��|B۴����'���$J�Y�8��6��&�����:��N"+����Z
�tSܹ(`�~�ٌ�b'
�k[��`*~���t�~#/ᶒ����4�۱��+�G�cU}���Ŷ(6������![h�U�k����K�d���Q���q_^�@mhC�Y��3rn���/�b��V�-fAҌxT�֣i�M�V_���l�S`�M�[4K�Me�!/�ɵ�^u��n��=�l��_V�@���F���yRK>�`���������4���I4��0�أW�N���͛}QQ{$��I�3
�e�>W�b�R?i�����(êc�z�T�p����್�һS�&ˊX_ûI�W�@~�6�;���tH
9��¡�<7 Y�3&\���{ɵG@E�7�[����*M�mf������2"l�i-:�'��i�8Q'pd��>�����p����1bE���tAQZ����^��$7	��\5�g�cG�<[k]B�R���<O���ǥ	r.K��Cf��0��7{��H�`���9 ���%�1�Xm���n���X� �e�_��H�>�Xm���ё�~؀�n'��Q��q��bu_Mo?�E]4Ji��u�(|�{ ��G}+��ؽv!#}h��RV �pL5�OR�jnS-`�<\�/D4Nϭ��L�!J�Y�|%x����ʝ9��_��4)8uڟ{$�[}��&`�Dʢ]�N��隄 �Mu�l#�����۶LC��Wq���ߠ���� ͩ�̮�q \�0��j��&:+��H#�xZ��$����OI�8]-���߾�y�Pơ3���{�""�:��
��L�0+%�p�K)�>T���#-X~Y��� T�{K�Q��+j��o(�|��%�Q���L7��ȕin�%n~=�Y<%X?���<D��f��q
a�������)�9�R�Gi
<�ɲ�U�XQ��fa��8���C����s�oUM�[.n��X�r9�Uq�h�Y4\��-u+%T9 GOB����n��d����o���8��#?}�yn�/�ՄD1�.:#� o�f�Uݔ��A�	�I�E�T���'��S�V��k����r���B�!V&n�}q�s�S�����1j�}�����[fKT�<5%����CR��r�Ѓ�h�	�V�xk���0��aǵ�H,�����#��Nܞ�vDE�ֺ�������@1�&�*X7����?l�G"ۺu-IL����������Z�5�u�r��U^'�I&���u���s�r�+/��8�.sN���^�1Pv��EE�-"#����}����A��W�^��fr3z����Eɰpp��)��Z�k��/K�#�#�$�L�_�DVl�O-񛜓{������{�m�F�2?wd��Y��6�z�� ޴����tڃ�>�sXj�s����5;�F$7N˳��9�;R�s��G����=�/�2"��!O\*�'鲲Yn�pRy��_�Z�i1��yY~yC"��<V��m�
����:��b���dJ�'c�m<��mˉ˃oY�8��%ݝ����MdҰ�K��e\�Y����Α*�yl��Nο�}l�:{�؃�L���-Ԃج�	x���ϭyö]�br����y�to�ɛ�E��5��1>�g��㘠�J{(Vq��(�D!����Ua�w��V��������0ھ����b���̋MN�"Y�tM�{c��gXh�����̭�	55�7�+7Ĩ��36&�����w$N�+��	&ƫ'2�$��b+P�M.9�R\3qo��
'*�&���J���g�:U9#�hׯ�Z�����y�X��_�k��YNXKee�EE ��;LP���%.t�iQIȀzoDm�8;Z������v�N�)��f."�L~y��
z��e�,�?�8�b>K6�I��ޞMӬ��X+��׾n�Žy_Y��4�(�H�W�I;����^�@��\�@�Q��Wr��⯅W򝡬T�q�/V�.Z=����<�յO������ ��5ub[2n�|��\u������ސ����t�b
-��
�X�/lI��o�s(��d��y�=�=�w�pB�D6Z�k�]`���8R�Ï��Lt3u�;�I"������h�{�p&�K�M��|�x�'�Q�0�b��v$i�I�<��5�7`؇����p-^v�8d����"
�����,e�i�����а���|�,��Y���!���2���o���D�-D�z����1� 7�u*y9�G�"m*ȫ�Ivʷ�Ǧ�^D�d��?��C�&�}�-	� �Rfp��l��wߐb�Cr��D�G���}u���P:.���'1��2���$Kz��i��e����'�]$T�&��`H�kaRS�g��T)W�
������d��MR��7��H-��l6Z+�2O�TP(HDFM)��G앗��- ��6��������{�P�	��F�`1L�l�x�l�;�b����c�5j���G�? �G0@.��#�����N&^qV/ɥ�<�'1�3F��Y�\a��/��T�n���{��-#@�h�_�����䑗,��Գ�k�O%]��0l(��A�-oI3���(]X6�-ZW����H�T��|����{��!F̽.)B30'{�S�u���;�=�}�KM��@D ���-��w��[�K+gV,�I�R1R��ý$U�� f�Ȕf���}�A�dԛ\6��&��m#�y���a����8g�Q�����Y��|���ɝ�6��v�%nڜ:�[�\$I+E����kX�a]�	o9�J������%��l)��f\��H͢�� )�t�H툒U��?� K�p=Ox��,�J}T�(�&*s�[�)732�����C�J1}RH�t8���r�`�$�+{���X�Q#d��<����_[�ȹ�dxNd�"���4U14a�T��(Wg��hK�̶���2�E~������}�k�ٌ�hr5��72� �r������"l,ne�(��J���Rp�
}��P`;�p#��$v٘_��{��Yƈ[0�H`a"b	
���V��/DL��;�����a��Bd� v�xn&2N �":��5���֜��(
W��δ��#29ʴђB�c�a�� ���+o�]:�V�l3���"n+�V��V&�M���R��"saG��Ң"ƈ!�T(�'�{����!f��;�e�J�. uF�B��*L���b33�,[���J��
���&dcYi@|A����i���N�D�6V��7�7�M`E&?z�+��6e�/�y�
.>�ٸ��:�-;�nze��e���89*�����+N`B#��!s���&�/�������~����^���A��#+�����e���zjqX�B6��ؗ�w7��$g�#tD#�+�ܺ��@r#΃�7���H��c����� �í[o,� �Y"��/k��<��N�(�o�����H�6�����F����9���P|�����+C��Hဋ�^s��Ӷ�搣���b����� ����.������E%n�*�m�F��Uy�OwJ��; �fU����NSɪO�
~o߁ c��m�+��EM7�Ŗ	�g�7p���]�L�u���n�d�;|�j����]�f�s?�q|���(�A:۰TI�N�h�K�O{]]e	3����)��V�}"G�����Y��h@�M��Yg�K�M�?\�u��
%ac#���Q��W&Ǳg��`�<�>��;�V��6W�hB�3m���`~t�ќ]�S�B����WT�#uCIñ����:��"i~��L�`v`����KLh�= ��Gf��� ���#H{�ʼ<�[�u�+S�`U�X����)�ۜ:<E ��Yԥ�n�������;���f�}5,ŸsD��v�P[ ��uM��fV7���{!��b�fo�����f`��(�.�ZB1n����?J�Lǟ�p�D,���n�:ʙsg�jB������P��E����`V���뒫#O����.����F׍��5&UN��N9�ܓ�;����}���u�r'�{����������-S�s�7���2J}���3�B��D���Oi�����m*��m��Kt�I�u��h0w{�:�eb���j�:|\tDeB��w�^X�W�=��U8�)�rSC�#�PL��=��@u�W��T�M�ݿ`5.�z�f;
��n��4u�<j�U�?�i{Po%��O�_�!'�����y����w��H�m
:IU��2h���W��j�RB5G!��'�եL���ô�zz��ꡁ�r������61�36+Gi����@����?B<��`�@��� O,�"$,>-h�|�M������.�S}��L�'�$�	*�-I�>�~��R�x��tn�Ոr���&�/M�q`�E�]g�6�Ͱa"�P��t]�z;|f�i�F�� %s��L���Q#����r9��Ėೡ��ڟ�Bhe��H~��;�"�G����b�Q��p)�&�ZO�b�uq��ӆ�l�рU�H�c���"f�=��ۍ��~�ꌤ�4 �''��6NkY��¨�Ć͉�z��?��!r��󊰬��0�ܼ۾�X����^Avר21㋠�����t;�:�#�ٕ�vF���8h��he[T��g�e�X�)򬬂�����T�3�@��9
��Mrl��B#u���u|V��m�`�|�|=�����
ݪ���AA����ԕ���U�LH���8~�"�����V�o1���2�&/�
v-�7ۓ�3��gVc�CqO��]G�����@��j9�V���z6��^�G[c����
�`�-U�h��g�5�9ԅ-B�OMΙI9�ID����G�>AL����@:.�����խp��5~�p3�:��5�i3g��/Ũq�C�yGd��b�B@�kԽ�>]�WP^d3�p"2^iS���;zRV#�N�I��ER�e��H�����T975�+�"���m���)S!��G}g�͝��ϛ�U���@� f��-7�uѿ"��!o@ �#��!�z�����j��y5�]���!� .�±aD+@b<��M�W���˶y�}��
�f��>�u�/슠��
�uŷ qփ\!�/QXsVMEC��/y���=���/[�������-i�����M�1XBZ6�|�-��l��7	c�2"]�H�$r�	�dx�A�-��<����$/��Ayt!8�RNe��;'�ů�IN�� ��A�����Ȏ�C�]߱��Uz2���u	�����M�r�M��G�((2��/H?i�)]�@&]8�&X�:����h�p�d��P�I�8�`�ƤT��zEuoS��7^��y	H��4kE�TtV��x�!h��z'Gb�h�R�##�S��+��&ҟ����\�~M�%ug��\_��3�Tv��-�d�-P����A�7H�� F�x�ǹv�.?�%�(�8��d��:�#��1�1��q?�h8r���d>��n5��L��J�r�j�i��Kް:}�:��W�Ft��D�gb��̝ݴ�I���?�É0�[��	�
S��\R�|]�ag�;
i/8�M?���T]v140l�}�C�֍ ��BI 1_���V�.!�9�^�h���n�tO���!����3��Ֆ�}fw�F@���l��'�����i'�茗@J�Q�J(bE&/� )+ab4�R�x�K^.k�=�0(׺��HY��
P���M�\tg��ܙ{�X�M�:��?V �+*����*&"u��ϸ��&����ujM�b�D�Y��.Q�V��M��J�_@�c9��JM���;�z��s�=�^Y�zX۰Q����P��'`�e`����S��rc����6x+�vM���J��b{�d�� �&Z�q�m�i���ϲ��i)r쌂��y~��4�cׇ�8�����=�cjbR�|E.,\N�����+L���c�2��]Z=ϔ�[ӼX�5�>f�+�0ߕeCJ�ع����#�tl՘�O�>YP!�䅼��m1|;9�d^3A�AMUtXf�bEԜCѿll8��d�&b+�?��Ÿ|��#xn6���zm$��H�g��/G�(J�V��Ǚ�~*2�J�W'g3�%I�^Q�}|��'��jJ�s�F�1�Jb{`;@Vm!+�N�pse~L�����I�Jg�\q-��B����:��͙�<�*�Z��_
�aD�,k1sֺ��q��w}(���UUY�wLw�0�A�����Nx��K�>91�z�0ñ�����&ݾ܂���n��6!z��O�k.��d(X�8.���>��r�V-���"���� �8���s�[����y��s�����.$��93_qU
�b�,<�������]\/N�Jk�4 [5ۯ2�T��}��ؾJ�H+[R�U�n��Iwr;�z�B|�VyIӳLi)�����ܶ{֌C�&ڎRA5<@��-��8�E�5�����7Q�`���Q�����������8��zM)��֚�P�1D�PcR��!^�b*��}]7�o"rVW|:h�o�9���cɌ[W�4U��aeA�3}r�r��moN y��ݱ9����Q���w�ju�k0�m���S�dvCĚ&�LGBff�#Uɦ"��;��C{�'���׽W����ƚN~��ٳ��B����J���z%9���L5Y�ch~7����U��z!&�U����I�~0��Lw|�G�9�X���L#~S*;J����5@/�㑙�4'Ơ��	��g�  RN���v�3-ў�u��;���sKnm�Cr�t!&o�X;�a�i�zV��q(f��I`���
R|��I�7d�qG&yw�[���mUg��x�T�����YS'5[��
�Eu@��Ѐ=}��������T�_}^0�`׼��6n�p}*T�h�N���+F	�f�T1	�)���d��E�j׍l�-��P�����m5!����.[ �Vu���k�c˹�9��S���TM~Ų�œ�݃ѩ ��+���蜔5G����(��!x�������DL�<�>UL!k7W��D���~���ֳP�l��4�% g�n܌}�����BhÊY���'�[�Q���+��]�G��3̑ޤ:����RN�UCBYɇ�y1�Î�rr��Y!]򑙌Q|TɅ$�'��p��'A������ih�����u� �*	^����w�}t0����eא���+{|���C�s�ȵ�ϪT���bh���,���E�8c����o!�l�|5h�<��M�Wk��K�������ߴ$���0��%f^����5��H��Lj��-Z>�ArI4��5|��?��+,�̨���`w�=�m��Dx�JdqA�� �C ����	`�7#���A$��8��� �ǎ�uΎ���\p;(gmc�m�W|����53�OZ�6}B"������A�eh4�)�����h:O���`f	��ac�iA�R�����������/c2d� Z"�.C��������U]W���l���[Z�m3�򃉫�(�O2^�lhT�o�҃���%�^�|o�t���
m� G{V�1�/�M������#����)��Ԓ�o҂��pn<�z�Bx���O�#ڗ��3T$ٽ��8M,���	{-T���6x4���{y�MpW�U����#�S�+Z��5֞�ޒ<�,P����G���J�3`��h�χC��/�_{��5>b��vԐSi���8���\.'�s�?�%gw�F�2K���_N�y���'e��Rk�vB�4�umNh�2�����M�|nŬa'�Cj���>���Jg��hm����� ��i0&V��~1�n���*+t����$�4����Z˞�G�$3�D�X'c9����X��i����� f��u��(��[2O~N�j^8f��RI�xKέ{���N����K��
���1p�R��)0؝$u�0:˞=Sb;Z�]Gxe[�>DÛ�p2���l�/>s�D��Q�����08?0�
l��/Y��;�|�-��֐���Jɣ��M���o$oS�-
�M(:埤���"b.�v����VLTT����ۭ�ON��&k�7ؙ� ��)F[]���x͢@�\�1�ц��ј٩B8ě���2Q�u�*޴RݱM>�;��O��K��pT����:@�����%�$J�����G�v���^eK��z��|T?���=��RUB�\�?��ʧ�qzEcS��i8�竘!�m=ձȲj���@'�%�[;���X�l�Օ>��H��8R�IXd/�H���9��&�����l��`"��[����wК����A���@\3�x�_��+��̑����)�\�y�<j\xV�vio�@��{(x2�j�7e<;t��터��=��i�P�D�l�'e��T���Y�D_92 �M�B��f�_%1:j�oelY���o�;�1��c��ه̆@����
�	�#8)l�}��l���Y�@�L)��c����W2QG��������EтA��|�����5B@�����s�F�޲�~O�d�����L^6B�^�7�2�J��:t�B��?��v�<c������п��o�bk#fI5@}M!��G�EϏ�����Sْ�G�k��*S�CC��嫮��|e�;?�������@��)Y��L�b6�����m��xn}��2�	�:-�#_�x| {��E@����׆@�t1���U��E��n+b4R���xfq�>��Н(ȲN�R;g��8�lѼV��� M�b��3�|��C5�A�O']6�簿T��D�f�������FcDu���|p��N�E��t%D�������/�U�>�RI����3�S�	+m�trN���&��]K��i�� ��<Z ���P�+�C?��nc�0Z$���~K��Vs��G=lqv#SV�7�����������v�9�}Ҷ6�׽�bm���|�7I����L��5n�(���{>/�Լu�,g���!�_����׵�T]�� �}��a��D>2DT�L.-G�#`�V�. g��%���[��Z�e����P�r[Q]�&���,�D3qHzk&:h���hs�����,d�rw�z�Vh%��UWϱ���O�ą�Yd�g�e�-{�!
Kl�S�)��8�� ������f}@�,�-G�(�b��kOԅcqϫ���{�ףB 2g���5i ���y�pS<,<���
�B���=��)x~b.,�K������/�K�Кol߳k%$e>�φ�`>�ڌ-Aw��O����T+@B�5����Z������[��T��Э����ʁ�֚@�����T��H�XV�j�^���{�岻��	*�ō�T2����s�*x� ��E�����m��6�N��c4�B,�~S����F6��A~�(Z���)A#�"Z����(ø��	]�i{��"�e9�-z5�����['6&������k�j1e̤�D�e�ě;�y��s*e.�f�ĿJB\��4�L$ʢ��~&P�̈́X�7�ctC�D��؍��K���'o���E�?޻�����̕�^���M�Kp^۽��2�aC��������_l��|�����C�k�p�yp1�]|�Y!9�{�@LXN��reU���B�L�n��L��h���&��(�v�ĸ-�NZ�?�.�7�"7��\8O�`��p�m{�Z���[[�B���"1��ӥ�,/�2��@��P���,�4*�tev�����R�=���n��NC-׈�7��z��E��� Bħv�H��@��%�#���RN����>T�6�b���c�>�w �P@�/l��}Z5:.���:�j���'�
:��7m��"Z�틐[��"�x����ځ�0�q�-%�*|��ZiԮ�xN�<�	Ժ>�Z��nJ"AU���u/G&�Uj�j���N�"C��ܶ;ϖ�.�dV���Lj������\�u�O>
��\9W.��?YP��@�"b�."��p���� W�;L���7��O�}!%�r��ܐ��#���\*��@;=�mڥdM�*z5eN�L"6�̭��C]�I�m���}?J��~����,�T9�&��	nr)#E��������"/T�M�G�kv�tp2T�����$��������H��ޯ�Ub��|���N�l�C�P���/�8Q��lj���89f��t�Eƭ���Ĥ��-I�2��>] {Ì���j�H~�l{����c��*�>�:���͓|'յeC�bä�K�!�|����Ћq)��ʼ�\=,�H�m%�����g5�2֜(����X8��,��P��i�Va����x�IG�D����j�v~)0_5;e��z���Z��ћH<^����S�����,C�_,��g8u�k���a���;w$��*9���|�b(yZc�+p/�&p�df�K�
Q�F��<�_Xuo����/�'��뒸�e{��y��7��\������o}��x[�Hv����z�U��8���^IKy�����86�*��������>��G|*����cNR�+[&�w���-`�����5ڂ�r6�<�GYl� �D����������O��v.��������x�)XdYD��蛒��tc���P*�Wm4^��vϤьx�/�ӭɨ_���h�d�;"��a3�~����a?<+�@��R�6&�g�S�8tn/wl��R ��3��S4�1$q�)M�Su�s��|x�)���$��9`�o��k�0�Z(������w��ZCF_�S]q����O���%�?��|�L��C._X�@3	|�-+�D,����IS�*=��p�V�x�LR���ջ�щlh�˯��|�ѯr��7/���o}���;���
����Cs��0�#:�+T���,�~Xj �#��u����]p��T�׀r���@4���
:Gq��ѧ��K���g�TÍK�RN9Ql��^�s���M����0l���q��m ;�L��C��FU������C� ���}5I���z�YK���b�q���5|�Q����g��j�,�_Q�Q�/�'T�!�>��i�����#�(�*�i�Q˒����:���	p��2xW�4�v�8I��;f�1T����j�}�y��_`Ӹ��������B����ǵ
ۛ�{����|����_����H�N�D�e`E�e� ����L?th=���U!�����0�i��[��h).|�~d�Vڣ��5�-���"O���ۀ�GUŗ)-X��ep<"�{��}O}<�
�{REX���p��1JYK5�ت$8
��ܙ��	BXk� ���7���$-�iZA!��w�����^���ԱW�(m-G�P�2� c<�z�[�8o���XQojdY�G����'�-g�e�g��6� �Dg�> ,��;_w���]!��;
G�.=�!��?b�f�8��M~�X�3*Va
˾��MQ��VFC4�`�<(���BDH_��4Ou7��g�[$Љ�$R��A�H�U����{r�����=�j;�(�Ҁ��1\��3���J�mbL�oT�{�?�%$\��=G,�ԜQS�e�ƲD?�,l^tI�DMuW�t�����5=b{�)~>�P;�;�n��h��{�5*�O^�o}������(":�J�w��L�bfH�°Tll��R3(y �yXӂ*�n��M,	2��1^~ۀon"�Xs��'�b�!BpLl��i��_8�U莬a���J:}�=S�����!w�Ñ'�%'D�ӏ��ItA�l~Wd��0�If�k���-L͌����F6B}�)��W{v��X&��Ϫ�߈�@���'M��������+����D.6�1�f���?�0����9���F*Ѕ8��oi�M���ҵ�?��n��&�TLI��l�v��O6<*�v���8-�A,:�@%_
pwRw����G�[���a��.�nw4w*�+��I�I�PV��=8���@A_p�7K[�Z�4�m�������qW���j�¶l�ۀ�[))ε�2u��H�����{���=�I���qi���8��+��!���j�nց�/���a=x�[���0&rwM��ځ)Jun�b��էatn��(��> ���ν|\Ԍ7RZ����Tt�.v���v�)��{�C�k#�2���efB���.%�����T���V]��x��!C2�>u����I�*�l.
�'G�� �c�~�1�r�
h=�S�7H�I��Ά��}c]pb��5����L��x2֬�櫨�^�dB�ή���.�B<A#�������1�)W�E���(NdKp5*].b8��:C�>N>o���h1����L4c��".�j���8���@�u�d��v:��΢;�WHſ���t��4� �\�ǡA%oI��if.�C�������e���[���k�_�T�t��}�'�"k��O�LPHy�c�A�|W(� ���|b.�K�K�\���Q�E[S�����k�=/�&/t��8�S]���o*Y�c���P@�c�qK��*�T2TW��/[�ď����3Zt��8�k��{K}!�����H�qs�"6;�����;�r�P�JXGQ��棧%_���f&�����gX'�
����4Ş�<�@ LO�;��K���`T�d���Ef�)��w(d{z�!H�[�/��+_>�C�\[�ߔ��<��]�Uۈ*ٲ �*�9dt�1�S�ƨ{O�lz"�>+�s��