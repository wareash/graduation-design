��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>hs�*�U��Q������5Ij@��voX�⑟MlyA���P�Aqh�ٲ�46�M �Iݞb����L�,n�	�ʥ�����ֈ��*�G�������|ՁＮ�g��n����6���ք�A$��M�xI�aN�̦�!��7�Ki�
W��|BB�a�`p�D�X��?��$���_SVˣ�u�.���3�tH@"�|�|��5.�h��0�D���i���Fp�����L�� �^7H�d�Ī���!M+鍡��M/�1c��߫_���M�<K�}Up{!>�!>:S�h�(�� ���_(��J=���#��B;�r�}�t�I�������/u��ޔ�{�Xݕ��Wt���[��mz�W���Qq��>b��!] ���d���{,�i�E��sXU�dVѾ��4/	�F ������ƽ�g2�ү�k��!#4���X�Zź��5�EL#�|o�vTF	
Y(�-/p���4�y��}��a&���B�������/��97ũ��h���v��ԧ$� px�k|���lg�~�w��ĸ< �[�Z1������X
~sa���p��
�3d�SR��M����ᰕ3���/*$\9����l�h���`<����R�Y�n^�!�qB�d@S��&,��o�G�L�-�L$V�u7���m��t��O73� ��2��p��]�u��є�9�h���&��8�k�����[5?%�n��o��vahZ]!��uz�8)� .Bz��C�2��K�������3�ʙAM&�C&��
�I�Q n��]�j���U�;���;�`�㤢�z1E��9w��D�BQ�=u.��&�,�4.,ھ����L;�҇��"�;���2����0t�7�]�����N��ID4P��]��u E�Yr=L^E�@���GC��O�/��H��f`�h�o��N�=���f�iI=\�@A�2�ݰ�=΢/6Dw��;�|���}A1;d��B~^9�콦Y�t�l��P]���{�����c�)x�������nx�s���j�0���?��LA�(z3���BlE�3���
����wo�e��^��/�!���b����\˻/�1��͙3����X��{}%����"��biֵY�:vJ̕�Œ��pP��<pNl�ο���d��è����k�9ӫ�pyJ�]�#�a{��b
����nD����q%a�ƾA�B�c��*���H
�Iw�3�v7ض�i1[;{׹����ů^��Z��S�$X�S�dm�b���]�}3��_R�e�V��d��-�h�K޺����6�)����r��~^�ч2 �+oy�"�� (&�O]�{�>�������X�/��daꡭ������ӯƋM��X� I4M�c���l�ML����bW,�)«�5[_�X�\i��t�$�}���KE�'_ .�IT�EPM��p-s�wM���P�	�����L�.�6@XQ&6��DLy�� �%p�A�.�l��Cj�xִ�+���������x���A�!ɇ�>�i�υ����J�������(������7��8�M#��\�(�#{ I�4��ڨ 9t'Q�X�X6�Y�� ��qɎ��Ԉ��x��%�U}[��3h��Ó`a�T�2�R���wmB2vH���7m�D��ak��=�.l�Μ��ľgr�p%�H�y3B?�.�MÌ��eT�Xq#���G�X���#9�5��y�*ǂ����:�8h�f����J�'�ٿr �}�6�ҷ}aT�v/�gW�3��3=��S�v_�{kɀ���i�m�Dp�Ҥ�.�Z��DQCق�F��P���m�F��R��4����NW�����Y�\4�F
��%��@N�K�pC�^=��! M �t�1����E�� ��@Ϩ��L;��V�+,��q��3���\���9��E"i�e�=�zS��C|¥N-�mܔ�{|�t��z�l�T��E��W�Bs�?ғn�����Rا��´�f�6�i��H�P������G�(-l&"�"��pW�5���r�E|�O%��R�N.q�cB��$����g����ۏ�*���������g�ӆ)�"���3��T3ۗ�⌖��Je��Gy��>gH��h���4ꖲ�ahB1�����׳���@T�χO�c��n������j�����h{����m�|��x�Sa)1�1��;�zp�\���N}w�y��֊�}(��
Kq�ei�9ۛ�.�7��J�����)]:S��x�{�T���Y��J�-�g2�" �/a>=}�\/��|u����J��_����O!2	��X���S�m�#�D�k�]2�b�>d��|rg�!���i�o>o�~� �F\(»桥f�V��LW�jH܅~���������ܤoS�B_d7��dƙ��6�z��˷��6O��y��aSH?�������-��a�B�V�c���Ef�G+�x�c�Xd�װ.���!~�����ax+Bh�n��:�@?�����}���
�0�������l�jF~� ����DW��1&��X�u2ٹR�!2U���qp��;���0���)6�`n�S�dC�ݤ�i��Vч�Q�6����DX�Nd�Gc�~�H0J��tpӕ7���܁��>��Ȃ�48���h$v��%�[l�k��q�7�%�ݷ�U��V�P�l�\���Ʌ}�)١X�]�G��R��n�h8�i��S]��9Ǐ�\+�z���y$r���Z�<�%`����N�2]�,3η<������|w�FD)�*����k�%Ӫѓ"߳;�xeu� H��O;F'*��68sg�%U$�ɦ��Md�4�����E9���[�ߺ���712A����(hM�Y����]� d�V��\���ɪ��N=5��ǌ?�2pI�$H1CN�#���-��a��� ��EE���%r��N<R�$��I۩]�(Jj��r�Z*r��W�l�D���PWG>h�o�@�S|����,�U$nT5%����#��#z��f����U�����q�E5-4è&�f+���=k-R}�	���9��0�(H��oo?	딣�,���Bl�S��I(�+���O�����pGuMA��}Q�(���z�*��[��?8^�-�5^2h�$��3������ɯ{;k&�!�F��ߒ�plL4吂(0XVK�<���&qJ��D�U�P��pU�=��-6����Q����X���y7Qװ����`�<���8(Y���^��6���bJFt�U�l��v�0O�8��c7��\�Ks���/�#�
��4�s�����fԗ�z���tyaG��*�{�\����� ��<�����X�y���R�V��T轜M��`T�(�f��An��N�s�������e2�.e��/C�D�`�oYQ}<�����������U��`Oo|h1˓!wO����nj�.��FQx������.��	+1�YǛ�}�A��(�]��"bB�D z���-&Q��A9�(��6�=�D�xl�%!��E�e&�ru��l:E_?���)�����	�֕���������]��0����B&����\��H���:K���������k꽃9H�a	t� �ְ�.��?-5�1b�q'`��P�͍��.�񻖁18c�E��T�2��( A��Xԇ�ͷ9#=^cv)��i�e�cA󴴧��r��ႅR���[Q��:WN�	1>s��qgJ��ȟ|c��q�5+v��g0o�:g@(����N(䰓����	��x�ir/�5�px��gSm�����Z�k˃����I(AL%����p_���t@f�����U�����T7rM~�>]:���~�]�5 �Ι,�j+)f�SA��'�������%~~/�tQ`�"������	�@�!�)��}}h5�ABO���QmmS����!�uGI�:�WEG��2f�d��y�2Z�����e�o�(����k�=�%7���7�:K�b����n��w(�#Q*�$x�b�B���A�
ʋ�{�OL�}�)�v�X�W'f?�λ���Ҳ?�#��\���Y��Ϸ"��Oa,�^���8�,�!�[sx���������NyTveWy��;e�4�ay�����P4Q������Ƴ��j�����ֿ���)�,���U�⩕�����m�a,�	�k��������el^�ҡ"}9�ni�Y��9�Y��f��ׇ)��1D��9+{K-�*�]��G�7hĠ|2�)yL����b�@�ir� o�D�����VlSo�EX���G���s��z�����t�^�7vȾHX�,�M��!�f"B�8��ӳ�cl�`=ӓ?��êo�B��\�!E˛^����g7�%e���:���Hh�26�9�V�ki8�`��J�F�6�ή�s�F�6��.fu$��x�s���(�T���T �~�����n5�A�%n�/(������[׏6�6������n���|����ĝf���G���My�V������N���:xz�p3�7Y�|��'��J��ok�L�(,�������{j�(��^�E�%��tr�x�g9!������$�ʜ?I֡9ݒ�}��TmQϭ�r�?�?���;�!O�7@��e>~ɳ�Y����竜���5��_ƃc���,���DD%1� �YB�Lo��rः�u��[�|:^ی����1m)� .�=�I^7@����34����:��v:S�;[q�������E!F�L�X��%�%r�Sh���XW.�G��Zׇ�[��S����P����x_t��������~o�d���Z��:��F����q\r������Y� ��_?��,A�)cE���S��aM�g9���je}�	`۷@M����ck����1��12��8�6
M���A�dH7r@�v<Y�����+�	m>����[l�dȵ;�S�w&K�{��m���ê�&��3{������z�%*0�g�� ��I9DB����Q;Eԯ�;;��������%������t:e$v��f�ڮ��k@�ӻu���������Dh�����!����֒����P�H�� ���k��M麲����W��o���
�5��}�$�L"�-�+0!y.
������6�b�)R�f�8��;X���&uF�Bv�a#PZ�8q��?��{��~�� m0�u���ʝ%�H���W(��/�m���^y�uS\C���ޏĉO֡Jy?=�ȫ���BD���
TԨ�h�π�V����Iw�Q��� ����Q������ɇ�e4 ��
�os�W�!8��=A��	1��	�/7� ��yS�|�u/S�Y���d���!_�:"�~��M
�!mc��r*�օ���B�;��a#0�����E�<|3�7��ZI+��w�b�����m�%8�V@�߽ib	!<���7V�n
#)v/�_X���
��,rLtn���ו���F�ދ'��RD�wm9�_��:a�7�X�W�Ywr�b^�\� (m��ǃJ�|��ւ���烁�����o/�֫��^\|����Mg�xf�3������i$A����=���L�2f)���_�]H6�C�}r�P��-[����� ��U��)��	1�&��k Trx��N�'!D�s�2��M�G�>J�����k�N-��%KE�b�͐<ꉁ	��d��k�F����j[e8��@�#����̿�'b�S��V�)�6Y���$A�x����#�T��V��r忴������u�
�H��-��k=�v�QK��	T��x��`ZS���u�G�o'\�Z�1W��`�B	�¼���d'ZJ��#}h)�%�~��A��wl�d���Z�]Q�j �b�Q_�7H������&t�e�P�ÏW,�����29;���r�ǉ��)&�[Qi|Uh�b2
��c!3_yG���{�@�jFj�/G3�>��=�si��k�ݥd�5n��Y\��-�u\�޸�|yL���_�|s?��cp��rw���b�����b�1t��m���x��8���|�o
V�~Þ�e0�g���3��	���'z�I�$N�Q�|����Z���jqF���5�#���~�N�˹��`��1n<���?���Z�)&�i��b�*���;G�����]ٵ8�V�_�d�BEɞ�ݙR!��A���c�5��B]�,v�L��Qx^��-蘷�u�C�}�㘿� 	�R{Ɋl�\XC�w如�9:R7T�t~�����$	]s��Q�uwr����n�2�s3�ݒE�z�HK����}n�abn�I���xf"e�0��Λ���K�%�˚�~���;��/ ��b�I�o0Nn[൵V^�r`y?c��~%�L���W^rf���h��S�W�k�н���B�������1n�^SUgS,Uk�(�=C�Y�[Cr���e�4
V����WrC`�!կ�#�w�	{���_M�- 對!�g!��ʶEI���TuLY:)��6��^+�a�F�6� �}ēM�u׌����M�k��á9�|<s�w����PJbo���=�3~���4C�v��R�a�B�ȝe�%��Mߘ �z��3��+��A��|Oh2 ���hg�>�ƴi�ϱ=�1�A���L8�������V�Tߙ3��Xt�;�@
]�=۝S��1��]���W��i�P���caZeX�g��,�z��R��G�gؘ�P&��T�ZA�+{,����E��q�ԏ�S?
���H������5@�Q�=|��q;~�J��r��7��c��(�`�?����_n7��2��'�A�۴+xa��1�1�0��%��}y���fr���=ㅑ��d�۟⍯J2�[ڝc���F�S�r��e!�]
^=��ï�N�Ka.�"��w"�9��&(I��C�ˆ������FHc���vy��� �����xU9�����L��L:����L�d��
%X�D�n�E�l�Bl(<�]���A�3��l�EWi�XG3�B
8���+�	���PK������ ��]�l	.�GZ0{�`^(_�+ ���|��})T��I��x��g��|�a�b�J�nË�4!���-�����ҭأ.t���5e����#��g�p9�au�����L@�ah`j�j,&�J޼�)`���)L�M؄ �������gy>㕝Ԧ[0mסO! \6��8�|�j�2� �5P�s3%��3ٔ�J<Η$������CHR��ߌ����D�>L�l�:Yi�����h@r?jӡ���f�U�=��d�vmw�]�Ga���lY��kIP+�3_�Z�55t��?����B���Ū��ނ���O���{gN�E�n��*�
��G��[,od�6�u�'�1/A9�������6Z��x5��y�M�i�Rf���\9�:ۆ��B7ÑS5cI�G,�ȕxY~���#�Z`y�Xy�,U�����X�_�m��<Y����1@�4C�e���&�+7j�׿;��eC�M�ꪩjG��<�d�jK?Ѽ���B p���^����`�F�>uv���}c��}�؄�AF��2��)��NE�ބ�j�v#i�J���W�>�>{�/J�hɡ�2u�@w���Jt�������j�2��ܭ�