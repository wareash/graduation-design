��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����)n �n�NP/x,�Fu��D,�C�)��j�vR�������|�]K�U;���A@A�qY@@բ���e�̍�gF<E�0�z� n��Yaex�1��p�+ [�B��;$ţ!
�_�c�>�Ή4�k-�e�M�}Y.tצ"[^`㻬Kg(5�f��#��D-s�q:�0eP�%����+���ݐ��j\�8��n�p������xo��|�v ��o���o�4,٫'.Kq��$�q��\�6R
4�q0����R�R� :P~�آ@�����Sx,[��0�$���E7ٷP�g����w��Ϗ?\x��%�2Ç�n�Z������eʔ�/�w(¦.o��z�2y�m��#��S�F:�..!U1��#U"�SF��A~S#��?;�
�~&�Ҝ*��N*D��bg�K�JsL�ql���dD���p�1�79F�ryσ��zp�+���W(`$� ���Mk�S�<6����%ү!LxGp�̓\�J7M��d��$ �)�.$JxK��\)�ZU�<!�R������#_�r-q�HJrEѢ�*�C:�&�D~�/���F�������^����S�C[;�Z�5����RŤ�Q�a��ߺ�b����+t��h�]�*Ԑ�;��C#��]�r����2���?]�g��Ϛh�D�;�<��l��W��4hJ>NeH.ř�!?=x,����p��dAdp��}�X�=���y �w�S����0C3U����&;5E�� �����>�ݢo��Vr�����m�4��q�=��Ҧ+$�HIgKp�PB�F}6��GXz���x��b��)~#�_�U#�=4����q�ȣ�&P@ ^\����(L��V�:�������e��`�R�Q*���=W1&�ݳ��C��b�k�,F3��2	]�]^�-��ʯ;fg��GG�7f�.��~i��������Fچ����I$�Y�@�Ӈs�d7h�)~.���0���t�h�:�����8m�Z�"��Oޏ_8��n�B"kk�|�TƢWv�S3y?��ߨ㳦D���2e|
���Z��"ĭt҄�X�����Z�W�Z^~wx]b�[�+i-ja�T/�"(���Ѕ�K<e㹌��N9���Q���G���e<�ˉbbN�ۀp@��1�b��Q8�u��?�����^�*���"��C&@&$sW���T��_F��ǌ~��X��cY�x��6�#����k�w��M�y�0۰'�������A��z��(���F��=��������]@c���N�m�mQ��3BN�,��|�oq]J�l'�+_SON?� ��ߩI�^�v��+G���t\�zR<ْi	w���	f4�q-��V�,��.9�KH+�u�zM�2ro�n�b���DNU2�X��[8��`��w����0dbjB'����;���l,J��CDSﻧ���߃w[&���{�;��D.ƀ�9�=A�PO���ԇ�	�&�e�{�)[Gw��~u�$mhL�L�
����Q�����Y���"pv�?�V�g��&� q�/��<�2D;����"=����R��6h�u���U!����O[��q%��W��q5�"��eP>�g���=#�,7�A4I��=tL8��Ƃ�K�Sv#�OS�J��yE永�MB��җ��G[:���7>,P�
�l|���&8Z���; ��ܮ�LŒ�I��X�F�C�޹W�=ɧ'�2#$����<T�^;ƛe�J�z����a�6����@Ŗ��wA��Ǧ<�]�yP�޽B��J�נ�ҋp0��ŭht۪�I��<����Nq�	�0�6��	4'�39qa�Ug�� b�?[�[r�j񬝖�yS��Oǟ��@�u�N����߲�: ��S̵�V��K-6�ۄ�t�ܞB4�>t����
�IX�R�S��d0�@�8 �РVPF9LC�e��?̝9����>t��n�N�jqTE�0�Z{���ch��&px�Ȝ2-z���s@?Y��uIqu�_�X�ԓ}GȌ��_�Ln@���['eYF���C�0����C����hy��>��.ppd�C�{��"�k�J�T.T4O��vS�0䜶��]�(/\�AG ��7�6�&�`��ʒ�5����������H�s�ރ�?�+*-!�T����
�Vg[�,} �🎽- %̲;����Z�􎢋:��X.&�۷B���W������Ku���gf0�4�� �/���L���½�>!�)4|y���<m���$v������)-A��s���`i�"��q��Ql��J�O��nb)Ύ���^�@O���>��	In!`�.Q�9	.����hzyE4M�� %�R��c��A�&��ۧ�p.�]�T[YِL�������������i�ڸ���>��HK�ec*��W���&��@�jxд�iL︆֥ eЪ|L��cTR�r����Z>tY*��2�NeHd��Cha�Uv�v�vO0����%eXq�6��׿��\0���(��IU���@K��X~$y���5#����ϐ�k�E(�d��M)_0�$��X����4�N�!S2}����l��Boi폯�-�C9"��;X�_C�
j�Wp�A�[r��b����;�5��:�t%a^Ѕ�nZ����0��~�[]��h�%㲵"��(�ѭ����
�L�z/~�E&�p�M���*q���� �ǜڑo�zh����'��փ�����
X7�����q{j���P�Ke��4r?����>;cIo�;�Ǚ1�R$[p�����`����Y�\�q����5�DԢ�-Z�aV�ц���y�Q��,vD�}_�jn��*�ٝ�v|ΚS�f�v�1�X�-���W>��̇x}iJ� #Ϲ�ԓ)ܘo�F͇�K��g9�H�R�<_�������
!!c��*�~C>���P̨���/?>��䔾�%����D����A; ��7O��F`���bu�~���nޠ�ˢs1�+&�j���i�{�wzt�@��zy�fs6{"	P!])O���mu>]K�Aͭ��Μu@���3���;��X(�G['�!.%���a�b��,���a�W�"a���928a���,�Y�V���{��H.*��˓��:
<&�f� �I� ���)��v�0m<�<�	��"L_8�Q鬵v�F����UT�z����򙨉�vT�M�[��<�^Q���wb3��Si����:,��+�����ku� ��>D�\�w=���?/�*$����l=�lU\l)�[��8���L$�#�e 9s�b��J����֥K��Z �����,R��,t2O��Ǧog���v�icH�0���2��'+(T0�ƀ���`���+��֛ߨ�y̒�����z��Lb����L������M�BP��WL֒�q��l���ؠa5-=.�#�SM�9h�8���ѱ��X���2�!bɗ	f�\����6`I�����5k)�Qy��C(�a��a�M�7����LW02����Qk�s\�'؄�q�ޓ�|C���ć�\7
J��b�oѶ6�������
�O��l���vҘ>�VI�����?�q*A�t�c@��b�md���^!Z��R<��S�3I��Mn>�"����E������Da��Aг�c�?�|��,{atM����cf��j��Z�J"�>%�f��#���b��¤�9t�� �d��\L��ޟZ��glc�)�n<ɥ��b��9.���9W�I?�
<3@E���Q��"ūf�m���sY�~0���8n�S�N)C�F;�m�Rv%V�=����`tWe�V���2��vc�.��&���ة$��W��]�-h�zK�O�\�?|�<�?Q�&����:F�OD���"�!���
�^�^�;�<��Q>�9���g��h1=P��<C7��r�n����	^�|Km���a���jrTO�Y��*��7�I(�F�:I���څ-�*���fF���Z>��(לG�P�¦h�v�tR*d�������A�H�1B ����<b������������^ @����~I�<.���HnQضXj��Gʈ!�Ł�q���˸Oo��B� 2�PV������<��@����Z�U&�H�ʝ`Ľ��9Gg%B��0ߺ10��ޢ�DH]�+W�̮�x�wG$�V�>�No���4�T[B���hF �$i�y�9�L>w��p���߲�{Դ�;�fU`_��fZ�I�|�?̽n��F,�{Z�S��i��~V�h���y��q0��oMo�.�Ig�G-K��6U���Y1�6�R����"�GbZ�c�5��Ǔ�