��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jåا{�\�u�?߷�dn@6�zf��r������;,��o+�[�"�<,!���I��F]ù�?�o�b�v\�O�����������3�5����e��7G�v'�;@̀ЭwSF�׬�
�j�J��Y���[������Q��ߌZ��X�-
�U��e�ag�ܔ:x����R)���ό������h��
�Bz��Bl;-��y �Dh��Om��إ8iT���s�,i-��J���Gq�8�F�w�cP����R�#��V��@���w�*��������K�-�������%�c�O����]��kw#�$�����ENq�g7]���#����\#3P<��܅��*�Y輖 �S�ϳ�̳5��匒���w��w�?��s�U�OD[݈yp�K��DY�VȬ���/x61��I2�%�l
�r	�'I%�{#�>�CO�_�u�b��B-�A �������\�p�zOA#�ć��c��3	("�Oe߅�m��S�ϲ�^�;��7}+���c�������u�?\oy���|2�`�r���ÞЭ�d(gn`q�̑�Ǳ��С���n�q��L/z�.N��n�!gL߰�ո:=te{���q�	�Y�F@�79��F��B�B��-��G�/�TWi��0Xɕ���XM�y��͏a�x��o���.��yv�bS�Y�Wg�����]�K�k��Y��j�!����'�|���:WO�#�O
Ƥ��ڱ��q;��)W'���<�,A7ӻj�� i`9<�Ғ~��T�H9C��{3 åؠ鸨G2���ѰO�=W����.�f0�!����p�,֒�L�ˍ�-��x"���P35Ie��ѷ�.����C��)R�P2:�j�O,����V#|I�3*&l>���3�X�+78?x#�ړm�j���;�	h�I{2�cT�����x�et���h޿���퍩}��U���[�O��谹 P�~Ib��xr}������H�gn�'F�v��{U�a8=N�m(h��0�z�xbwnq�C�x��K����m\e�#�Ҍ�!�$�y���~|^��gʅ���$($:^�{��?�kj��4�+��n�E��B���G�w�����٭n~|��g�In̈́H�5���I!����%��ֲ*��s5�Q���ray2g�d�p%��]_s�1xn�@���z,��"�@�.��s����}&�����;u���Y�F4qa۴���gH��8��,E��r��/E!+�qU���+�Y��Wi�0*.�G�$�(�Q(��KX]��/u�a5@�6�F�G�������_�,=�w�6:��.���D:e�������`��]�	�����߉%�j�:i��)�����:�߶t�(�ٵ��ۄI��*DEV
n�jz�zz����U��{#���d^w�$���'�X;#�"�Z���~U���ӭO�9��C��^�J&�{'$B����&]����ȿ��櫛��GQ���s�:�gY?���K������ɉ�J�޻�L]vZ�+D�f�^����?Z�� Ɲ�r������rf��q�j��sd��?�IG�Sу)��HN[C��o=���%,T=
5R�.x�ӹZ8DSL�[r 36˱�7�28's%�OQ"�֟_��o�������%u��_ ��.Z8Db�����K� <{ޡM�+B�\h�w�	T�Ǆ�2�}��Dt@2Y0ng����Z��|@~���k��I�������*+5y<�$�w��E�W���}��&�C���,Ƃ���"V��9�k $D�\U����w׆!��G�濞�{=|t��?�;\�k�Cl����7_��Y[��t��\��?��j��٧Qu�����~Ho煰��M�|�Z�g�V㣎	~�O��S�)�u7u���~�zu7��b�S{f�̀1i[<
�ʎQ��ޝ^�Ȑ��c�O��|.A��Y��(��M8	m�4Nzb�ٶ�w9 `|��l�kw~���ҟZ\�a{;��Lu���~bC��0^L-+�O�&������Q�,
��:'��]�������*Ė֑�BFxmݰ��K���L_A���-���Z��g�D�V%�H�x`������R������׾�Y-�Q�l��۾:��'U�~<-�yŕ�>��fݎ3z^|�Gl{Mރ �Ͷ��iV0q�2�v����;M;��e@m����ڤ* �%?ρ�]j[��L�����Y��ã�jy����'�'Ƈ.< ���6��C���B�B1h�f�|$��H8�gZ���:#�a�89/Um�g�DD)HN"�O��q_��� }|yM%H
��&s�틛��h���xN�x�?d�2���D	PѲ���\�B����RB��+y�Kk)�rKhUk$�%z3��[�	�g�������~>�JM����DD�+���{�]���Q�8��@Z���p޼b�0y���Q���v����}�~�Q�n5
����T��|jJ>�r�*�����K�r^�1So����/s?�,�Yh��uE�w���[���jcˌ"L���4�+��֙�~�����)��Ȟt���<�ϕ��9���-�ҹ�|�������W����q����=�Jq�룥����qf��W�%'W�������!U=ɿ�8���D �����U xX1�_�z!.�����zг^�J��d���9W��n/�1��tIQ-���C����To� �!H�hPǞ��J	A��j�e r�B�V�pj~޴��}:>G$v*��X̮�.
U�jӟ��z�u�bP����d���9�W"Լ��Q��ET�,� h���ڴ}Ĕd��ުN�ҡw��Ubl>�!Þq�qd��h�2�l���oݮ_Ϸ�E�Xc���Ҋ-Ne?��2�u_��ʺ*�I$ ��d��ދ]b�~��_��j���Bp���ݧ�����!��2���X��Ax�?���H�o6�Y9:��w^�<1�@=d�-�-mfx�
� ����g�w��e=��R������߫Lu� �o��0>n*��6lut>A�s���Og�G_���PZ2v�q�X��m��D�� ��O
�A���>Lq&���ɗ�k¨�`sL@��D��P%m����b�a���:���U4��է�m}�0�#�����b)2����c�eu��"~�<a1ѻH����֖�1v�s�vM�ʄ�7d@�Vt��{��	�� I��K������*�η`��"]5�5[w�K���mU��;��"i�:��HƉ���&S���Ƕ2�ܕ�����(�[�����|�@$Jx�j�o`�):���Y �i�C�������|;�p�3�û��[�u?���VB���W�L3ޭ#�`��G O�SA\[�T��W�u��(��:�U]!	\�����Ő���YM�[!���&��$��<),;��O[מ^�I�e���5�fj����#ŉ�NN)���`EjG�p��f:���/�!4��k���-(3�uN��#z����u �O�q��ۿ���Mcn�<U���"�u1+!kW�O֓�,��Z<�A�W���Yk�}�5�I锋Ad�	�;��%c�e,	b,㬅LK��Ib)��!3rq��(��֫zX�zS^$]&��j�!.7��4+����fz�I���S����ز qL�˸��E[#�ၰ�L9���r�K��H��L���� ��L��M�@���R��E�,E0 �~���/�}�M���#�|Ty}���4���A���
ռ�>���&( ��X�L���?�0�e��Zܽ��DP�����a��	��$�󆇉0�U�Պ���M�/�TՋ?���,��4�t4����A��_���>�mK��z`�X}J쒦�A8>+��̶�e�/``M�z��i�&�����w����&��ڪ�'�l �R=(.�:��sUf�_5���|��(S:���*�F�X�S��)A�9�o��!�:9�����V��w:E��zƍ,��'95��:��ꁞ6�)I� &8�`"�[P�YZV���ߪ��.�O�_�蘣��R��)E(��:|Ǟ. 7�t��:3t���#��i�ȐeB; FH���Κ�Pa�:�K�5�p+� �uҍ(j���'�� <|5�Z����y�N%�H��؟�g\�v�?�粛f��$��ch���5 X3�:<��b�3��4�*�C_�8RXŖ�=m�JP����[=�s�x:d���E�^[
3�Rc�\��E"�y/������:�T�[ �)}�.J�eҖ)��=R�*7~�|@t��6[���eD���X�<�D�ъc:L5�v
0�H��C�2w"7e|��I�X�E��;H�]$W�Z�7t���X#���0���_S���n��D6ހ�'}쥖�qR�ud��&�M�� �bmer�5�z88�і�p�~��3�iy$i��P*�0 }��c�r��*�&nK1���.��$G�P���Rs���9a]d��9eN�3����A�;җ��uxѳ.����C��V)	Ҡ�����_�f#U�>�.�#����"_E���ab��f�h�?i��5��}n�7m{wq�M�&a_J����h�H��'߼�^y��3|�L���]I��˅G�ϜMе^E�lU.l#��@(vU�6��B�F5�`�i���i�7�#}����s�o;O$z]�����{ �La{]��'��2g������t8WV:�n��F*�)���;��s��YrSK�y�k�*
��j���4\ uR�g_�Ң�`'���V6FnC��mm��ҟ#����xK��Q�Xe	tB]>��j�ȡV(�=b�i�����J�Q}l�s��e�xцV_G�(��r�f#�e����Oϱ�����D�S�r�M7+��ő2\�w��go.�Is^�j��ĉ�g�d"��άO�D�APC�m��"k�WD�a��%Nm����z� ���,I�rZ�A���*Yi�T#<J�d\��R�L(��x�*=����l�#�Ac#��v�muxS����#%�����!v;��(��HvCZ�_t�(�:'A������-_��}s�9J� ���� �
��ߝJ��oD�!XqeEy#g� 
J�0e�Ê"�^��fgq�~�gD�|g��td��h�ʂA�t�Es��Q{������E�<n��߼?�u[׮u��!A�3�ܑ껆�w��7ui���H����>Jv��s(�����Y��e<�9���X���N`���b�ɥx���~m�8|Ǟ���>$q©��B~ 0�c9=h@�������0�p��g�A���%����HG֜zw,��*cL'�ׂ�$�s��,,)5��z؍����c�PrLI#�h��Ps��7M��u�2���C�j�ɱ<Z'	oP�����x����!�V��y�M�}����j� ��Kԏނ����"�'���/�z9��)���拘��A�8��[fxZ���������ޭ� v<�,.���X�iC���[����S�E�(��Ms�Ƣp�8��XޯXh&u�X���t�_�W�O�юv��g��=n�<4(��L�繆�;��K��鳷Ǡ��az���4}���Y�Oٻ*��WK�P}-�}�����`[/�f��W_]������i�VW��g*]_�!E��j�Ƌ�x��4$VM����j�ώ��.D/��͠s/��>��8�K	KE�G�6��λ�9� ����V$&qz�+D�	 �1im�F�
�`���0��H���H��(j��L1bT�Q���q	cN/��u�^�J׿az���g�l!uȺ�De�q�ҥ{T0OݬBZ�A��o�]�,������[��Zo�
�%J7���7�� G�Q����H��X��>���ŹĂk���č�2�Z���u����P�{�U5�E��� ����[1I�\�ف�X��M't=A�0 ��s�Ȱ,n�,{NK�W�h���P(l�t�r�K
X�j�9���3��5*=�?ՈO�q��z��X��6v9L�uRÏ V�u��ܚ�<��sF��,䀗����{Q��|"�$c�S�4�<�^������H�b�q�]%�u^9@^{�#E��@�a�^� �^�p~U�ء���p�9+~�b�ۊm��y&��OMhU谀�:��c�͕�UΊ���fZ�%YÄ0�8^�"������Z�n�^�7�(���"R�0�HZ�zq���`tz�J����Rp��:��������H����V�pXm$D�2"eb`�B�Y.y�q�0���--����ն�s����*�ԁ�a�Q���(D^:�ס����qRgw��O��V6LD��W喝(��et���t��$�V��?��K���Rg,���$�ϭ����xݤ�v�(��;��1�[�M�mJka+'������Qx@�}�A&�p����2�Cb7��PaȄ�
�|q��%��*eU��0�!��F�T��	%�+��s	�� A�8�=����l|�韒�mq'u��h 1���98�b
)�X��YK+��Ж�Y �*5��2)����||��o�e�ku�hW��P�#ِ9GQ��)�=@tX�4�q`�b!ץpr�xi�v�i,+u�ZhF�V�qV�)�/eW�H��N��[��Bi�c�!*@���	�(��{W��w�e��p~T��.�7Y隸=K��Fr��%�J[1�/�^���i��p%\P+��:�y.ߝGY�P��M��Fcc�~ntb��e����,[�T��5i5,��kOc����|]�hN�>���%���$H� Oh����6���Z��ed�;VQ�U
�gu��G�QND���,#�f�;�4dbt� U��{�e���H�ưM�7ӳE�A�a9����/?��.њ0����%a��qH�M�/$�)0����p@s1��i,��h�}-q��E�غ�9N���q&v�8�[1GI�d��CŞϘmV#W�����}����Ҧ;������<�%¸��W\���E~쯐'�^��8�t#`�0�hxp!._�{���%"w��4�����z9kγAg3:�R0��؋�[P��hɪ�Ia/+�}֊zI�ȧi�V^���˸��$�֝ᎆ��X_u�>Kz�Y�,a���������M[>��3"�>�����0e�4h�`HjJI�^PH�3�����No�!�Q����N��o�jt���:){�_��,��'��b��p�U�A8��M���{m5��Q>��'V�h>�IuQ���x^�$k���M�C���/��'��e�/�� ����~/��!6bT�;��/�.�B�������X���1�L?
�'��
�x�\�l�U�.G|�W9��̲X�˲{C�� 4�/� �z��W��,B ��;y �V�z ��,��۸��Eu��A_kC�S�(T���]�<���:g�d�^��ݳ�f�P��_����Kuu����Ja���)����z�f��Ԟ�{􃆿!�lX�����:'���іr���89�+��*3[[��jt��sAf�4�9d���-T�����9ڴ	SH1��Wb�"�M�G��<2�y�G�y�l�\� ���%͵F/�3�ڞ|�׸1@A���B���A�=������nMk��h 	*��U��������0z���@g3�`�g)�㇯Q��F�,�1�z�^mi�;�V���4���4VJQ:�>{���ۏ��Ov3:Z�_X�l ����,rIk�.���Syի7�	f'�籣jT���ƃ�w��ߙ�$�G�{��돭��nb�J���[-{�6�l�zͻ� s��e���*��Ӎ�^�Y�vi)#*�A	�ހ�ϫ��T��D�Z0#�ɣUs�2�,�Xb��K{��*-�Ӱ(�g����k� �5׊4�W�_��d���-K\1R�u�B5	`�0]���{�S|���b@�`���`���V!�=�[�yk�{'���9�b����l�c))i�l	d��kMz�	����Pdfz��!�s;|9��g��e�X�����a}��8����.`^g��7�m�A�o����X�� ��4Js�'�U�
�Vh��LJm��E��c���r�r�~4ax�N7����p��� �`+��`S$�1�'����,�(��U����� ?�6�(�)����g���e��I�Չ��9^��z����H��ʑP�P� 8�G8�Z�@hi�뚝�)�f4��n�rǮ��8y�Y�^�[.�gS\�����f����`D�f�0"��7��3�V�9Κ�͞o4'�K���!f4!����#�w
 8�O4���u_s->��=���g�L�Ȳ�&����i�<ʺ�C&��5F���z(6j�_�wZL���q[lWw����FX<ye�;p"�(��@D�Q�Z�iN�Π"�4i{�[�CC�\}M2^ K���cW���Z�yͫ�KYUW��'T����Z�F��9��Ll(hUM�`bR �8(9�<0�� l��>�s+S7�[_u�8���TsHEq����� �&�NT��k��N��mޜ7p�c���,��e4�e�v����n4r�lV�Db$�Ԑ��)<a���"{���%I�C�V���x����!)f\Q�_0��yԫ�f,{�T���M<�?�uW�"�yw_6�+�G�ׇ��c���E��D���ȝ�j���#N��/ۭ�ޤRN�X
���3O��&��g���﬈+�����$(媫��Z���e�i]��> �2��lU�\��J��
G�)Ը�Pe�ר��=#�-�Q��im�\D��5Y�����)�AS��^��;3k�����/ʢ�-"Y�ʇ��$���Z1g��ւ����#�3�a��_���!���n���W�O�yM�B���#������\�!�<uZ�F]k@@s��,�8�t��c�"t5�T 5�K�^�2.��w>�ɮ&�\P��͟�J�
����0�Z�+�-
O�.w��4S��,�������b�~� ���]r�	��+)�|�$WLk��%)��t?����:��p��y�4 to���@7�śo$��aҔ��@�y�kh�^�u+�F[��!׷�8a�T�a���q\��ܼ�Wu�B*3�Z��K�ٹ�����E7�q&��h����H�8Ud&�n-�֧�kΈ? F�����yQ���O"}$X�s�Й�]IʊN�G����ޥ#,n�&�t��D{�����l� ���cl%���wJ��*;|��k*�:��)źbTLm�E0{�
Х�W	*����h��z�ԃA3�/�k��S��O�/����S�����a80G,���	�=�J��b���NOW}h�z��U�����$ގb`._���'R����n
0T�^��s��],XG<^Cb}�%���ܽ�ʼ_:��&�YC�x����#&�DH���?�|b��֭��fd�W�#�pA�d-�yu��I�vv�2-R>���2��b��uh��n@��-��\Zk�V����^#����u���_�^�llЧ�+u���gTp3����#/�>�!ZZ`��H��f�!ľ�j�#wDv��	҄s�m�]ًx�N�+�ϭ�'��7Ł�p��<�l�A>���ǑP�VB���i[�i\W2���y�	�׋,���9vz�	᭏�#����K�E=ʱU>C1����#������Β���fP\����t����|�@%07���<0tʣS�z�đ=F5fo>���#��u�yj����7uD���O)|Pl��r�Vy@���\���X�r�$�1\���6��b(�d&G�-�@��z��v�l#���<���A���!�S0�Hv�wɍ��{YeG.I�M�n�A�2-}����g���\2�H	K]�N��fL���=�2��k�*�ׯ�0�y���3���!����]�L9ͫX����Npˊ��	�&��U���L��\M�I�Y�'Ę��̨�*9�l��W��h��Ҕ�c�M~�(UqO9It���;��$��~�/x�� �4)�*&A�~"+���sN�KLe�s�7�G�]�����ܣuI��������.���	����-9y.�L\
H��L�(:�*HJT�jd(���=�Ƴ �,�U�N��LnG�<]��%��c��eվCN�&��=�}���Q��"A��`�5ե�^h�dC��(��:���n4r%H+c��N;x�}Gqd*S�,��\� �h����)���)Zt��
R�I<֎�18�GT�o*k��gZ�"�{�VA���ך��c(��jhߤ��fٟ­Bz�)z#�R���(O>W�D�-���]�"���س�j��ggڌǬ]1ߺO��@V�Fӳ�/���q�����|���;��2J�W�����+8IR؁-�b���L$�\!�u�$�1uuh��~��)��U��E%oq�"哵v�#QMi9X�|�L�6�_���_"����:u�݅�c-�ex?ތ� �Iu�*�>� ,��c2&g{��{Z�rujk-���۹鸎�F��6�Ė���'����a�ؾӨ��=����))Ϝ��B�巸�fP�*����(9�	c�o����+������d�㕁-����o�ا���ף>+G���& �J�['q�m!o��`��輡Ej�
�`u���av��֛�>A��l���?+z��ىh����}l�$��}M��"Unx<��i͆�5 H��Ѝ�׉{]}�����w"˃q�Pea�h��h��?�&~� �D_�@�ø/ h�u�)�;��P�;�/�`W�ˆ��$�Qi���WE}�٣?��G�+��s�c.�-E�m��q� `�Z���T.*i�����VI7p7�e���瞑��<?��k�CC�O��*��t����i�Tp���E�/Siq�di��E/c�̂&�	���F3.�w�!�ΈnD���1����zI�;�3��q]u�yY�ݹ�Pw^r5�$c����U�i��U�O�i���?���j=y�����~���xF�pR�zSb(�ѿL%�E||�D�&�Xo�W���=��y�\n�7geg�D����}0IώW��|�i9L]-L�<�{x���g2�*X�n>���7����݈�>V�����(�1����ͼ�C���@�=>1x/DK��'^��Fj���MuA��ȿ�l���C��?�~^yN�M����L�{��=q!�0��,T�I6Ԯ}y��(�G��zc���7�o�Wl�z�Z�w�fi��К#���BSP��2L�(���Ks��I�~���6��F�/1�%��&��icv�������[g���=�Z�x���Nϛ!�JM݌Mov�	.������Yj��t��D{v�zFTz馓���n����1YD�ҩ���ċ<��`�'xDV�Tc#�^e��l��(�M��sR�{�m�L��ѹ-�k�wƇ����~O����;��?�ނ����`��`���4�]w�	o*��w�Z2t�J��x���5��~^�iS�@�*����1B���| ����1]J78����q�i]��Yò2k�LH��7�/����X OK!)�We�s������%�Uv:Lbj:x�T? )�2=F��l���04o*�ׁ�A
$�^�ה"�u�ML۴�K��2��������prG��#���P�
Ja��%�z�g˫T��r6۸�ZN�����biU��߈G��J9%QT��q72���@86���W���b�Iq4ۆ�DX����u.75uG��������*C���4�>�1۲;�<P�#n���Զ�#V��T�폒����^3� ߩ7�#�X̢Wj�O�I\���6���o���Cd h������� ��R$5���T���?���ݛ@�D��b�e�u��ۿ}pz��{oR��Fr��6f��M_;jJ3�M�Y_)RGj��43V+u�m���z8hgq�k@�^�{D�p�O-�U�۴�g����R���c�����
�F�فL�AC.�dH�C˗B�6Ӂ��:]��ً�	�#���Q�r6oh��B@y�h�u��w�f�8����\/lT�)3x��	G c3T��*(,F<�[���'`���QLyM?��/`���!<х�A��y�^�RCot���\Ϲ�1�:y��L��G�@�~ܻ����݁�.F�xo��P��RY��g���I���C�"��d�`C/����3&w3���W6����i���ŏ�gΒ�O't0�(��H�7���{hp���A5laue
tn|`�0���x��C�����{O�B�6<P�����k�pz:�3��Y��UBBi	R�qZF����i�c�_��fY"/[]��P]^Y�6��+�@6J���@�,9�!�%)=�$!��ՙ� �j	��ZV=��[�:�7D��2@XI5J7�AꙞvV�*F�P�M?P��g!�C�ڮ�ːH�86B�o�iFl�������N�������D�ԹJ���(����Ip�i�+��3^F�I'A��K$6@Ҥh�ho�D���O�H4H�G��}\�EQ����u��|����iU���D���w��G}V䓁a�f��5�q:��� ��\��OK> ������܈y��BA[�5��P���<�	J�s��rdb+^�Y��e)���R�Ch�%j���1����4���D�i���I�a�Q��oZ�"E��F ����l��{��ѾY�T Co=�o�V��U��B�t/��n�sg��������@��o�jC-ޣk���笧���4�Z�Y"�l��!y�9�:���F��a�[Ǯ��/���f����}���28�����Yh��f|�&�,Xo��:pIq]��1d5�*���j��s�B����wwXg!����(��6`Фںb��~�2���Iu3��h� z����,ЫJ��>3q�+� ��JAi#���e�mr���I���ҳ9�l�%���K/e�Z'tj��fU��>�-�VP��)q9<�e�����T��3ǅv�z�8�Vyh�")��o�V����ρI��v,;P��d.�V8�J��8���d�}xF^5�'���E��ɻ���I(J�+��'O�T�DD,�"^�r�ň ���x�o"�f?߁Zf��a�8*{��=�R�)p®���$�����pB�o�&,Q@�",b�r���cL?��{�Pb\��y��GoXID�T����n�\���.�C~�rCs9��*E�}�����
��-�Hצ���>w��(H�l+0X:����v�a�*r�V:��f�/q�����>��$�U�tY�)̭�	޻���F+�^=%P#vA�[R���ޝ�����N��Qԕ�sms����PN�/}���kh��7���7����ɶ@_Z�v�A���n� �`i�H�����[�"N� �J�F��4\�jı�t�t�����M��nE��H�S,�<3.!�Gb�\C�0e��kBO}��(;~�k�Wf#i�Z��7�|pA�"MZڒ���R��.�	J���z�g�e/Å���l�v=��$v����(�6Eg�����u�H��;��H
���!ȼ���f�*5+��JaـN�����Vw�^G�N�Ȣ�W����U�7r���	�N�@�k����jM��2����FW#���0`qƄ++�v=DG*d�F�,8��O7fC�(A�U��C�1O�7^�G<��~��>�s�>V3���w��j���g?(�
�d��еЯ��bA19H�A���% �|��a���4�o�L\Uoǈ��3W0��(�f�����^@��TpC�Lͻ`z-��\T�!<����{_6�-Ta�|�ꧽRS<�0.yf������^U�����OXQ��o\����j�������(oʞC�a6�า_>z�*M���>�,�B�q�7���a�\��O'�&Ӕ^�p��e^l�v%?���=���6�9�z2M�0&�#@O^5���_���2�7�1�,Vx���9x1q��4�mEH���}*� w*/5���x�^۰�����Cb0J�}��a��skl��&|��SN�E^.o�@Na,Z"��q@	d����w:��P��<B^Ʒ7v��"<�$������e�����)��i X���XR�:xV��g~8d:c��0ܜ(�<�̝��^o���5��޵q�ծ!��AV�l��k��*�����i|/�əb��߃D��q'�&�������������F~8�"{\�U��L �ȍαv�t��F��36��v�K�OH����7��I�{d"�5�Z���#�CL��ːB�{���PGB���Ex�QZ��m.�d/�G����s��B�dV����"�{r=Ckɪ@�]kKٍ�r�[��$��iI�?����,:&�Ɠ�����γܫr�*"������u������Vn���XI�d��-��4+�g-��i׷)�����`����8Z�?	�����n���֧�C}���=9��aҎY/m��^�-퐹��،eë��Ւ�ͭ]���P��h��G ���DjN�:����Pz�V���{w�E������w'�K�n����)���qH��ҳ��WB�'"��@6���z��Tezᷨ��R�5J_:γꜼ؆T��_iv!�z��\"��K~�TX�qȅ͏�or{�N�g��Av���l��h8MК�aa�G�^I�1_�9�k�������a�9���◗�%��U�.�X�ĳ��;yP�N�e��n��8V�/._G��Yև./+�����G�_:�>HV�DM��#WŌ�����@Y�QF���s�@��f��-�����p�!Ĥ:,@k�32<�rd�.p�՗(�>�+=��U���q����R���m����� �cu�|e�^�����y��ZoI�u�fHZ�L������M-���5r�դ1�W�/����d��#��s9"�3����Bڡ��F���8�&��#��~Xؿ�?��Z�nAh��#S�Vv�9_ק�f)�֏r�`!���.@\`���7�v0���p͎�7<��m���e�}a���}�&�\#�J&�lk��7��:	���%dl=��,�����aJ2�H�����n�l{fUQ+�g���`�Ca�K�򼰡��
���k�����k�
�h�@0߽�)�f9I@Q�D��7#p>P��(2!
uS'	+��?)�깅�6�bR�ǹ�TzR9����9�PX�}��[��=ׯ��e�+P��V��'WK����G��Ě(O�]�z��a���l�����Uܗ�b\�޺zy�6s��f�#QZ!1�
t��I԰��z�c��`g7��h!I�Sf/���_N�b6.�p���<4����u=��Q�͚6�� w;��]E狫�y\���u�ʷ ;
��-��{�Ƈ�f��}>T��`,�������ɶ�v7�
rZ������#���~�t�ǯ����Ts��R:hjA� �U-�E�c�d7���ḭ#�-\-��Lo����<���Ck����!�H¡^<
�����O(�A#b��"5�;��dH/p~�`��@�T�>��IQxt5��%;_��Y�v����p���~��5_xM*��6:)�p�/�QT
����ɗ�Q"�8� ƛ9*��~>Xv:�r��N�R���� 
5���a��{tT������q	�;t�lWñjv� 	�D�]�>2eƗ9��=������c��]�G�� ����J�Bבm����6ʓb��,�;9tS����kS
�Y������G(�4���:�ӓ�7�pYP�"c��E1�Ǯ9�x"��H��Q�ǈ�*^R}f�HV�Ɵ��=K�g����b����u˿�0��_�4��l�Ol���^v�W�Nsii�;�AO˒�}��ߏ�R�N�W�|0�͉�>�s5���6�R����ԟ3x��	Z~�6�wz
K�Cm��K�6�e;US�{K�ru�
XxTZ����iQ�x������4��焢ы��]7ƍ��s�JUyhŸ�$��u���
WXR'�+�"݇�U����z�O/�=�v����&�Uۥ�^H��5���\/����r��N�l�U�bU�g��-|�`��9��0`DX��������>x��O���=8���dh+H�BX��̻�1��H��5����v6g�,P���7X��e-��<�k��bӬV{"����x�T���!�jN�� �e/��\�r��XTY�h����td���']+Pm���R��3B+��
0�=��U)\08��t��/�,�3���߱C�>�Aܛ4�,���+�2��"�^W+ǁ0�8|l���d8�E�	�Q�=�}�.pK�5N�l�jF]��b~yK�f̎٧���bR��%/ĮD�J4]����O�*�� q�"L=�@L��N��3��4�}�ށƹQ�dϞ&Usn�c� �4qę^3��І��e�^�&��\�h=��~���G���#��D�(�ςi�.�lF�g��m�`O[��W���#7<˿dY�X���Z�M���F�`}
\�q�CYX8��aY4s���o,��^� 0#p���-���M�C��\�_�i��.��_.i�A
�)d���Щ�ٵ=+�����vE "�ฑ���4�?ɣQ�?zPȁ��[w������x�Б[T3��3|�q�f]�d��5��_`�~�ۛ�z�3��A3�c~�I`�a��֎@��,w���ђ�~�~#�5�~�:⊻�t��J�z�`u�|j�iI�J6���{�~�������cģ Mt�b��j����l_Cv�x��H���E�zn{�۰�.��,���j*"XNL��:��H<�Wfd�y�G^�!�.�u�1��t��fi����`�1���m���il��`X���La(	��Q�/U�K�x�}�*;fql�{�G�f��*������L�T�T'n�]�-��@�
��ӻiR�&r�[!mV@!�������_V���ے����j&�>�0p��t��R�%pb��:�A1�Z�l� LpM�i	��#��?)j��Z��ӡ����RK�j;s��?+z������K�'���@�h�R2p���L�n�+�f���ߡsy�+#"  �������̃id�C4�Z�8t�6�ğ�|Y>��%&|�A$����hQ�� *�O�x��]�D��&]��O�rڂRq�ol�q	��$�O�ZaO �ZPk���3"�#F9���V�SmQ�`j�ty�uUT1A��	)l	9�l&V��{C[l�S9Tw�Rl��s�X�5�w�^�a�ex��u``VL\8n�8���W۞�d��'�	}�����4���.��B���5�G���0�Q��S䘸�b.���`_���ՠx�TϮ���;��Y߱��B����J�^�Ǌl�	R���Klft�B{-
�ė(�h'�e.�Y'{\ة�uz��nޭ�3Z�xC�q�@���dd v��v_�i=��^<&�pz�<o]��cq���������^7f�qgsJ�P���lS�ҵN[��z����c�\������T%�\�O�f*���Q�>�7�a<�B@�}ЫWD�E��}��}����>ʟ����]��l�*A�{���B�����Z�$�Ҍ���DF}>5�U�=f9_D�� "ҫ����ߞT�RԱ?8wz���?��8�7a��E�n������eAa�RR��& PR.�%Vi��$s-4>JX�m$���۰���6�}��Y��ًfU3Mb9���|�m0]����CD�m+��6��W�a:f�0)."Q�"4[{��ʰd�F�h9V/�J<��O����H׈�������3�}�ؑ`�{c�[�Y��~���:p�l�d����O��dk�����C��ጝ��a�U�#[z�=]�&�9�i�X��0n�uLWan#���F�ݬ9�����hc�U�;#�+�W���goӗ�D?�h�>����r.Y)�od�N�C��*L�@< �(��|J�&�S,�jr��y�D�9��x�����3l���o�}Ob!fq�����_:��A�,> �|9ĤNN3.�q +��eZ�8����9i����q��b���>`�\݊�l������`�0*6�!W�Q��un�(]�w���踆����N��@�d�ބ�.��w�����i2�"L�G���V"7mX�Ke�+��������,�>�"��k��0�tZ3�����- ٥�}�Ҥ��x���n���1�;�ͷ��Jl�W�d}:R���ĥ5��ƥA|�_�6�ǋkt�����G�sT6�Al3�H�b�:s
��	��h�������d`Q�Q`�1��l{�{!�1p�3E8��0G��a�WDmSk���-~���<��=��g��ʥ��<0�#�2X�46|�.M"���t	��`���K\6�����E������"^�#�U��g�2�HH�!�cbE��5>�T�3�Ҝ;,!8����N�Tl��*��@���~M�9Z�x�u�����N3��mN�H�I���U_d�$M�R�>"R�`��5����>9�D(A��7���V
u��	Ns_+߆�*�&���AMĮ*�7Jv�̌��j���OU��a��~
��f ��� %���ϬBT���(�FM�j�RH�1��C(�Ed]:"��i�{�7����,���$�w�b�[��`�@��(�HJe�xJVZ��%,>��Ot~|æ��눂�C��~��7��_��x��X�^��-��s^je�ʟ��OO�|6� ����/m��R,eoT�;,n��h	�����(��Ђ����QˎAr4Z^
^f����lL`CSϺF��-a�rc�"�Y���ש�&Pp��?�x�\�5n�gZ�P�h���Q
���v�����9�(�������Q�&�T�i���U4VѺL��5�~��,z��1X�Ђo��kC�Fo�뽈D,�/�IV¼M�G����~������Rt���yH��{eAă�Ad�]ƢM�8u 'P���k�3�����^���k�)M�U\/��23��:"��Y޻�E��N/�Ez�*����P��y�x:�PL-B��}~WD&sf,Z _����cgVs�J� �w����^�.%�4�ڒ%h($�ד��ڜKc��M͵KX=d�;��� NE<�T2$,���i�F ew*�����T�k�n�'������]"g�_���xx���|3`{9�J4�^x�x=cB��c.�̞��z�;�O]Y�2����M��'{wC��\_9���i�r��k���� .̜�?)�lBj32ԋQ͔z�X0��Ʉv��\�(��&W^���	��|�H��M. ����� J�����p�q5b��������B70�Ejg�*}��<�	t��"W�K�5��K�M��N�+i��Tf�%�dfBR�f�L�2A���d�����c<K���0���b5��?�i�Aw��Ch�n:�4���/�1;��s@,~5R�����Epv�� P\(?^jc��RGi[g��|�]�S2��R�����ձ��S����!"�0��gګ�!�p@��k�g�'`� _�X��t/m�d(f����x�:V&U��d���X��z�����7=ؘ�Y�U��x`e����|��`sr����z$�_� ?�{}�A�����g�]��6�����\�gP	�S�V����˛5S�a��z!��vO�w���c���rAxi�3O�ڿӎ*`�c)ׯ �Gk���M�d��p�$�ږU(�SI*��P�`Z��	�ɤ=��ܴ�0�R�\X 8�s��NF
S;a"�5�M��IL['BX�ؒ}���n�f��x��+���&I�Jx�^��(�>ǔ fC+	������+X����k��Q*�E��˷B˚(`�iԕkB2̭��D��7.Sv-�]�79�6�1	z���(\����~AW~I���雞	K r��Bg��r54��LI�7�r
�.��_�;:';�6�J2p!Q�.��0�uDQ�z��� ���leo����hǫ#G4b�gC>	��m��:�R㟁&ZS_y7xIݝr���'h�:O�E��*��� �T���DG�g/J�����e��qr1��t)([oկ9ny�^��qڢ�v �̮��MXVM����ӷ�&��^ѣ��M�${+�+O�-lm9���BC|"	r+��6����VH��F����	����\�[�V�8�DkW�_�;<;��d�T�j#��]yTj=17����p*1G}�@s\l.K46���K���	h�[s(��2u��N
h>��yN�׹I�J;��� %��yL� i$-nT#+�zaJ	��������EMOa1�:ϵ��fdN�u�/:�S�Q�Ҙc[ه���?�8x'�\���e5�o�Go�-[j��(++KeE���Q4Q�/����P>��>K���.�P2׏��J�Q3�g�Z�����2�)a��.{�\� ��������%��w���FԘew��-{�+�\#�%����hO�� �G�"gi��e5rK�{�9��,�����������U<�2g�m_�V:.r�٧�T}$iX��24���[�ą'��|�c�s:�.'S(���D���ǻ��+����K��ս�MLwaYWu��#�
"y
����F0|�����uy��$eN=����4!��f"�XF�<o�;t��� �ɵ�*Lx���!��:�5�G$��F���e|;�]FU ,��_5�S��rJ�ns��Sӑ�����$큒U\�͠W��K��D�i���Y�LG���΁�v�X�֢^����2���{'M��8d��C��}R`�᫁KÞ&��� e]l'D�:^��=�Fr�a;æC���)߽/�|Dd�|/�����
����pK��Vn-'N�eX$�a�(��"�x
�JTU�\U�P<�ʦ���)TE�4��"q��m��{��%o/@�0'.h�R�K��R�����܀�zҫ�%�K'���VlzwY��x�b�o�5���IZ4%!ّ�-_({P��F���e\� �xty&����8+im3�b��������g�Ҍ�H��s�� o�6]]����I8�f���"lb,�G��O�J�n�t�ݭ�'<�8�Ԙ�3����b��}֟�7����^�i�x�!wt�z���َ�J��*
\�G��(� �+;��JD�PNMr�ϐ��#��p��Ju�NՒ�<Pqr���].��b�d���f���95R�hg�!��Nd_mւ����	s�7o�@1X���u���S���]�e����	�<�@�C�$(O3�o�ڞ{2;U���t�ƙ̱>C|N��OV��V�jB�v�R��l[��1_̋��N!0e��i��ۑ|����6Ǿ���_o�b�6Հ��\�(�ƎUo(Z��0��|�/H[>C.���˷X؟���Ì�+��S�
�K0��N�F����(.�u.�ZH绡sG��O��/�菟,�қ�Y���
�y��� �]c��GsڰLjm�z@G��:yD�c+@�F��4��M*[A��M�q���l����c��t�w�L�2���);*�1��\xc����Y�v@�2�<Ȍ�l���)6iܭ�*�脧eǼ����]��g�EN���U{���(s�i������޳�+ɶ�.�{/��=���| 5���3�oN��A��i�z�P��_@08�d�vc&�J���3|��R��uZ����C��P��aO�,P/�ai��=�Ǿw�/_��᫸����K"rˏZ{�n}�X����/�I�{U&@�f��`�4^t>��\ֈ�~`��̤+�&|��6&��6�{/�DV{;� �𗇴����PNYc�E���i�ǧ�����(�$?��S��;�g�i�*|v�ۦ"���<��-WO'�!cWp�2�bTVof���ul��mf{�<�'�0*s�$b�l4Ie:w�V��&
��JI�|<8�����R*/,�s���6��w��h�s�\���o�Ѓ�oɝ��x���b��t���f�YV��-^fi���a'6�q��'�R$��r�-y�=���vm���vP5x�����"�5�_��(��`	q���Vf9�Z�q���S��I���]g�l"� ��_�<9��J�)��o��d�����U��.�R��Nqa�'e�NY"^��ю�|�%��v�^��!]_ӎ*�֧�z�5�Ja����s|����⍊h�{���"*c>Y�x�u �EMQ���3V�I����h^��N1(�S*f^N�iI����g�.��s�����R�LY� �G��'�oS�<V���R8�p���tI9y8Ǡ7]������e]��"t��	o9�~{�J%���;����j3t��ɓB���.�)��ѧo����CA|�<wI�M	���n�#��G��LX�ޯ�����ga�4�;�d]��З��M(]�VԢ�NN^��f�ЩS5UZ�O�.��:���Sƺ�Yp1�j��&���p�qi��rI��e�:�� ﱋ{q�U�;�DL1:Z)�V��i=���ڗ�<��,�(g�ijmֆf�2��'�i���P�q��e�d��ڕ���O[kq˴��H3P9[+�r�T�"[�\�W�v�[ �}p��{���?R�v ����=K�,aԝ "�����#!n�ٗ�cK.,;r�)p�P�GI���ь��������3$���N8Y'�F|A�@;X���D{����|�=8-"���+��0 ��ge0��I*� �V
r	f�%�/A_J�����Q���5�1N�qX�T�
��g(rX�%��Ϣ� 	����.��y+!���]�����r�r��u��a�IIq�(���}4HT1^���F�lm����/�1� C#��u�к�.�vXxn�>��?�	Y�?��l~��`�H�3M�e���������bn�Ylu��&c��np��N�g_��ba�U:��N���+߹�m�������ک�V9ҷ�ɘh��������Ni�Ŗ�~HU�ՃE��˱�Y�
��h�h��	9\Jg�)F�	�P��y���*�#!>[RQ.���,Gd��,���oP��[�Z7١�f��/M(�˭[9�4 ��c:����"��d�`jU`�рDu���Io7y|�Z��i
���0Q�C7�/(��iG	�G����F?ҡ��tG;͇@1�l/NH�'E��ٕ��٨H�e���K�B@��$2$;}S���X���������>=��:�e���#R��Y�N����b�u������$�+���@pLr=���޼�g���Bb�+��֖���g��;V���)����������w�IK�.�M��uR��ۧ��h��$��ϑ�O�9���Z�"~���H���3�z�٪\�/n ap�C����.�lx�U�,�$	�\�H�C��uJ���)�O�@x+�A�!x+]G|��zK�#}rG�zcF�}AA+��r�l�tRj�?s8�m��f�����>O?�^=���H����q��$�߅�C=tK�'_�D���U��,�{�m>�`�I��U�Zc�<-��:н]17]�8I �6W�Pgj>G-J:'�Xh��ט J)��}�6�X�^|5Nx�R�]u���x���)O���Va�(R�Z���9��Yo/��#��B�F#���Mt��"�l���Գ׊a���x
'�/�����V3Ŋ7���G����F3��mC"I��a��}�ď���F���f���ޝl�$4�&�i��A Q�,�K�-gp�v�wL�?�t�k�5N<���ͪ1�Q�ˊ[�1�� ��c�Z�e�������Y�Gz��H�x)����	�m3I�'RD��]���5a�����`�<�r��.^Ia�j��}���k�4���S(bIa�R,Y�1����%]��7�06 �&�1���m��;<�Q�e��G�=�͸��3����l��3T]}8�栮��R�t<&rG�-�op���Վ�z�g~H��ln����g��w��\��^	�$���B�ĦI���ǑF���ѓ~�W���f\v���0��M��h>MC��˸*�\6��3̭��Ťk�4�%�I
9��5��H�jk��&�wE٩���ggpm >�N��S���M }5�L�-��!�/S^g*lT�6���fRi\�D��ij���8�,!��*��t�����ޡ���$٢��<� s��Y���ٸk����2�(b>�����t!D�|\M(���l/�/R�=ִn>o�:W�,�ED�x��f�P�4P2	�#���6B.�����aR�]:?�RA�\l{�_���l�Gz�b�n`�W�f�d'�����'	N?��)����+�j�~��Rg���<���ER�e�h,l&�??�O�jD�3v����=`0�j������`�ڌi��f�"�"qt�^��bK%a�H7a��iw':
�P�Y����)HPl����Gf����h�U� b�������n�j���D���y��sK��-���;¨@7
q�aD5��=�=4z~�a��g�Z�6����;���_5I������S����D�D�{�P�d�H;��
�Xsa"OI֑о��ʌ�W�$��<u�醆)}{����RR�U;���D�Jx�:�|a��E9S�W�R4
?��h
4;���_-�u������z���8͙x��%��6Xys9�5z6�[��©Ĝp���k�o2G
���v,X����<A�R�`Ɩ���J��5^>5f�b�>�	����Ɲ=ډbP�Gޱ̹h��/��R��E���C��8Y7�Z�.`��Qu��n�F##��oAF�F�y�§������m���VN�[���R6���5���n�Z��rJ6U<r�.��y0���a���4��V�O��$*��H�\l�`�O���(f@3��3c���O�Oh7�A�@�+\�l�X.E拔Z��oI�q(��$���Ӷ��GT
mz��K�z��Om=��+���/��Ѣ�ZdJf����Y�o�CXْ:�A��b��1eh�N��}��:�%��[av\Ն�e<���k�%E��_c�J��5J2����!9��l���]7n'f��Nψ�S�9�) h(� ����~Z�'�ˌ-dc�B���g·����o�Х���y�UoZ���QI��M$̗��u�%�n�}>7Y��Fm �;Y�m��z'��ye�8.�u2����[U�%#WQ\��H�ݬ�F�������:c6X
�~Xv����&B�d��ڀ�Q�miJ�M\�I�FzV��!�&�CT���[�� "��� P�j�<�e����	q��j-��#���{ ����L%�	�;�}͈�G��51��<�XS��4��#�	���4�bx��x��Gt1d����T72�t�S�L�E��a��1��RI�(����T1,�,XyĤ��x�Ru�`��f�UJ&mve3C�)�Z�Q�<�a�~���7^�t�ob����wdqt�ݐ$dz[�,͐�E���t9Ԕ��!�v�̰���B%��K�R�9�19�֠������-N�3���Q���7���,��B��i��o����S���9�	���q*J#�\YB4y�s�2�Y����E�j(�Ɇ�M�9e?�%S"aݾ���]5~�_�"m�s�?3��	�>ү��nMҏ!��������VF'�� �Vy��]��x#��O})�*�1��N���^0�p_�1{� WX�V���	.��+�Pȣ��z_�#���;g�{�&i�=x�`�f��jc(�������L�DƁ�6a����S��F�Y�+~(�y�{��D�9=˿Y�τ���2n�+ݴ#�v���n0"09�(��y�X��/qi #.��=,X�;ti��k	�pS�zҒGg��䚐?�q[�n�j��z��	�Z����E���b�Z4��T/_c��t�+��8m��2�wo�U��J8� �j����ı�>P���{��s�jH�D/��+`�(+�I3��,[�A��kk�{��)�n�u5�}�a׀�j}�UYd~x%ͣ��R��Z�W��׏�ء�gҜB�$'��W*�-؆�]���y�k����c��c��q� ����շ"�p���.��C� �i��En�����{�懿�!5����I�F�X�ّ$�0�t�X� e���O���Te԰?^5%�����D7G��d�i��2�\lR��>�c�^�T�!ػ���
P4�prr���#*);�ث0)��OR�w4��)��,��V�mƆ����)�%�d4(�%P���fH���>#���g�_�pOb�*�b�ɳ����kZf�����9�%g¹n*�W���p�)t�k^I��Fq�RFZg��xQb�#=��BE����|y�N��?�ٽ�vRQfi;E�nV��t��ˠ�]8���Ӟ�+�<���/��P����W9����	{W&,�2�\��V@�^غ�b���6�V�����^����P����X�o^M����F��4a�K^�O�����h9�c�J;��_(6>�� ��b�#���j�k�	��I����Ø�����xU՜�YKQ[�yT�,8h�Oa3<L�d��n�0��:F���x�Ҹ���O��[�pV�Iwm|�z'śGI�d�xp:��*��PXs�W��y}ׅ�l(esx}�8���q&1XM�Y���g��&��`�܌��#��<ّ�6p��~�`e� ��,��!�I!��ߤݞ�{���`��ҢI5��sQ+ !��QaFݿ�*��pp��DȨ��Z[�'�"k#}D�5<0�O��ac�-�z��#-�L�:����ȟLq���&���R�Nqj����r���=�	Q�^�i��K�v�jO����~����v�p|������W����<�.��>�s� ����98Z��R�C(sl��3�:LF�����8�=ڒS�y2򏚧��X+{9P07"�2}#��+ۻ��\Y�I��h��V�!U%�-nde��"2J�ʠIϊD��K��T�+3%ꮞ\�/aQ�[�Z�����=����% �>�k��Ҟ�4L�N��KXem�]��rSɡ�uc�,3��E2#*V-bS����$LE8����Z�O<N��ɭ;t��7�x'�{����9���� a86{�{��x}3/�T5PF5ͩ��2��Ϊq M����0�I�"I?�̉v2J���AC�\pB���sc~��I!׾"e�r�"6h�VU"^X�`�(s!R����6�&�~GA��@��U ?�@'H�>�p!R�e�u�6r�<M��1ͨO���|����_r͈�,�z��qB7�d��!�#+PS�%���Od�=�_�v's$�<�ٯhv�AB�iR�7��\��]�Z���f7�hR{C���ZfB�-P���x�����5_��i����r�&M�B�R�p�[�����̪�H*$��)D�8Y~0	�ν�8'��i.!�۟5�.�
iq=��Eӵԕ����8.|����ߴ<\Y��GX}N���ۧZh�)��'���8�s����M+�{��敼�a����%�Cx��;�=\?*{l��5���MW*�S~�{a�zmެKb�k�u^U(!I !]�>���!�B���-���������q�x�f㕏�x�H٘u.����c��1���Oz���"���V	(��_n��%M�p+-���d��� �ﺴ�O�kx�'��p~5>��Z]����[na+вu�Z�����J�av4w�P��ݎ�R뽩����%r�)�G+{��RP�hb������entXXF{�E]��@ž��V={�ɚx]R�mp�E-��w�������bq�a8�c��%n���L��m���r5.z�5!�C�� m�8���=��}��5�q�QVע�s����磵���L�YO��"����%8�%�	1���ʂA�))C�sՂ���A�!@��\�X�x|�/A�bN����,�
��] �JzC����)˾SE/���Y�H�/Q�c�niɦ�k�ֽ3?*+( �skո�ͺ�܉,���WEG�;�T�z=H�Q;[�3���0%����6�`9�~e�D�Tĉ��%��u�
8KN�|�LXnE@�����}�d������1��	��=z��_(#<qAn�2�(���g���h�M J|#�O5GZKY���V2�Z��f�!�[Y�<IA�7[<���|���CE�T�ʣK�_K�^�{CU�`�H������
����q2{FSwK�>[%�_!��f:�g�G���G�K��ST�el���⨠�rǻe�k��a���u�(E�&.KsC�����ۦŹ�i��
M	-�R�|ZvP�����+0��L	���sx˿�l�f�B�Ș���U�1!"��5_��,��徥�ӦÈxR�:�(IOB�0����Jyz#N�����S�u�lS1
1��۩ƍ���Lq�m�N~����~}�����<C����䈗��P)I�s������r�B��=�X1�����<��l���yC��>�pW�(<�,ï���"g��T*Բ�M��)c�Uu| ��70�I5e��91f�"�Z�jc���
�84��זS�nF��NV��-�L��R�ok�-:v�5�(�[4��Nf�в�BN?� dZO׭� '+Çw9%s5����l��i��qCZ�a��U�?�M)�u�<��8�{�	>�;���8C)��v/T�����X�zғ�nN@��t9�t�,]�����K��s����%���d`�':�L���Ǿ~UV/�Д>�����I�8��R�u?�U5Ta�'0��a3w�^a�/�A؊Q�]�o��Vs��ⶠ���{�R�� ������&³��4e���_oDo��V�U?X�Е��,*1>߸w/@A`n;���km" �:S�3���D�ΫKI*.��\���|��QV[��+J�v "��h�L��ݽp�G�0RR�;�[�n]X}��m�:�]Ȗ6��}�l��9� ��p�����*����$��~j�N<��5Q;ƛ n�����(��
���
#����1���ҟ=���/����`���q�]����D;A��l��8w���W՗��e��mD��l����9�����Q{�hn�k~�T�ꜮH�lG�������㝇�i��OH���"R[ʤ���0�݇ց� H�Ip���`���')8,�K1����Ĺ�y{M���ǽþ��R3��D����Wc����mE�^*!�dv�k��y�ON`c��iU� �>f%a�(YM߄�i ~T��yH��#7˔��dp�\ ���hVr.6�}�K�oRV��o�1g�#�A�-���vY�}@z������}`�_����5p}@�^WE}I5�쮑X�ڹ�ع#WJ�k�~�0��'�b��mڧC|@|toӍ��C^oj�XuR!�M��A�-"�rCA�&y7�١@�G[� �8����ȜS.���	P���zT!+���}��d��1ҕ!*������`+��2|���P�nn�\��\\Tl�C�|~�n�3n���v9���m��" *�		�;��c�ۼ/�NL���)%��ɷg谒wF�P��u��G�	<k�,cձ�T��F��P����sQ�PE�8���n[�^��pke��Ř$��D>�p �:R��CѝQU8�T �:�N��1�j�,`&���s�Ի.{ ?n#CV3*^y��~9]&��q��h�}����[�q�"���J�M��N��fS�z?�Xg�2�ZZ�,�k���oш�pnD
�CMQ��1�|>CP^Ij�O~*�]���E�P<ZA�5�[�Jc�fU��l�P�T�E[{���v���3\���C���䗁+I��36��&��d�9��l�A C�l���WP}�*�^p�TUm�dǚ~����a��$L��ul���0|�\�ʡ�f�;��n�`�Xl�S� b��%j�O�+nB�я�HUτ����:ۘe�^4�� RO-=d4:��D��y�gJ�	�J!NW:�!��}_��
�ω�7�+,8
�0�)b�s�^�dJ��}�z�_���8�VJ�	���5��V6ę�k�I�?���/�Ht<+�t��!onQ]�M�N�J�]���CX0Bu�A]���g����l��֨~����I�e�ޙC6n]+)��+W�`6H�RyY���A+�%ё]�n��׍���+�,���U���8�4P<8��2?U��֫��	5O����{���lя4@(2`�O#I�G6�1���	��m��.JE(뾥�^���˸��2?(m�:dH��Jk�%��Io��=�h���z}D'DHD��4�f7ݘ)�/����}7ƛ�o��qf�����?�ac6��z׉Oí��(8p@����9��˂^n�n��:C�ȭ���98٪�qa��B�:�:T��nۥ:t�)��沄6ʎ��hh73�y�xQ�o˫b�5Ѡ��0��;ݼ��1d)��@#!��z�A��n�//����W�̭'B���s	��͝�m��d^���f����6���+���b��-}!�`L�?����%x�vV�K��Dg�T6�Qa�u��Ȫ��9h� 3	dbzP�t�����6�-E�l��f.e >�k�����=%uv@j��+�����OꜥE�@4�z���W����h(��4QN�����2$jb/������H����*�rY��Q#L x_ʪߴ��p���v�[��4��d%�z<?/R6�����C����b����_�sT���s�o0`<8�V���Q��! ˓͟���a�ؽ9iu���0��8V���Ӛ<�*P�Hi����{��LW$�]i0�A9� *q�����%��uqI1���Ƨ���p��J���u��7�6&�^�Ⱦ��_Lx
�G^���1��C��� O�i<���I<�E����ϣ���P���lf�ӱ祟���A���M-����t��/P���>���Ui�Xu�5l�0YFQ7��P۝���Wp��-��_g�����k?Ş��Zʌ�#�T��A��vG7SkV�y]�7�p��j1��5���ݟtm�D��gXK���l#��Ӻ�����q����x�,����T2h�C��n)N��.��,R ����+F����p��Cf���8W�F�D���%�3٭(c]��h�)��X�â$%�ߝ��`V<M�MQ�h��.���s9���>��n�����?-i$t)��<o�x��ig�^UQ�E�8��˴K����@�cU�w�1��O��׻�>@�������Q���4��_�k�H<#F���/%�:�u&:�Fn�Wqx���$w~<T���w�Ғ8z5Q?n��*�$�Y(B�Ht�XzǺ��V�m"R����Sغƙh�C���)�<��6�[�߷Xt��6���D]H���憤�^����*Q�ݸ����oEfza��|+=���=9d��ZH,�ސjjZ/iX5Ϸj�$�}���� �R0��/j�烈{ڈ��� �R�y_��NTU���!f���
�H�����OQ�I�i�߷}��49��!�(-9�y���t>Zz���6���N��N
����Drي��B��׺�7���AWW������'b3�erW�����:[���rd� Z-8	�I��H�w�d[�P�$��c�jO����s��;h� �E�m�K�L��	�� Nr�
~�эb+��+d��MV�U�Bթ9��/����iG>8[j(V�	ݏ�t��)N�f������T-�D;�����"E�4m�7*0���:W������3�q9r�~�}έ��c���	���s��0� ����U�l� �֫�̫�O?�;��{ �U�Pm22�>��(�3"/U�w�FѲn�VnW
���q���ީH��~��Y�^��3Zj�9;����8#��^�� ��#�.s
�.�c�W�O���OL�� '�G� ���j>WdaJ$�;2�n/EY�lOo�2��wT�X�	`�V��_;�M�k2n)�1�'Эl�V�G&�Nϐ��/���R���c܅�X�)�ؚL��O�m����jF�}���t�3�+�d�Z5G��n2^��=Y�s���V����xG�[�w�HH�	��+X@�W�D#vʵJ�ީK�|��	�Y�óO��ZO7+�?�鵺9;˓���,���g}�.7�b��Q\!R��"Xܖ�$��g�F��k�{��z�����l8��"0�"����EM�`,�C$����D%r���4U�LK�[b*D^�����/e�_f$n��V�GS�Ƒw�,y��2���w��}�5Yn�zg�����.�����Y���2u��Z��N��E���f���H$�u�L��?�9�UJ"��p��4��\Qv/U��uӀ&m6��;k��m�C�QN�J�Z5��a�(�J��dϐ��ktT�@�H��@\�@�B4lC,惂�O#���tV%�o4Ї�B�����bt�	�]�|��O��/4�k�����7��]�����vBh��붍p���#�[��a�x0�M�6Z� �8'H�6��$]�uk��.�T����ӕ�qz��s����`N،͋\2�D��ea��*a0Q�p\�գ���nJf��X��,L]N�l�;痡��6
*�c��o���5�>Sw�(�-�r�DP�C�Ipн�2PǎP����fJ���K:��.�CMt�4A�'P��ր�f,�)�N(�f�k��'(����"�W]Ͳ�vZ�f�s̒��2�p`��!�R�a��s���x*�i�݇v׎�Vl д|"��׏u����$��� �K��ȬR>�i��!�����V��ۮ+n��1!������)�;_��{�YnuJ*ŷ��-�"��_�����o�<g8w��:�����g���@$�G�}C��L�*tc��3DG�;VX|��T�~9�!�p�5(�v��S]ma%�H݉����u�p��L��Y�3i�+�5ğ,uh��V��*g�3V���:z�=R	�%�i��z d��8)���d��А&I�T�x9gI�C��9�B[���ư!IN���5T�'p���h%7i�����y��J=jC���m�i,�m���q̟=��b�M3 ���;�9je����(��Ei4��]S%�xhW8�H��;�Z�F��J�Ë��\yxm5TrW�5,C����w3z	���j�� ��:�)�o:Z��A��DI;<gV3z��09�fT/���pM{/	�{�J�&��4d|����s|Z�|�\:��|���|n>� ����`����e�T�EaG
T�X6x��H5B�:���p�h1������A�.}u��atB9{�Qb�(���e�1P�^��P����rI�5�^En_�zzC�N6�6A��,���;�?E�+uw�~�-ж��և_��`m`�����H��]�m,�����(�e��/��͡� �~xt���|�J�";~��VtM|(5����Y� ��ɩ3F����dEc��"���zc�w�<bw� j�h�R�ˉQ"�	Zi��)�i���4B֟b���?>=�͔��^�"����(�Q�v�`J��ށ�{���xp,_7Ԏ=ܮ���T�\��,'McP�zXLu4�5B�����F�&��hh@n)~Ԓl���s���'>��qWӫL��@��=���j��^�?�%�,��-���;�6&�h�PG�¦����x�x m��	z����6��i��Ŕ����(S�:�e�J���~��n�{��j>�KM�1f�=���̦��-Tk�����Lx�=�)z����)UA^���6�pن,	>3GF}���M�_`�O�d5��
]j�˺V=y8a��8��5t�K����Ŋ���@���D�2����cp�Ez��A3Ӷq2;G����1PQp��Q;w��s)��ol0�ۗ�D�I<>OϞ�`�zy�܍H��x< �~vr�\B5r��Hc�����Ue��!��\�U����:z�Ս��W�z���[�����:�T�0H��82n�Rp�?���z~z�Puыc��U��΂V�8��\�4V�4?�ȉM�{�[Ѐ|��.��46�\[�l~=7�&�h��ơ��?�+,o���'ŒP�hW�VĬUs�	���y{� �w���^l�7�矺Ov.�&2TK�bG�L4��>;��5��3���p�xyX;�7z�
 `�]��V�遹��`�T4"�)4��x�_�3�r�b���9|��L&�R���)�U/�ϋ�x�N%�GG�V����Q5��~|��y�wguX��	��iWd�v���U�0�s���} ��v�*�O���NOɜ�%�%���ωZ	9:J����W5s�p�>2y��ny�y��%C�_;2��&��O	��毫z/��>���J���)8�
o3B%�w�qQ�g;����It��лC�)�=Z����h��+�M�4��X�děZ�	 ^\@�>��s��#o�:��7~�ԇ�؆t�Pȋ_�v�>I':���TNM+�� !��pR�ηp~>v��%(��xˈ�k�Hw{v��s�W~i>�VM�C���￭q@���I>Dj���� MY�3�w�
2�^d��������A�J尃].n�8��J�V�V3���c4����D���C�k���e��p�� O`���-n:����oy ��F�)<�w(EY�1A�a�r蜥dH쒋����
�ZИG}-��>�ۄ�)@e6k�s��=b�<�2��)��`C�J�]���y\��Iz�O3E�������w����8=-���a����u��#��<��e����|��Pi�O{��:�<!����:�`����F��8�\�A�׷g���p%X2��$�����N�5�b�`gPk��" ʶHJ�GZ�2/�J���v���T	���x1{��AR����@^�:ty�Ui)��ۭy@��sƆ�&H>|7^��5U�u?!�r��5Qo���Q�䍈�ާ5���0�ҕ���3U�s����p�ɛ��(E6�?�:\IJτϹ��{�
�h����[��i�tw�Xs���h�����P_��q�۱�nܞ��M�Ys3\ =v�.:��Zu��,{���˅�ү�T�ox�'��L��������s[�#�Q7$6�/O"a�#�vK:�^l�O8���i�c�E���_r�H�K�݄N�}��gy��n����>j��4�f�O��0�*��� �E�G���C��E�h����@�����!��gd9����s|��I����j���l�	��I�7��0��7З*����?'�-��	͜�"�ȿ��Z>w�]�Q�#�����ö�Ct��V���A8[����/I��)�Cx�HH�j�e�=VS9A|�3֥ [Y�V����ph��Y3����w-[���'����f��*��^6�"��3m{wء����9���Q���nE@t�\b�GF4� � �;�T�f�&X�Z�[�zk���C�����3p�粣7I�`�&*e_Wޜ0������8�N#��e�Sj౜ÞR&�c7��C�Ӳj�z��JC��㘦��m)�  ���� ��i:��[yEsa��(���@�s�׹�^u�$I0K�^w���u�nӁգ�C��̻}`��Wv�.�/����%���v.4��t����?MU��ו7.�O4����B���d�#� Ｔ��h�z�f�x�1�օh��b���Y${H��j.<�g���"Gل,�LAO�[5�M����"}i�r�
ȲOu���K����3���2�d�����sG�������u
$���Q2�H�Z˕+�ieih壆�/'݅-�����vb����ĸ�*�W�w�˟%w��n�kW��%4$='n��*���ݭ0��(���{m������V��ʴTS`e��H"��B�/Ѱ@�}⡓��X@�@s>3��V���Q�<�S��Q&���}o R��#�ܿ��G���Q[@�nl_��3��=��:��9�P-ы��iC̬̳���m��c�>BtB���}P�p�<ٝ�&Z���Ľ}�����OY���Ӆ��M��C˙��n�9�����|����b��o��T�B�Ɋo0��� ����v����g� �?�-h*�㬥^�N�yYh���ihV9�1�Q�,k�U��@$�����7�]_k��ԛ
L6�Yc@��d�N�ow˥���]8��=	�Foj�̫bu�����+~*+�C�(���t�`�����UF4K93�����ʵ�]
D���O8��
���	�%o(��������R	�<��]u��0��g�����z���C�/�'� ��/��8D�65n�+���]��fJ`�e7#��gbv[��Xy/��Y�}K�[��֠#�&҈��x�ڈ
��,I��|ڡ]z�wf�������!NI��o��"(A�Q��9��4��~/���R�	y�"J�%������l�Y>^`%��ѣ~���D�édF��@��ՏlT?Dj�zL���v���U���=<=�=�g�u5��'T=�h��~&3�ƽ6MȆ�2 ����9O�n%�1�u�z�Q�dF"�hL��	r%O�Uef�LU.��zl��t��z"�읷�=���W�����[ EU�:�Pc��Aj�Q+�a�pX�F�u�y�%U�,�h�����$}�St�U�:d����m2�#�A0�"�� *ה����'4"UZ[a]eiH"CS߃�@���B�;.�\�,���w[]D�v��bUw��3B2^(ڤ��]�x��P{���^�����+���.�GO�xi6b�Rn�$P���,f��Tj\~l���ˈ����T���8O���X-�i0� �����'/p3u/pvrZ2<��]Y��#�7m?,p��OS_0�������$b�E���"6��
B� �g�m����+aQ!x��Ow]J���y��`�ٚ��`#��Qf���|c1)��^6��)�齨m�بa]OW����n�H���1U����b>
�]ǜ&��
F������[�z
�[%��e[�Ň#����_��;���H'J��?�h� �׌�},a�sS��*���j��Xi���mT�DW�Vآ�*I����u$O�����Wc�1��kۊ:�}� cJ�\�"h���c�e�|
��������~� 
��M#�J��(Zf.W������7)�⫺p�n�T}Y}����M~9&W�T����߱�>-.�E����AA�3�~�8��Ǐ'~h�X2A ���j�(��#9�܉�� �'a������S"��1��x���|��~����Rn|6������h->n%+���Cx�����O&��3��/5Y{�˪W7��w�T��:����q�\ry����O>~�e�S���9��k�b�S��S���-*��<q��E�4<��W䩒ҕn��8����;�Z�y�s�*�^D�_S<�lY<�� ιz�x"�=�Q5���n{^�������^��g�@��_��z\ʳ �% y�!gVMaA�d/��H�k!�^��V�i�W�L;��\!�f�YQ��)��l�j)M;G�;Dp�h�j�k�r�2�|T`A�=��Sr%���m����,O�5����۩���/�	g9�n��4h('5���e�7յ���#����ߑ�4l�|n�g�fT֔���6s����ϣ�	����س�M��!���7�LH�D��%�-�m���iп�j�d���);��
7g�P�J���|��3�ͬ៫K��>�"_ͯ2��;)}tӎ��:���^ّ���=�r�$����4V@zT�Rd}"n� �B� �݃ ��M66�����"���w����f���+���A0�`1��K���IK��X�$��.5��N���?X?%ϟ%z�_`D���v�p��>o5��?����#�ӭZ�$o1��P}-��ౄ�/G	I�Q]�JY�._H;�-���l�X�Xe���9ڗ��7}�O�5��|C�N� �O7���6��(��ؽmrs��{����Cޟ�7�r�s4���[�M�D���@��y!����Q�ݲʨm)���K���G�r�e�XB����.�����d��$3EVR���(��)�~��i���������璍�h6���Z?����!f�L�2�s��cZ�U�.鱗Y�\�����!�`��]��^�ܤ�D��
�JW�`�;��T�����Ռ���Z��\��͑�^U�a�4�����5�M���S���a�]y5��P0x��o�q��j6��pD`��:?+� ��t���x� T��m�"�h>����2�v��>@�A�;��y�_���LwaT�F>���t��X�ٳ���A�����9�Ͷ�i�A������T�qȒ��Oހ�Ηsr��P�� %�%ƒ������BoM��1HS�m¾fבx]3ꋣt��a��	�,�A����e^yK�
e��Q�o������g9��>X�6��eR��dx{=�ťU�;� x��տ4 `7B/*[ș�����4A�[����D-W�6A���ELhcr8��nB��M���K��T\B&��H�����w�
�~M�a�E ��-���d�^�3��� �3/���������2׈hC��O�d��2V|��7�ZU�@$}�<5�K=�$���,�z��P)�ʪ|fu���D�K	<v��1J�)~�"���l��#�vT�r�Q���C8��  d���N�&��x4�.���y��_�.6XL�l�Hu��^�'�{] ��[�;�P3���#-`V=Z]�l��JM�����(����+D��;��ׯ{�"a:�dB���-1��9��<����[�5�v[�&��O�6{%f}�;�h�.WyR��+�@�N�ܿ��n�R!/���$Ҽ.�V´��vЇ��E\3�+X5�2�\\�G����[��9m����)O��o��;jB��C�R���a>�RT�k�����)�R={n	�
F��{�V�5�!t�.��L��H��7�/�`���b:YM:�l�y��!�Ab�@�j�pF��S�H
��^2��qP��i��{o����(����~�_�~i9UZ��0�C[��F�'��sM�_��׵73V�J�q�Gu�kfvtE1���b��c�:��v�U�ݣ���ܩ�n��v�;����=��>��$���n�����:�H+�1j�\����0��=��n��e]"��ì=����y�X�'['\����y���k���Te1�����rBaK����J��ڤ�*��$A�ʮ��0a7T`��mD1��_��0L�9QX��`,maDتR��V�~]!����uĐ���c�5�@�����e&e��V޽P�Zoi��}��k�vI]m���1�ݔ��;�|�b�b����;�����x�H�C@�#��bg�uK����V�0��=[:$��qB6/����ùN^c�
rZ!��}#!}ie�/�O���A�3:�ң|��M��r�\K4�i}�e��!�0Hc�ʂ!G�H�P�L
�,�86�+��&�����LE6+�ET��2	�w<����n�E�4��(x	r&_k�]�TOi1Dg�z���86�%�W9'LU[�QHD���+y�#��L.k�xٛ�L�#p�U�+��=�b;��S�-�~�����N�|��Sp�!,q��N_�
��9���'�W���/4�R�UߗSAJ�I~:2�3��&�!��8��m�I�ڢ�%&;��D��Gn`R��ccY$.�v��rUx�{k��~^%���Q�,��x�Rr >s5���U!�@�j>��cw	)���$W�O7���Bf�XXdoh>b�x;��gc����J]��|��f(8V+�F��b�^����F�Y�ߙh<�#��Y�SjuL��L�`'W���hG�F	�I����V+���*.���N��",� �)T������I==K�`Xp?�|ѕmʭ�w�߬J�1G�rn�����ݪ-Iɚ"i .�w�3�d!}�#��>$�*p�<Y I��VL�1q|����,{�W"52�����$>I�'E0�Z�GmG���8�p��������84�q��$���4y&�ItO�o��=�e�g"�q�g�2�T�����og�<y��E�~��u���5Ff@�g߈I"��낏̺ŝ0��v���Zq�U�
}�z�ZzR�i]�7�d���H��	a�N5D��U/��
�&���h�T`� ���|�'�+���)C��N�Z��AA������1%mA����z�}/u+��k&�P���J���:t�(VS�)T�%e���N����ar�Ƀ���6'|+��r`�D��T��MY1b��#{-� �v��<��#4���1|���'o�^�6��`�
\�� �;��u7�1݆(�3(HTX����m?Vn\�PR5�\e���`�����W��wamB���v��7Sz��w~Da���- ����A+���*��䄰��~id\���5�Y���.j9@)4�WJ�%|Y8�Y�b�������R"���2[?/54&)���,sK�yY78{ٿ?�����^�M�#s�׍31>�H�8����G8T<��� �
�����<�=��@F�������l��5Q^z�\E-!��̞�;a�Nn7x�<J���t�Rɰ_JdS�ܝ���jw���⳦���#��u�����3�Ћ���:�4F�M�8\ex^��#��"p�l�&�P�U[Og��;1��3�z�=۳Dd�>F��FЃ4��6���{i�Uy[[�S鬮ʯ���]��Y`�2w(��GR�÷��=��i�ju�!uLy����l�dr�\Y�ݖ聧[��U8ްpM����	����
jeL.��uۭ|C��D'#r��.�s&ٖCK/���<y� �����f�NҶo�|ĩ@���]��{��fu��}Aa3;a]�t�=��w�g���% �z,ljY�4�}ɣ�e�;X����O!8�������s��{��H?�ם[��3Y����H���C)��:��e�.�0d;݈@�<��h(۱߉���ɛm��(���J씡��cq�xLw����4kj��N��!*p�*��_-�iCF�Y�[6�IW�t	�h<2�6�;z��H�j��[* X�q���P
�7Jk�����o"-�v���t8)��$���&7�.��~~��hu�z<g}�R-{_;7�ur6��;�p���CKǽ,��9`�"���)}��2C�D�J� ��/�9�}�v���t���ae��k.���*�tG+�Π��
Q��d՞�2Y\~��.
�4]z.����b������K7ȴ�*�|_V��0�N�{��.n܏Qk�p(;�0�Š$�D�7Z��>u������p���J�p!����X�~q��d��gj#-���pr�x��{VW���>��� H����+���H�|�����A��Y�ןDc>Z����a�/�C 	��"Z/| �$o��x`�m�z� �ЙI�׹�7�xo��4���5��f���o����뜤9�i(w�D��]L�zQ�8</�\\�hA5&YD��E�� 3���i��p։{����x�36ZbB�����羒�ʭ��${֩΁�����y�}�e�o|�HKZ�/(�_X¢<�!l�Qc#V�o�an��yH��d�a�h��� Ǧ�D5(���c�i�ԑ.\��vч�ϡ�!-�<bz����]�7��;ɩ�y ��	v���!0#d^Ev��TI�Ʀ��4bD	.X�'�Ǖ,����ڠ�K��LH���Sc9Lؓy� �<˵��3tZ]%Qr�#r�9�л qꐫ]® ꓠ�=���UfMi7s[���6�S���ItM�$* e^9ơ�����č��#�����̋�HyE���F�&94~���غL�-�Z ����7��]���#��Ɏ�x�k��̿L�oY?���r'����wJ
��Ȏ���u�S�tĔ���Nyo��{x[�ą}��[�(U��Gk�P�s��s��P�Xꑩ�'1#I#*�����QA@1\<.T �ݭ]C�Y���+ 8:2�[=��i�<���j��UE��j����9���t�b$����k%���:y��.�k�
Z���C#6��Pڐ&��׆�ժPݎ���Z���'��S�I2W����{2&,6����9�>`��@�"+䦫㑐���o� �)�9&��o�زEm�����$X`2�`����=h�"�9�̗&�t�rH��^S�{������n�Ƌ2�t	�l�����եd�zŶ�ْ����~�v&��)��
kn(36/׼�b���/��7�;=:~�M.V��db�e'.��
�o�`yp��P6b�7S�O�Ʊn�Z�Kn&VL�7?[�.��)�V��Sd�+V�*p{k��+�-8]��!�����lPb�ߨ�"lް&���0�N�5q�_����γ�Sj��Z���m#��,w��J��#UC�/S�ʹAr�|5�$G�;�	����Yǥ��Ş)5�E"? ��*��8���爿X���	9��;�p�>���koZ`��Rx ;��'��/�Y���.���]<.1��\��e*������(��x�A�s���h#�k=\e�YU=�L4�0��H"���l^�2�Ϻ��(��y+�R���n�钎�8��C��N�u\�),�Č�7���L�dt]aj�C[���Upv�u.(:����R:��u�������O좹΁��"*��q;��ܮl��(;�.(��,sn�/�8A�e�4�T;$p^��| ��c񏺊��͖0j�H�O�����j0*N���,�Uq���k�4�w��:0�����9���3^�9�bv���8����a*y�C���q:mX�À�A�i��S�YP4o�u��ƁE���1յ��_���ݦ����{���h�\bvH�<.hf���k���;T����
�D����	��L�Q�kg�)�a	s�\ ��C�Fo���O�Y�\���y��|[ۙa�F���mlɟ&��5m#�_�ow�а�0��������րm���/R[��R�ӯ/j��~����~G�x[6!�^�F�"�--7e�n9R�e�G�#W�}A�O[.g��ia�[�z�eZd�u�3�wU�߅�/�['i����S릔)�!%�k�������5Ll�f��$Y����bmK�g�U�j,J.dl�5=����!���B[��V]�bv%�mΏ��R*͒#B^ZO0��%�~�[���<����,�;���S�u��<��1�^��8D��"�V!ƪ�L[L3�)�Pc�Ng�p9v3�ÀAG��lH�ܫ��a�$D��5��	B��
�К�-Zh�bZg���0�E*p����.k�/v���ՆM��zN�?|P�p[r�-�~�Jy+�Z��T s���i�fw�^��cô5��R1���u�����ӻ��Io}�U�Q�,�&K;B\����<�]\�g��W;�ф"@�.���;�A�w��qRW�t�ObuF�tu(YH�%
`��QH�$����9��A�7�\phq/�-����U,���o�v�E�.�un���w��CZ�L��K��ԍ8!�
�:�����N�m!��Ą��)�RҘP+��MV�x��H�Ay����ƭ����2]�&Z�Q���џc;�d܆�ph۲(`ae"�x��"}n24�+��{���Y���'^d��[IV���H&�ϊ�*dk"h�Q� ޹�'�Fb�٪l��ý�s^�'/�iTt�XR��r��w�^PG�*^�%5XYXjsEf���?��+�y	Y�Xn�'qc�)�d����x�H��k[VF�(�e�HH���*�q�64�#u�^�K/�D^�Hk�>��ө�XU�r�x��~���������sXΙ��CҎߛl�E�R�����\�����)o�̭�s(�O�t�DX�׭��u��?ڝr��#�w�?�w�M��\q!}�gL���9p���)�%��6�����%8�aN?�"A���1�����C9]���yB�6��#0��=߁�$�r�0���@�0�0��A\�
E^M�|줟p�+(z��lI��� ��z1�:�~O_�6<y 0��O]��'K�	ζ�����N�6�m�)�|$V�
�2�ևz"_� Z�V,�-$'{$��ia � [0�$��U�]YU�2��Vv�e�%V����#���YI�ǈt7MLd=k��>���ƌO<`�S#+��ɍW ���{s��H֠iQ^����.��*�3�0�t���U-ڵ�W�= ZR���D��K�@d�;"�yq��V����5����Ey�굍���rd�0��X=)���IL�O�S �QWnf�O���D��]ӥ����}�ބ؏9x�px?S��6@O���hF��)T�#̳�B�����o��q�
4�G���c�#�4?M}*�4�΁�R���������{(�+��� �M�@�Q�oX;�ᣠ�ƅ�O��b�n�D/f7\n!�@��G ��c�M���2 ��o�8%Z����bK������l�v���	���<��\�'(|�,v���g�3/�kd"��B��AI�����X�:�Tw�x���]l�V�'n�}�L��2�9�z�.��{g�����v3
0:!߳
�;�kT���b�k6��B���˻�x=��eF�_��`�a��r�FD�59?dX¸+�BYG��Na��A�!�<�񾜺}#�o~w�����13N������0���ia�K�R;��N�?�X�$5�a���"72'�ѽ̫���a���� ��De^X��06�kz%
g�I��r�6ΓG�bO�M��q���4��d1�q|H�7`��&��s�_ߧ�����[q-F��V1J���9~�6�;��p�S�O�B&�&�`�"A����9��f�q��Hu����8�of��e����ˏ��{*�"��i�͘���6��צ����%��rR��ek���i#Y.x|��󐴨�^⡀Ds�1���37���7�X4��������j�# *�y!�E�^<����'b�˴�s�ly�Uf@˂wA]�O�1�<��c-��0���.�>�R'<�	�&N�5��KMQr��ԾZ��d�ˎ��1u��N��P���tD�G�$t�1 ji?�Ƣ״!;�<D����r�Ʉ����À�'�Mk�Xд-���{BZP��i�� ]�������i���
y5P���LD��~i��D��^g��g�k�� -��)��p˝6L�t~���nL߉�u�z3F]5��t�u#�#�SaX��Y��F�m��0�;�0Y;��4S��6ė�z��4bDZL�/z}�v�!ʤ��:�KpFr�~j���Z+�F����!��%�s��T~��),�7Q�����q��mi|<P�ekk9\�!�)?�]��O����{]ڳ$d��%� ���טK�Ή�$2Ҭ>���Vy����T�f�a����R�f���Q�AV1��8/�O}�íjpM��ėIm?$N��`}|�>J^F$�{C�,~Kq&O�$�Fv��N'b2s�'6#�1�a��R��e��i����/K�=�U� �C?%�#Ь{�+l6�6�8�������(�?��X�]e�![��T���hPy, B��&�P�,�/���g��%�~�V�$��b��O�=�00�n��D�W�cEaV�W��w��6n���ac��Z�,�#L=Ǯ�{Zq���3����s��"��INh-,Do��h������o�қ���=Y�T��c.���jf�6~P���7���>��a��i*�ŝ�,Tp����M F+j���/�r���N#���_����������:�!3<!�glD^���*�%y�?��xa4e4����$Y�=L��%Ť�C��4�6C�"RR�02X�t����3h���`�oV��+���7���J��Q�%�����I���SmP<b;c2u�el>'ahB�	��n��?\]@l�*xugh�۷O�g�Kd�?h�b�D���R��>�~���U j!�H�� �T�Z���.����������_]��3q�	r�Z�8z�\�lb߀��fQ�������^xY�1�M�4��V����g^( �,�D��1�1U�	]H���M��/�%R4��i���3�9؉���} %ԅ��l{�p4��5�c�K|�"{�hlM	�C�����uX%)�{ VP�,J�
��̐ [��]�<�����K��I��1��w-J��3��r����O���!�K��ObF�f44�_r�j4VPӍzF��J`A�W���%C�zݠ�=W�x���M7�!e}Y0I�>Xg=������]BSm�?R�>I�\%7�ѥ�z����cF��
T�$��<=�e�.h�ڎ�
7>?�.�kiSt���<}Ѽ�(�U���ʂ�=;�brZZf�$����Ͱ9��"aJ�S��
H��3��lr��T5�B���[����0X�\A�,W���6Fb��s��)����3�G�A��`�-�������%N���.�n��6�u%�Q9����k��\����XQ瞑�v��@&a@s�mT�48Z���-�7xK@��{����)�<^M���\�3�K�$���_y�^��#�F���&¹�ҔR"j�A�(�uQ/���%���q��.x�!]��^��A���(>�	7���O��F����hkP<2I=�f�/�`�ڭܔK|P�%��|9�W��w'_n���DY�7d�k(�7>/g�,� �0����{�$�E��*�pY�稍�tC���(��pNf��i�t;xysxmo�o���x$���dOkY����A�h����]�m�m��8䲇�:d'!f�\�a�d�HO�>4�6�:���i��{n�u�B��tnX�`)�cw��� #6ĉ	����[O &����:�(�;�V<*�/���V�	d�����e�ˎG�����0��sx�����C�-ƫº+)�y��ob-2�"$|��$e���@�RG#�%�Аd�b��sv��I�W|C<-Gӗ #r׆8j�l����꫒ ^��7�#�a���q�q�)���m���x>�c���x&>���X�"}@E\MII�3��F�k�xB8�/ޅy�To���d��
��a�e6Ȕ�p���&h>�r3<Tx.2m����� �-��[�	+�w�����'z���,У�pA�۸�u��"����'L�'5��|N�H��(`s��c�G��M����NR������Ub����_��s��&����~��}���g��>����F5kHdt��*EB�a��2�I�E���*V�i(M�:����Ǔ9��t�	��'.����td����!q��v�%UYp�p38O(��zWj���i��UlSt������68Nh i���^w>ߐ�R�r�_1�]ػ�����x���ي��ꑸ]x��%/=�8�$c���=�d�o�	.����{.�1�v�\�T.?� 1��� ��E�^ 2v�X&g���5�n!|,S������\�$�z���[جv���< �~z�U.��flB/5t݆-���ӆ!�¯ۊ�t��3_ZL��3CD4Ss�nF�Gm�5ⅅ�KU+�Gt�V�a�;������r|�����̈́�| ��ܽv�}�w�<�������~*|	�jCnSb��r��I*��zyP��n�
S�`Ju��LP]?[̧�{��l��虊�VM���Il36�W�)�:�^��pv���lQ�2 &d��zT�k��;�!y|������@Uj���d�3�}����8����P�;%g��;�q��#V�K��>D�D���b�H{.0�¥n{�O��2��7��ttb����vd���Gj�g�\h)��KˮU�j�r�d;�(�����[�"��-o.��;t+x!aD�����Ŋ�b<zՇ���Di��kq=38痷%Oh�6�d4mh�&1?ֿ7(��.N:��$�`aX�Ý|?���{ճ.]l��#R���ߓ^Fa1*�
/{�$�6DL���a� ��u�j�R�׳��bͦ��3�t��d��˳dY;� �a��@u���°Zi�m�UW���M�ӊ���V�a X�֌�E��M}��(t-"H�^G�G\�Þ��� v�ѿ�dx���6W�dxL��[����zY%n�=艞
�<;��To5��/mU��p��\^���B�h�����d�k��eqb��\�+��8�F���`�E#v�$r3i&O֔vMM2E��ꘀFs��c��sJ�so��q��J%$Ȟi��#��XfU�}�1�gG���U�aX��޷�e�IۣR�k`d���Z�4��V��1��z�ڢ�>�Y��+
.��(3�G�=|�?�g��Q7�n�L&E���k�H�!,fǡ
�-Z�uJ5*�h����dԇb���u���Z��>y�v�@n�|-��Z絎�y�W��%�Ρc术]sQF1��,����#���zY�5kn�
��Ug�K��pso������Pg��d�z���<���lڬ	9�/�=����Ω�����ӏѕ��%��$�BT)���觓� ,N�E\=�.4�s�+��<�&@� ?̕w�� ,r�0�$L1����x-���%��[�"�ڽ���Õ��/���۱�~�)�P����ts�i|���P�k���������	��,�����i�j��(,N�Yg,�ˍ.�e&��HW/�|�(��Z�Lp��1�����6	Ǘ�.H>~��G���\�e����Ѐ���]�MK�jt�zQ�.��>�[��;��<�f��R�R��1�~z, �-����4����.���$[R��w:f%����\�A�Hyfgl� _��W%W�0����Z�$�Ӻ����Tw�`7М��p�{/FK�����L薉	
@4��s{3K�#�F�����5C�Z���\7\)n]���[����.�O�?���9�a���	}}�d�z����'�Q��x��2�q�3��rR&���a1dH�����YVHG��PTI]����,�q�\�Lhj� ❽ht:OF����}���~�(�#C?R���N��όf���k.#�_��Ъ��/Cn�1�G ��-7H^"�8���߫��o�&nv�C\U�n����m�y��^�:C(�y�%��?p�W��WQ��V�_iǙ�V\dKAD��*�D�ᓌn}J�I� SZv�C�."�]a�4�X��4�&�g��?W�8���9���tK��[�i�aTĚ�ZzcLf�gα��r8T`Z��)��*�*��S-5x<je�̜�8�1�79	Ĳ������?��qc���-Ԛus����ptQ��]�`���>5�<��f�P�v0����I/�4�XK�d��+�7O��7m�ТXZ��s3c�Ћ�JV؜gϋOe��6X��ƨ�'����H�'�p����u(�d���0y�-�Nw@�4uQ�e��k�U7����J�T<c_p-������OȌ��"��o(�$o]�t�l���`�3g�W�ơ�l����V/Μ�ӈ��Y���fx�Y�w.���q���B&mx����Q_�Rs��`޷g���������!4P��=�l�E���]�~2(H�2�^B�-�63��i�F�2<A02��-,���O}�,O0�*�=���[�ꛓW���~xG����#Ε��/X1�X��'���6L��6�ߨ_M\�B�ѩ7���2��qr�Dk3������s�m�p�Y6F��K�lˏ{�������:�~0Pʆ��U��B��������X9���Bv[�9�pW�GH7R�n̵p��.W+:e؝P5��`�*�;��=Emi%5��_�/�P]����e�ʥ�?�(��N�qJ�����@fw��ݜZ�����cr�W�gv������7���{�v�y�ڶ�%NR6"A�cE��l_�	���"��~�w�s��^�j"`Ny�c}e4�xcǅ{Ȃ<x��Jt�Y��G)��Q=z�Cn��7�����lyi�1�*q�Gu���ѼuU�����l�(��,dZ`e�N(�[���qb���ޱ5�F	"z!�eRGxʆ?���c���;�1٧�F�#�)r8�����9	� x�-�O�'U���zK�7ʟ,��_x�_��%߮��0Kq��UHp{�Z2���n��y��T��y��Jk�-~�Wc�\OC�U#6�}O�K�QSV)�i%��+E�.(��y&���=P5K�,LBd��B�=a ��D*�-^"�g�<o�� N��}��e<]�Y�?ub@z����z|�0�p�9h��+���I�>mDO���/�d6&�cm����������5���|w���<�r�ؐ�T|]��6����J��0��p�a���x��=O�;�bԒ���чlZC�����j��j����������O�3t��9����4A䦾^��n22�O� �k�s;��~�6 ����NoF��f�$�?��C 	n��M��N�nI �?W`Rv��jb�OYɩ��`*�P���fOh�+���:�f����1��KB�����1�u-�#���+E��t���+���vM�ZM���:��E�zݒ)����P��� ����ָ�����Fz���ǂ�v̑C�tb3 ���	`+�(� #�L�Eߵ���F�\��#x�k���^b�R¸��c�4dqVr�ͰS�8��y�m�POe��	����k� �N"�W�S����r=�6e�p�N�����l��+z?l�e2D�I��[V^ڲ��Tz�?���^&���0��а���{>�=�V�|��x��W��U��7A��MRjVn�	k|�����`��)��g�n82��)V�t�
�-�b���Ij�����6Q�o�/װw�3�������.���,	��M�j��J��������74�Z�Gl��Brْ]տ���O	�L��b �(��Kp��V��� T�ʑm=��{6���A�a�N�+T5�c�<>z�d���\�Ө^O/�%���0�r�Z`���]�mf&��.�M��>4�Y�t�_F$,֟��
�ĉ mË䒤'�*�yJ�uC�.>Ė<	no|����Y��pD$
<M���a��J�" r��m�S���ã�qE��=S��I�z����#jOL0nT��bf1�R�+uW`���6YY'ٝ�oE���뮝jca�XV&v���
� ڤ�V�9�b�p�ϧ�,��#-�-�]Uƾ�Kҁ��Z�^�d����e���v��h�Y� 	cd@F#�*gdu]ߡ惖@S%e���ݵ�@�1)���?�6;�����G�( ֭5c�7[�`��Xy�tz�$�4�
f�Ba�A�ݰ�'u��n~m�(�֒d��d�8t��FqT���N��D.uׁq_t�,c���c�[CE�zԏS��,��'�������fp� A;�`px�Sd��K?�&O�`��,���$�^�p����d+�3�֊��
��H������(b�ͷ�h_��yu����<��uo/X򹜷4�91}A��\�v���߾����M$��E�r�d���g�������̡(��� 
�b���Z����^��i ���3|L3����܄�w�p5�Y���r�ךs2���D�+��}E3�e2��������P*uO��Jf'�Ԣ�`��Y8�T�Z�}bɣ�˓q�d�-��#�����F.0���$��|���-TC�] A��{���Pm$�\��(��$���!慒�J�X�8i�̦�>U�;*�-,�Ap�'�C�^i�Eݺ�u���si2q5�X����^�dر'���AP�T����Ӎ.uP�zH;�Gn �)-U��ׁ�������{�4+� :Xz�-ਤ������S�F#^�_�t��\�r_�t�s����)�����<-E�Z�
D,y&t����7�>����<����{§���ib���gl�>���������i�dzl�l��vA �򿲉���]f%��?�E�Л1#��r+65��	���-�(�*u�� ��΋����.����\�}2����-��$6�l?�\��^97Λ��l�F���r���>�{�}�<D�����mr��+@��~����~fτ~��웳����5���P�D$+�~���`�ʂ�abs��A�ȧ3CD��%�;f]���[��7CbĤ����B1ʤ*�:F����ÐT�������1^��К)� L�,����ᮍg�m�-c֗�D���6s��w��p�3y"�V�3O��/p�����]ϙt�2�e��ʋ�yX�-zS�7�+��I����0��a:C��=ܸ�pu�I[�����nX�!�X,P����p5�{�]B5�*ݳZ��Ng���Ը�������s[����Lez�vr���,8�^�a�K&��K��M:塱c�A(�����)��36�H�-A�8�o�^�T�B"S����~�D�˳,I���`��m�L�׆�25���3�=�����qT`��|���Ry�D���c[�:If�hF�inq}Kq�Ą��M��%�}j��#r3"�l��!�2�=�;{=�)s^�uL-�ӵܰ $�y�%�+���s�zU�lJ��IW����d�M���D����2/Ÿ������b�i+�8h�;�H��><ćy�k	��]�U�^�(�,�;��/��
��w��V���s��~��ޣ2<����~�3�1V	t���v>��.��%�e������"���O��-G���~\���̟���R�����u	#���t�
y*�N� � s:�U�j�[H!!�v���� �Zu8��{X_�L���gW�����
q��C�0~�U�
'N����u��D������6	m<�mܜچ�#�ݎ��ztk�Ჽ1|�@di���ᷧ�,[��7�&�vb�v���5�x�����o@"��tK�TC�|�1�Za�
:Ӈ<��ᦔ:Q�y C���򶂋�E>K8����{�mx-]��%��J����A�1��.�:*�Q'�@�R=p6���nv���!�J3�������[U�rl����;)���$���{d������
u�2�BRӎU$��	��n}��hd�����>+�~�`���=�Џ��$6ݵ3V�4-x}�_���F*&1�&q6��o6j
O��ǲ	Vg������č>oPc�7�ա�,�Ǹ��8/k��'����TG�Emm��QN��T�:��D%H?�Qyƿ�	�
M?����K,½c��Fל��9�S�Wb?=�i2�,w,U_u�jz�L��3����NJ�p���?r(l�����X�Đ��r��e�+T1��;�%�]�c�J���b`aY:Ty���@�{D±��dFQQ��O\����__w-p�{y��=/�bIk�ބG�)���5�giY�L�8�
Z%C)_���y��5�i4�Lz/+$���V�8�YG>�*������T��`�pt���Q��m)�5�I��L���8��f�1ȡ$���d�0�k��Sny�R�qX�����ws|��p���%e�RRw���W��3�|������\6�t;ZRcm�	<���t�~0��UrY���:�p�5�k���4Sk���P�lk+{ӓL)�V��g�=w���4����s*��s�^��e��^Q��l�I�{B�ڳ.�^$����:+C�����G�Mq�`z��bM��Q�
S�L9��SLT��5�1���_mS6�JS��ӷ��I/�-c���zf�=t>^, �>�0|��;HW���,ɿ�e�ӻR��"�ɥhnyC��H�1���粓��%'t-A�K�e��u���aY滣�ݚs�=�]�z>m��Si�	#�4����"���&ul��(5��>���Iy��\DVy8n�0��Ao��_�}	v��j-Ur
Q�7e�YvÝ��6��FLy��nj�$���O8��:��C��Kv��HNd�Ĭð�h�F	A�ۘ3�:%E6�}q��`���@�a��5���J|�6&���X/"�3�($ mW��b�Lv�U�U=�9�(�&K��2i51�.�ü�ny��}%�? ���N���2�,�^�7��F ���Tƕ�t��;	��*�;c �U����?T D��"_4q�XԘR�q��%�tr��7�����e#ɕ'f^��8��V,4^�^���8=�^ܖ��f���@0���b[��	H�*���lx�h��"��/�9>�|�3��P)jb?��5Q���&G���JI7)���# ���,h ��q��N��	��"���֞��e|h��}�2���N�n%�`8EgI4H��mZ��p���%uYu�ߺ���_q	cٌԁ��X�	ڿ���Z����0-�!0|����hhe9�~&r\v�ǫ��iD^�q�'E<��s�����m�	z�	�T\n�Gн�]�Cz�f������\�Wn�0���$�y��~���>�f�۞P�	��Ul2� 3��_����a��"�d��D �� �� Η������Wj+tg������nAa'�8�
�Hm��yU�Sh$����|�ˣ�o\^�Wt\��iD����ь3�(L�ḹ���~���R�
W��JXF�z���K�B��6w-� v6�3����?#�"�f�x���-�]������-�a���Y�֭'O����w׺n��t�YL�6�͈���B`7�M�I˾��d�>7���O'��b�#�LοQo0Bl�9I h,�&���EH� ��R9vd�+V��^�8m�l��ޮ��h�{�/���%��( Tg�z�d�O�s�'b\�)��1�
?��!�q-��=����?��^Zo�@~r�Lw!b���9q:y	R,ϳO&�k`&���Œ��3��V3@7�A���p$!����~�Βdb2Z5YW���
�1�@X�� ;��[�Qs�ǌ�-B�9�uT{��k
q����Y��� 	vC�k��r7C��H�w]Q�|�S2�����Y��D�t�k�@�;(�M��i`Ҡ7d:ӈ�
�O�FǐTV�&�ۼ����Ζ䯨��e�˟Y�Ŵ7�v�2�e���m�/%�����'P˛m[����:�1Q��i�-u�i:���}�簩���� �3���o�d1EJ3�&_�z֔]�2wO�=����,�� ܪ���ǉ�j�C��	�r�C���P@�ف*�/�r���i���Co��8��*�I���_�.Ğ��E璙m��B�E�v��.�$�|�-�!qW��!Z�~H�Z݁���l��l+����;4#ڬ9i�A%ޏ�!��9��nƤ�,��[��5/�"��f1$� �1��5@���\�f�Z�dk@��c%|96Py~�c����̳��v��>r͙v[R�Ҥ����|���������-��[I���R�h���o~��I��{,��'�l��r���>�6>>i���a�^��*�S��U��0�Tz���S��Ǧ�D��}���ҹ
< ��XE�K�8f�q���ʿ͂\E�����yL8���em��%mi{$1?L֫4^�S��*��cUL�~��A��$l���&�ٷi��|01{�1�ڗ�6d&��5�1��JD{��9�!���
т���^P[�G;�9^���J��?�q�>�g�������!��93w�M�0Wr�6d�k�;�eWQ�E?TH�W��9x��5B;���H_�A�^��f]�^�T.��3�?Uي#9ֵ4���%JF��זb����k�%��}N��p~
��.,k[KH,��N�F�ӊ��ĽI�>�s2
��O��J��f
0�5a"f(�g`���S ���~��!Zj�ԋmA�Y��D[ d�U) �|�凌l��$�!�#x�0��a^�"��@@wC�meO*����~()Or�G+?�Vt;q.,TݗJ���>a�$t��I�T��cDe̩3��fOòw�Ѭ��Y�I��ո�����Ip?g��;n%��7ٽ�LVaЋmR\����dV̠���6x0���C�������]
��{�4�
_?}�1��	վ�-�5��	��Z7�r��h�m>��ܛӚ��[@q��ì�-��u���GI�j�����ڷh��l����Aǯp���ճSv�_�s�>�0}+9��I�?l;;E��lZb�th~Ӏ�z����hٓB\��sh�q�qK�u�x����1T.�T�q� 7��s��m9��H��*+��z@.�	�I�� 4�ZB�Hf,���D֛K��Ei�˽�>a���'E�(.�O�q���Yi�̑�t];�x�Bpv5�R!�#��#Xd� ��x ���l�A�-�f�޼n���Ƅ�K��)�r�!� �k�-��τc]Qv����:D�*�?���ɢ ,/�6C����Q����3�<g��.V��A	�����?M+/���.#}����AEO2�w�π��B��t�y��V���+�t򕓱�V���B������A�B\�R��0�a���A��3�"w8�6�y�S��[�Ǝ3А<�����o���Uus�C5&���Z�,����2Z�p8(��6�Q��q'�/��D�w�'9`��l���q��o��ŝ�<:����Cˀ<'�ئ��s��N�H����=E�%����)]=����.=cl�
L[h����*!������ �@�_[���Vbٌ�$�C>�k�}bn���+YS��V�$�E|��h��n��[['��G{�:����w#�u\�xdQ�gH�U��Rk���#e0�pD���OX��fAP��O�(MԂ4w1*m��$��H�F���K\�)�X*ZDab�
R��� �d�b�}Sذ�ً�%�8�I`%��5�8â̍�غ��%�"6���ؚppvR3q)v4�^$*P�P�H�_x�����m��g�G)�]{/H��{��`j#��:�h8X"���]���%�&m>�}ֿ�Ys̆y0��z������G�I,� �&^����8��HK�ծ9����M1�=�P��e������hS!bm[J�1�3xhqt�m~aH�U4>�~�u��H�,�gSl����QV���!f���Cv������r6�M�r�lO�:!���=��&�fH�5Z3fOϓ�^H@1���d�izi�k�0�.]�Mը��5��F�?p9.��:T��j�p!�����>[i���u=�:B�>@g�0�Y-g����κƜh�
6Q[�t���������m��w�e�t������=��`<D+k�֌]r2E�a�.9���l9��bgs(�9"{h���ផ�C��X2���aU
)� W� 堹��[��"��nO�}#>6�ct��}�4��H~�yWH �>,J�xf��A���(�}�3D���)��˖CX+ח0@����\A*�R��,x����|ШD�̊|@�0�%ϗ��!�a�����{�P��F��2�&a������M�$27uxJ
�S}	֝�w��끤tqx|����9�]R����i@��$�bf��_�$�a�c-)���?�iآByӳN`�-���@ӨP�(t���T�mn'�C��TVObzM�������(����j�8��晸�-�g��S،3("��{�ԋ�}r��?s�67��H Bw���1�Q�(tg�g�t(\��>6L71�{��Y����:�� �ĒƖ�El���v�}bVs���a�X����	2��q&��+L0p%G>�=��)�2>�X%}@����Y�}#�As�����8I�!�DBz�ϳ�d�_��FX��d�Y8�	���E	�l{��j�-�r���[D��0$�,��>��޼�k$6�G�G0Yh�Zל�՘m��@��ĖY��zR��Qh��k�nTA��BH��! �� @�B�"c(�I��a`�\��9�Vce-���Z�=g'Q��H_�Ǘx��O��*�H���L�]z�3�I@�!��%WyzP��JdD�n]R��4��W�o��YcA_7��O�)�mql�T�pdJobT1D�4O���Ty��C��H�TLt�s&�'��KSY���7/�
���{0�������9�Qv�xH5�8�oF�Fz|z'������6�C�ԂE��{�m�޾Bj�#3��������am�����$:�{8���w@k_���iB_���������-�����T��"�����U1(V ��8yg
;��2�i�i:����XMl�_�����s�@�i�^���B]��R�B���dj5�{1��4��$pl�*F3���ӱ����V���U�0��sN��!�'�o��
 Z!���m������2��-��R����b`��u�n}^N��+ȫ�+�����e2p�(�a���^m��z!��ȵQ2Ɉn��U6�}}�p��g�n��6yC+7����+2TY�7�T�O��kpT]ԯ��Ѳ����Y,SL���ԭ�� �k4���7/�tz�����w��T6����E]���m6��E�,�����(ܯW� cP�������י�&����3a��.0t���YG�>|�3('��l^���y�gPC�tC��l5���B�C�Y��:�ói��φ�����P��khcK�%h1�m��H\lJ:����c(J�:V-<�~f�����D��C.�LJН���-��mH��g~:�@2T0�×�+m�SkP��U�d��D�ȉ��cE�Ԧ�*F�O_ګ�?��7�"+ҸFx������.c��گ^S��PPB�����@� P��+>Ў��]yʕҸ)�'"e�t`�&�R<	6#�̧�VoW�_���*���;��6d����˭E�=_l�4�\�-P��7h7|�:81|�G�V w��"K�c�`�ӟZ�Q+�Hu���u���$C{=o��d?�ř���E���Ao�.	������ V>Y	i�
�G���ѱ�H�/-9�YF-)Ȋ�B�	�٘�
�`�+���!�T�X�c�
�Rz�����H5�Y�-�d��\QT��B%�v���p���������3
����TT�"���E���R]Sh��������+�S����"Z�?8@�*��+��qn��vc�AO3�r �/��2��]_��_ �>:��JK�]z��XB,���sh���o��Y�Z�J�t�oll���r#9�Te�/}T�.���o�tĜHK�AƱDǦѧ�����'x�;oAgGx\>ޗ��7յ��w!�����EXn��c��f�����q���t)��,����f�����˦�dj��P;��܏�M�Wl�>c�X���H��{5/9*����TT>N��~���?����cס#��BA�u;.�MY2�e��)� �edz�
#���y]��o�a<Ǿ1�!��C�[<-�Ue�~���4h/�+q�1��V�\�.�f�S�`_�ٛ5jڤ�p��[�ܷ��LzA��֡�8�Kd�xz�?�O<�\�ԡ������PWض��ꨋ�B�LRz�x�Ɔ.��j�T|�]�H���rO��9TwU��Ny?A��_)�ʀ\��;З������?T���\�K2yQ�J��d" �7a����:vs��u��ъ�VS�������i.��?���e��^�_�V0D5bUA쫤�y�h���v�^�F��`�DZ�!�5 ����O�H�ѲTFl�<Է�kU��K'.���v�Zf��U��>���6s�8��+��Q�ƣ��$M|AV
�־߁��lfb���~t�I��4Hΐ���%,������`s�^��ĈH×��yBW�"}R��@�� �%��?��$)!!���f��=�F�Cg��p8�C�T&�ɨ^`hM�饀u��'��QL�2h�b1��x�u�W��6M�pu.���έ��!/x~��'��7��r�����ZF��}�Hr_MI���0d]P1R���}T��"�Vq�L:�Q�����?3P�!����E�C�-�~��j��/U�;��֨*) �LL-�tJ�b�
��0?�(#��-.�=x�����TߎP��L@}5l�����m՘H�X�{�b�T�io>޺k}��I39"dw���|����lw�)����%7T�F�/�	0ɥ��V��;�a9a�ҵ���+Y3w��I��V?�ӻ��3p���1��Fռ�3m���͚�v� ��h����N.�T��*x5�{؝a���
<p�yֲ��K;���"���x[5�Or50}�V&/wRu1I.�4�.���MꞆ�t�P���'����a��-���ڋ�t·H�w��q?�V��Xn��Z��qV�*���,M@F?��u���֌(V|g�M ^���*��K�L��-	�R������E�%�e�tED���>y=�Q�c��
U�*��/��#N����&7����vu�1s��A�-� a���`	"���3�Ern�	�S� m�[��pTNoJ���u���-�g}{:#��ɫ�u)4����1Bfd;&�S&��]Y�5R���u��W҆Ea���3��|}�/�^1�m"�[�@�
[d�E�z�Uՠ��@y[�)$���X�:d��$b��[���PR��9��_ث�H�6b��?F<G�k�s�fv>��?�c��_{4�+�Jg��-�K�j>S��ӕ��㎫[�-��3�~�qz⤶-Md�,P�� �Y���[>��m�D>��{}G���·l-߆�e\���h�)ȽE��8l�H��5��)���}���]�Kg\��5�Ø4��ޔ�\Z���B<̒J0R��>O��噦�\l0�S�8T@W��,�C�7*����ƙ?���M�GB�tz�KUӄD�N��ל])X��A��*���P����hz����"��b�=�)O%p��I��_j9��lH-�w赊r �K����Ҡx����@��Ig�6�FKP��B�O�<��I3u��}�U�6�?\��`�$��ab�^B�s�9�Pʂ�u>��٠=�A��.�e-�T3 j#���j���*��%O���j�s��EmeB���[�����)p�h���}����'wpp�iu$���lӡ��o~u�+��֥��)Au5�[�;�r�f����eg20��G�Q�_����Mjc�jgX*��6ګy�tH���3���Z����%&�Å��x�A�͓���Z<��8ּt�m����%����(��t�As#2C/QD��(h�g�-��oJ�5���o���tw��H ��F�%��ؠ�=��6P�Ʀ5Ypԗn�K5��R����R�z(�g�E�dG8�71!�5����T�`�y�@���/@�� t|�?Z��}+3�����^���TI�K,��
���.I{�f����<f54�zƕ�Ysc���4�����6�r�b���A�@�9+zd��:4��[3O�mF�L�)�:
S�.����l( y�$�����y�T�
�Br�ޞ<d������(�1O��"�D�e��� �&�T�-}�62j�g���������� M䝿ဗu�	ql�*Gr~�Y¦}L;	�U�>aW_n}�o��$׭&e����o*�����W��1#���H����r�,}vv�/�f��}� ����J�>�ƞ*�C��(�\]���ƀ����j���Z:��l��L���}���b��Q�B��cx�����軆?�Z�V�6Y��3�Н���l
T�T�@q�^�q�|��h���"y�S�)A[��-[ ����ۇ)��f�IX
1#��%��*g.�m�e*=T4{�>^���ͬ q^�i�>.T!я$�_���Y�k#�g���V:Z�F0&����3�lf�;���}4��h�x�_!(@מL�����ľţ0F���j�Ai��C�cP����ƒ(c�br.�ʲHQz�bm�f����S������2�2�ܘe#���H�iR�n=Q!��P!�̼;��/2�� b�<�@�	M��t�XC'�a�u�!fa7��A��ѦZ1`����{�2C8��D5D��h;Z�nJ�_Ĭ��E=��;�������	� 3���Shu����D��Y���c6��̖�[J�9�#',X���ZE��}����)�Y��}� �����TC�g{��"/����Oqu.ֳ�O��i+�h�!����bJ�I/@e!��a��$��U";dQ=��4���w)�{��c�qU���B {aqy���
����2F ����m��IY���r�;ْ�ڌ���5��i�W�B��5*�p��Z�k|���S̈�u��X��0s���g����Q9�u�tvK�;
M<8�`0tw���Գ^�6>ɢ�Y:D��s��"$`yA~�Q
 ��/�������e�*:QrL��`/�R^E:�p�ϓb��y�J�v�Y)j�|kL�<�����F��O���A���O���Z$	~�yܴ�P�74�l(��d�;�h9�JQ���+�8KY��o����r0��P	y$e�?K���<�i<�C�c�#b���Y[n%r��ci�L%)��Zr�X�i��֟�*To�GB����y�7�@�X���<���&oΊ��&P��N�`�A]]���(���	#FmSsFY<95ڨN>�mx�͝��raX��p�k�}�cĶlM���:�F�D݇��ޜ��'�z�ձV�e�TH�!����lX�N�:
am���U*f0"(Y5�w�(9�"�c 6����.}�M�Hă�'E����w0��3A�Z�j���-C�*�K�@�gU��9n��vL�0��f��>O�����2��W�������G[��:Ti��L�/�7��X�%3m�w`0������rl��W�[K�z��HKp"��`&<,�/����{*a��$da�̆�\R�h�̑s���9����B#]u�jI�s��W�Ga=�֪��?�3���n�z˫�1��g�.�x�����J��b˵��_LD�j����G�úD�e�c�To��Gl.�k9)M��8��v��O�g�E��P�S>N��;�^]W�ӾV^)�g&ސ(dvk����4�x�R�����e�y�i��1���Ō��Dr%+)��W�f�M2˾X���̄��P�a�+E"�ՔTE��qw�X�i��U�]xӺ��7������c$AA�`��'Rb��];����mBS?'���q�7�F����|D���	A������f���k���_��5���A��SU2�|s�c�Q�J"^H	3s֛�,���"&����\���+��'�7jc$c�Qa]p��t��R���[0��+��P��><t:�N��s4�6��a�BH�h2�q�_�u������Dߍ�Zd*Iu��[:�p��N����>mf%�48���n��J��[���R>)$Mµ��ә�?�`��~q��y#�e7)H��
8iY���ݔ���Z!�sM�/J��ഩиFjؒrT<��Ʃʯ<��ݞq�;�/����) j(f�f��.���H�>�ph�.�.1�[����u��a��(�Tl`=*KY]2���n T�=�zo�y�'�z-�R�ek��HVBh�I�dP�����L?�cD̴�,-I��ޱ	�g=�v���J����=��pk�#��=�)�����B�8z�>�8~���+�E_P����3:��Xw��_�
�r�������w��##x��˅�\4W���.����)Tӧ�pyf�qa�m�t�֤�����}sm�X����Ȝ��io��B�kH�#dv�Y`v�#`��zلL���'TK:L--}q&sqň��4��aS��D�@'���/+x�s��ÆW���)�	�|z��8����_�����6������Z���:�Q ?��<1�I0�z�^͡�>�qy`ط�ݐ0��;�1k0�11�]�
�C�\P���ȚK1?�m6��3���<�����$�ۇ�!US�w��U���nL3���;�,������:qNH.��k�U�&�4]����0+��牝��QS_����_W�������ċ&��R��5��6��ye�Y����7r�:Wp���V��vu�[�&>�6�.�h]�o�O �)�:C����?ed8T���B�mO�j��"�/��\e���I �/Uu4�a�(�W��XV�z��STh�ϔ^ѝ��LT�fxˋK�r2%ȕ�R`�s��r�Y{����!!x��ξ��F�6^��sg���:�f
���<GI)�^��rBZpg�����^�8_�رЭ葆q�p=/?f��/
Hlz�$^�������1�{���rz՝�e�d�f/�N�g��ު:�wDd���b�?��������o"�W<���΃b�ϙW%�@�C�""P/�/���)���+�&����3�QPlFu ���8�T�3n�*j��^F��27� bY�`�� ��A(-Ob}%�ƥ�Ab�|��n1��?S>ѣ��F>�#�Fl�xf;́��x��f3p?�BG��n/������Б�����R0�Q���z����LfP]v.U;���U�U<3T"e���d6��A��&+-� -9��Q�)���f��Y���'i/\����,o_J��'4�������kZd��I�)��:q������ah~xT_�E!���,���ވ"���"��q�KP�%yu�Z�r��ZM���Jd�ܶ���t�͒u|�k�,�͇��Tg�Vv��)�(����`9$�����/&\"�A�B�LF�y(u�Q�..����M��z&��M�����5�K�,�@J��}ӬM���B��9p����_�HŴ3�%�O�Z�q%�es�<;I��H7s�(�����=���p��������&�UV�oWb���l!]�t���L�
�̙����h�YM�:�������@,�
�wz��暥mmrȶ�s���4��:�:��gl�/Bk�>r��A��\��jbc �����\�=��������U��j�P��]̞��'�W�()mx)��J�2�+���C�>�帒6�|��D�`*uzg)�>���E<LHob�Ս����i���i�����w���&A�/f��vbx�͊�|��X�f��cZZ�^w1�a-h [1]�j	� ��o'Dp�]q9Rm�~q��j�r�f�Ҁw
k%\����8��p�9��},�Y&������͐�\�cS�h���Ɉ�F���,�y%%�ĲJuJ��u�:ީ�FI�W�����7��oK��=���'ocQ��<p	�.��Zw9���s�@����C�j�<ӦW�(�8�Ad;���I8(ܚ8'�l�{��i[\�a�+����SX�K(���v q��f�O=�T};��� oó�e�L8��eD��\�iX�9)���.`A�dW�C����~T 
���z��V��1�� ��`~Z$���`���?O�@?d;\�
�Q&���[A�vd�Ƀ1�@+u�,�Hg9Ɋ���u�5X"�x΍��2FP���C%fe�,��ˉ�>����b3hO�:n}��>o��Қ���C016�*i3�����@O���q���5&���Cv�o�Aw������
��2n��=��>$~4��Ӻl'ѳ�"f��������1������R��<DHŒ/�ܾ[	����L���L ��?�����h"M�h����Ax�s��C�N��"	b��@dO�P=�p�a�B�%	#���)Ճ�YYW/ԑ�.	#͊�tα���l�D9޼�*X�h����*}�lpw��-���A���o ��T]'����h�e�I=���� _����h���	&�0�� �jKh�V��;ɲHk;F��6N�؃�ۗ�����츁:_�Gb��@Nnm�/��7��&�hD����s�S]�L{���������Z:�
ͩbr��[�Z6�ج��~��M�M>��"f�п��!?Q���E�AP��1�%���q܌n��:ט������R'Y#6�ɥ
��63J���u��n�k�y�f��K�_��3t�"U�����_&ؕ����e�o�T�'l���&"K�&�9�9���m%��&��(�LL�2뤒׌��(�K*@����ZU�>q�LR�e�D1 �d��kfx�ӆ�k��{��bQ�-@ⳬ��G~�/�υ�?�&��*��(��f"��D|`�pSX�̴���^��W�F�F�5U�bJاY����	`K_ݥ�cK;'e�#7L��@����C�j�B�^rX�R�6��b{ޞ��5&�k��A�����x������b�|"`v�uAS(&�"ǘ�;}u����\���^��'������h�=�m͸���qKj����퓌K�x8���Ev=X3Ӂy��4��pR����^%�	тʖ䮝w	f�"?/%�&�[���P�rWF�<�˚ ��Hؒ��%8�]��T�a�_g��p�y����9�T?�j�������n�J��MMčЄP����$@��dHi�'h��F�h������=��K�4������Q���zM<�|:��*��<_~(+���-_�����Th	��$�5ȈK�ě#E�C�\w|R;F�aP�������m΋Q�U�:Y�^�Sr�C�Ï�a�H�4��Mqzpq����#���w�[L�m�}����4�Y���@d��z�0��2�T�u!��#I�i? �۾�I�|�w��A���؁�;q�H�8���ui��@��K�t.h�\QQ��0˞/�p �b�{�QԲ��ף��� '������O�Xx���}l\���=6&�F1S"Q��K7�������>�a^�
Nʆ�+V�:p��*.30��+����.�o��r�F)�� Χ ��	FX=�� T