��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jåا{�\�u�?߷�dn@6�zf��r������;��1�ŏ�%!�W�pWF"���S6��6�[��v�V��<c\�9��d�iw�� ���=gݛ���L;�1H�����+B�
� �ŹL������v���8�H)y2�ּ鳞#�Ơ ��UBX)j����o;�ȣ�B+R�MGU5qosƓn�9��y|OOT::��uQaD
5�}!�9��	~7�Ҝ�?�:�ո~�	K�#����.[�yѰkN(�v]�� \q��]&�c� �( �ӏ�-�:8!���з�Z�S[c�Ϝ#�G�d(1�Ǥ�dnnM?���B���vů�ײ�yn�8η��U '��. ��@�,o5a,`&��[�(S��$� {����8�yD���"��r���L�"T��i��T��^<�$�0Z�̬�=F�j�tY�wiP��v馩P����S�D���\_��6th#��,}�T{���9X�1���)yH�֑���H��zC���P
��X�)�k�x��c�s��������Wj��n�JV����-0�q��w���l��_xf����{��tqQړ����ǬP/�a��O|����(�=)<�����f�KR�~�b��M�����V{����ʀo��/k��9r"�&���㵱��'{�q�h�A�;� ��_��:�����X�4��Ƥ�{��
�����C�����#V����<�TŅ��;�ҼJ<[:{"(��K��I��)}\k�s8NH��>g�"?�f1���R��F_�\�[?�(�~��S��x5�6<,N��L2e��qW���W��R�X9N���Oq��ìQ����9���Δw?%���������49y ��u�	fe�dZ(�pS����O�:���I���|��n��쾫ES{�}��T� �M	�(_i�G�B����`�2.=8Pa���n�Z�ɬ�!�^Q�mN���j�N����G���w5�D�X��?�� q�K �'ޖ�t�������س�+����B�6ۨ�5E)�g�A�@��Aj�����hV'V���ȏ Y+�S!��n{�B�,7:���f���w@�U��[�$��f���-�,`,�{8n��\n]r�E���-ۺ�f�#P�2XrH�>�1D�r!����N)���
,fY�O@V�d�3 ���"}��Fk��oNz�����ٟ��h"IM���|�nf�,M��,SI�=��:~ľ��+bJ�nE��p`(�E���tS��Y�N#w��Iç<�9�J)��c�s���x�Ĭm��K���yd.�i�3$�$�fVH��@B�
��.w����g��������$Qi�x��,�9,%�y@�ȒVҀ5��Mٺ�K��{
��ٳ&���S$�u��c�3
�8���x���ɐ�U��<`L?Ƶ� <.�Gx��k��7�^�	ّ�,t%�3������2�~Bvg�K/����GüXqi2P�7|�����Kh@��@���ܾ��r#3�����cI�)�`�����l�h��o��.=͔�D��ECVO��$9�G��R՜�Y߂���~z�>A0iܨ���6�Q��?.),�VhmFGG=�U��`���Y�^�BCyt@��Vx�bُ�t#$!=1�l,� ��-׾�h�̨��<�
�O}�]BY�	<�ݏ�>ڧZS�w� �D�`����D8i����Yʍ���Hv��H�Շ��)T�C�4�h뚠jM7��\h�3:�K`Ŏ� �i��:��G8�n���aGKi��
E����Q8(ώ�.y��"�&e(8��ᡅF��N�G�Nن���(������"1��I��r��ζPd���J���At[�!��<��ѐ;@��
>���M��2��J���D.���/�,���������f��y���C���өF�q��|T�hQ�/��]ꂹ@-�$P���!��ǲ�r#���$1��~y��Տ;��)��.,��u���
�x7g����,��6cz|��>W�fhg�v���(�+� �jǡ�=�<F.���6�x&z����Yb�uT �/�>�di�q����e�P�Z���J-f�}��b�zfٹ�F��j����o;�l+���r"�H�O`��.������s�X?Ƕ��ՠ�TK�UNc�kF�
������z��>�-���]��L��4 {<
�?��pf2�b3;�]KJҿ*� Ir��:"���W�PvDKP���M�|A�[ߩ�"Y�|t�OE�N��=�O틵�ܮ�-T��A��n���W7�1�=M��R�2��fsx�Q�C�Ɲ[�8,�Y3�t�t�H��6�\$�����T��g�3�1��;�tޛ,)�Rqz��4`�c�\!V_^��ZSP%țH^ظ���-6W)B5WK���,K�Yro����O��V+�&�C�`����HG{H�`'��>� ��l|�Y7k�eL��/+�l���긛 ��q{��Qળ6��B�s1�����#]�q�G�'�CIК)��ٯ+~�'M.����/�2�ϫ��[t���s�T;��fEC��V�5oX?���(1�u���m<���e꺢b쎦��}��(�bo-W���I�� ൰C�O�zt���fԂ��Q��'l*�M@�ǂQ\��$�p��J�Z"�M1�4��#�R���)�������8��+���"B��Ve�ie��*P@ʠ(�*e�'�Uq'ヹ_�f��q>��\!:0����k�3�NxsK�h? �xq��Cځ �3�~����g�r�2� ��Iq{r�./d3����,F�T`�.(�8���)(��aa�VOة�=),E��NC9h����l�q�,��{߭Qrk}Ci_0�u��~��>�.��_��Ūt�h��HQb�Så�i��,��=�\U�F�v3�&	\rK<=.n�}ѩ@}|�?���M�;�����ހ���ۗ
|�za/r�&�6UX��j��*"ϲ����|Z�i�M��G\��ܪvB7SM ��=ž���ғ�^nݢ
��P-Ŕ��y�^��Wh�N��X�f����}�cǬ$�8�9Z� ����K��}����N������jﻤ�W�)��/�8��&�Ԏ��l�E%o���h�7C��H�����T��E@�+�e.{1��S~4�����~H�&A���M0���[ �9���E\�p��yx�B�vtFr�e�l^d�㽚N�0��?�ڰ2�
;��a����l�}��&��U���u0B/[,��X�f�L��`���P1������u��{�'���]W�IG An:��ߚ~�����w��r�����cʲ�)�LÆ9�|/o����{3 8��ӡ1c,�%�!^���u�rR�p
�����B�<��TÛK��Q+o��<�W�����o�J��{J�OV���ɘ�X^:���Yo����0F����bI�/H��o�� _���k	4$e{�Ay�f��ی���J�uE���_�������jMa�c���E4O��.^R^��Y�yi�2�I��ރ���M����Ry�%9Նp�	b�%_�<���@��x�S��B������m�������ԁ�T%���j����nZ^����	ޯ9�G�{�L�L�}8�P��Z*�H,A��{�"K!�F_���K�p�U���L� �vuC%�'�Z�/�m��L��;5��%l��e�S�+�)�[լ��h3e��y���f�'~�[Y��~�²�3�ZjC��֭�gʘ�Z� �h���� Yg �
�B'����
�P�.D�5^��_i������9�&Z:+Jo�b+��Y� P椬�_�����7���^Z�� �"�L��� G�u>Щ���g�ڕ������wљ�s�"Dq�]�9�p���#�Zz���jp�QH��?��*�:�K@�WD�+Kr�mDs��%B�������;�I��A}�IW�Rkf�W�����9zH��/�{	�pD�I���B`��4Y� %/�,Fx�$	�"�M��	�]�o�+�fk�ɘI���b8?�4sJ
�i��m��dD�*��4 @��8U�t5��_ϐ�6?Q����A�1�\�ܥ�n�'io�1̳�ØМnmA� :���D��޻�A�Ƽn���u<��k�XA�;s9�@t�N^�CG^ޔ�����C���2���B����v.��z�B�y�p�����U��[ű^�������Y��:�o�Hu����#�4�
ʼ�x��+=ph{X��{~s�2�9����9�E͙�7މ�䬱H@�c�R��e�b�M'�=� F��Km9��y��ɚ�Ҭ�O�y"?�7�� o�^�RՔ��<�_uE���	�*"R)5�g(f'��S�4�QG.j̪rR���f�_�TJ���exߖ@~�ݥY��T|��o��@!4Ah�������S���K9��v:��N�-r�ɏ!���~�J�|hk�
�x��жp�4$e���c�8�%f���o�7�5�t�ߍ�)]-0����.Ǩ�/��i�<��(�Ii��N�iQY);�� d�D�<衧���~da�wc?�sGW��!��+�m����?���#��R�A���K�3�����W,,c�>V�LSXh�V�98�}>3�P�k8(�Av��-�>����I�!-�IR=��u|���E�y�җ�{xf'��̸�f6M���)�k�2K��if�J>3vғ�| ����!f�Gϻ�w��ʔ̸�Jiı���'��4� x�[kE�+�U��р(���^M�GNƗ	�uUrN}�w<��k�	Ӟ�3��;
�����5$%X�k]G�h��(����c�1��*���t[�
B}]��$��IAO',�r�l���mʟi(GI>�
+��Np��Q/���톌���ٲ~ՏFu�J�:���Ԏ����}�V6=]>>���G(���w��W��!����*�į�5��^�RK(f�}������Xi����A���FS���o  �V:�*��(%jB���e ;��v�G �Ђ6Ty�R�7�gK�;����YC�~�UH����r�g���|K�+s���[�{�B5p@�����{�7�nR�R�o�Q�C��
6�B�9���5{�!"(���S$s[6z���y��,9W��<��~j�R��B�[�S��0�'��N*�.��I�鼪���F�N��/��{�(Z�an�B.������<�I)�Ū�䑃�1��7*T��O�s���E�"*�W�^�䙔���U=��h��1Ӷ"G�eN�R@��_E��|��'�}G�qe	�p3�K���H&D�,$E �69hض���B�Op���׮�R�
�i��d�T��.� �:�\�nf���j9ٰQ�f����t�o�q�v`:��2�|g%r0";�oV=�Z��1=؈��zb�5���ٱ
;6V�溜�@և�j����҅�\��@��u]���ô0���9o��8<��Gu�b��Jғ�d���4V�,39�*ܞm��DlQ�{]1���QU�\���gE�:6�K8�����ה �W�7��IG��&T����+�IZ�٢�;/{|�^������ZEtD=�)��jm�^B˜�\7�4~eY�8� �1*,��ĥ]�;3�G#f�4 l�����ϙ���������t����m>L�hS�J��n?�����ڛ��$IS�,�AV� }_����ݱG �;����0��GC��1؂b������>~���9�X��h�G�lz^��l���������)��԰Wd-^�P;�Ȯ�`9;�s@w%T=��%��7M���eg7��yt����e��a��4sB2�鐠.�Y�)��Z-$�8|K��h��7�.��H����}�A��s�LO�zD�_��-9�E�CXL����$Jd�#��{��ۨ�-�3��(�S2m%Sh@��'+*���lR�VQ?2!C<%[w�/��y�(�,&�qR�ek/�Zv���)�<PKT��
v�ٲ��rV�P�6Sr�Я�cC7�vF�(j{���$`��:��ǁ ٨�����?�j��Rz�����2��yyILrt��l ��2GvN|S#Ǟ8�d��#���%�xt���Gy�?����w$xY�(
�'`K�Ԑ+,u�P��J��n>�vLo���r��:��;���Ϣ��8���8�y5��~H�R����<.���H~��qЧzya�$۲�p6�>w��dh�	�W"Bd�^�2�_���c��:L� f)ua~��~9mI���|�N��:�U�쾼]%��[��'+=(|O���;��D�2�J�Δ�s���qq�"�(���������'P��� �&��tT��zi.736�!x��H�r`����\u��y^�V���ϸ���:�e�@0+��Q��8�A0J�e7���W2��̾�o��+�0���/�����2��G���h��3��s jRl�=��i�����8�����d��u�����Oeҭ�n���å���"���9�o��NN�Y3����;��%	���P|�zC{� '��H�O��t�.�3���	�m�Yc���)!�y$*��~y��ۗ�������.���V����ÃD��J�呱*��U���1�EG�N	Lp��s6c�1�y,ƄG���A!f	�	��':q.]���r�O��;��k&������A�-��-
m�u��>���[M�+;_x�ՏD/&U`���[%[5?��9q
}���9�v]S=�S�f+�Q]��ƪ:1��NA�x
O�\+T�o�1>"�ZC�6&ӿ�C佯��#���:U݈֜}�6�/�6Yb5���K�� ��]XC���;7�������9gZ�U��@�m4����K� ���|d��2f�K��aLj�Ɗ�G�RqL�	�+��je�S��`j��n�����.��V���Q��!u���^�Q`K'�ę���Ĕ"���Ӕ��ܺ�T�'FV�~Y��5 �'/	�����"�N�O^����oV�BdZ6��h���S6u�{��r���d�*n���HB����e�F���j��lAr�����W�3�j��P�w�g�^s�36w�Y�"f��L����Y>���n*����I�@��]!�4v���8��K�8�H��ϭS�t��[�6��q��"ஈ����㄁��p����й���o�=Ȃ�ؕ�P6kB�	'�e�Ό�xO�y������g��.���:M �9�j�����h%��%�5���G�|�D"6���(����Q�T�{�(e�S..��C#�,�hp;�#G+�	{�DB���'�������LPG[V���[M�&n�2%Q���N(2EW�K��R��U� ��fy&�0ulIkH�7+u�1�u񥝸�q� ����0��ʘg��/>�(d�ezE�|6Ǣ8g�zT�Y��G��GW�fvG��:%'~)ԡ͜�x��F�8Z�eb�@�����$Ǟ�]dE'�%�m:�)ɾdZ��-W���w?w�[��S���[u�2��0�e52�h��
l�_�p�PR&�ì�����#0̳0�#c����K{�Z8���-G^�> �gTL\�KU��Y�I31����t����&'����^�M��ڭ��!�V�a��������ʓ���:X�i}j~��������M��,?�� ��S0O��z�X�߸C������%/9Dce5C��|�{�͸�ѧ���R���l!)Ͱ'��з��pa�ԏ�]f	�o�6F�0��Kg��Wtdy(Y��g�����m�B��k� 3`��MWR8��^je0?.@�-�{�mE�i��2�(D����C�����`�up����ׄ�ư�p5|��/��l�* T�`��t���̬��d������^�m�E9Z��zbzʑU��w�ng,0�1�P��wra��G*����6�\�����cY^M�����l�G�$A��r�`���qI:O�`պ���(�|e\o���LJ�]:�ǝ�\��TG�Q�t�:��.�bDvj)�*ݰ��{�����A%G��м�Y�/���c9�A{�
'u5�Ŧ�t��&ۡo	������-F<˥Uq@����R!��W~s�0���P'���7�u!)�-4E��E$|`�];�(d�$��s�8v8Z# �����b-�f
��1�s�>���_�Y��/��"������1��p�	�#A�x����r�&�fH��v_|�5��[��d~����-{�0���:�>�Uˀ�������]���.���p.�����l�5�wT�(Y��H(h��0�~�&�=�� �؜��s��(N�K�K~T��<�+�R���Cn��		��5���PT�߷�9A|��ޤ�W�'�,J�knl\K����tƃ����"G;�䆙�,�DTm���G���Լi�0�קgf�PG��δ�-��Nx�K8:Rޕ1Z>���!n�Ǔ2DO�wS�E,��́�x����b��xq}))��;P/�,��
��1o#��.Cu�m+8_��h<���j�5[{RV�|��L�ſD���(q�{c�&�;�,җz�Q��oq��l5�~ϰ"CY����H����e��0��n:��J7�Z�.��]�ȃ!������<��p\
%�L�PL��`�8w�6u��)��	ÿ~d0@��_@�S��bL96�l�th�JXx��M��M%֚��$����=k�Cn)��tw4Iݶ~�pT׾>�c�"W\�}��j`l�|�C�c{�3��7�}_�o&c�s�-�ʈ���t��$�Wv�T�Y�W�N�Vc��`��Ә�l8����Y���+�y��ʗ��o3�ǫˆi��p���)���@��
�'���F�_��|���0�?��Lre~\У��}q�&51�7�3_Ja�k����-��K!Vk�ѻH��z�]'�A�^�˼�-n��J���X����99Uһ&>j��){�bq�hjtwĒ�G�ཾP���uk�I��=���=A��ӆm���h	y�^���B���>X��������K� (i$���jׄ
���JZ����`�R��zh�˵'��/���y�b�2�qq���K��T��e~��7Y%�¯јI�I�hQ�rM�&g��Nts��ꃐ����uQJ�o�9��`��U��F��}|��rkm�E�o[�D���}��	D���;ʹJ�IȺ�l��Jr�}a��(E���D�XE ��%��,�+��-8��'A�v�H3�����d�ɒ���-NB�G�+�������|i6M��h1���XCq�.i�+:��R�g�/EJ�G����K�s�0�:P���. ���Ɇ�_br�
�~�'���s�Z�7H�DUS�nW�I<B>� ��'�F�{������.2���Sْ�L�|�)�F�Y\=]��x���6����-��+O��̆��Z��#��m2�{[T�}�J���Y'�)5�{r*����5�+U�H P�w`G��֮�EMO���__��c҂H�*�y.W�#�%�z|;�_� ��ȑ�9���M��U��9KX[P�R�d��c������ �j��xg.�c�;���hi�ZǞ�5��z°��I^lƂ���a��c$`�=��0�)��%KtV]+{꽽)5�%K�ģÙ�����c�λ)���ĸ��������w4�
�S"|��9k[U���ބ �G��U��Jj�(g�ɩ%:�n�vT�~�α��ɎK�t�_f����<�K��A�8�4�sw�aP�J5}��)���7�����?�6���ZH�V���B�?�إ�.F��/�"�1�z�ˉr�~"J���1[���q(�P�ZYl��J�y�u)��hĔ��۹(���yd�-q�la�9���n��{�@}��X�,^�+�R&NI����;MGZ	�-m����}9*q�8(a��*w������^m�`���n�/.s~/vE��^Q`������èë8���7p��T�d�#�I�z4l�� ���ߔ��	(~+Ǝ`жՇ��BKA��yD 9\��ũ��"�[�y�{;_kʺ/_�K���S�-|!�?�m䙨���:W�!�ga)�ǯ��+\\U�C�������-���3�5m��G���HXސQL���}�t"��A�Ïv���먦�����\˅F�(B�k�h�\�H;��yu�c|�,�ڿ�Q�/�Eg�"M�o�Ƹ7^�dx���:���J���⼒��U���gB�%�6�FZ	�-�+�X�x6ʀ�/��m��EL�Ę�o�ґ83�����E�Fj^�l������^�K҃���3ػ/N��.u�~� gh-��'�3ʚMAo<{�L _�^�4�[��`U�v�^�p^u��٪":E�R�Ts?����E�4��Of��Ǡ�1��7"�C��GdP��z5'����`xF6eDdDC��,���������:�G���Y�B�b-n���.�7����x���7����#�������ay�D�x��B�Ϩ�<���t���˂��M�7���a_ \��7t�?5����fMf��}'o��3��9o!{!
0����6()���תcR�FÞ���������.B�|���aM�����I���8K�Ɛ�7�~P�h���by�#Ї}�����Vj�R��Fن��0�$�M���QE��DL@$yZ(,o4�u��}����o��ٞ
�ӗ_$t_C̨|��� Üp��|����.l	$Ũ��c,k�D�@U��˚��щŽB���P�UQ�(�:/��c���$X�t�<�Qd�=�|�Sg��[���[{�A^�`�G�B���|nt�������r��D�VXs���[NeW[G|`ב�����jW\�/�}� � �n+2��#ϫ���nG��)^^���vflu��x����/�<�$A㻦�H�`Q"L�s��ͧ}&.쎃�o��<8����~�F�p5!�щi�锗R:h�x�Z��."�&�H����f<��`�J�!���3��x�P�{K:9E��%c�n*J��n,�v�%�����o� :��{�Q}L�Z�VfP9)nY���[E8�}�a�J%�\�d� E��v���������(�C�#j�W'���Y;W�r����W�NdǊ
�����H���w���WfKl @�/�T$jij�x�c���÷>t�s��9��x�!�J�i;i�?�7^a�E,<wD;8��ּ��f
�k.�j��Y�\%@:Z$GT�pQ���+)kpۧu�;;�򫇫��j���"S���Nwm7}��}����`w����:���k��r��1��*3(D"SLva��R4 V�a�~�|�)�9�=\���������Я؅"D]��~5c��u�����+��� [�
 ݗѠ�$J��IȄ��/�Oþ��={3SK�N��5��q'�.��	}[]?ϵ�3ܩ���c�=�tG�#-��	D�]`4f�v1���J�y�U�?������������O�B�_�"�3=փ	I9�~�Gb�߳Ɔ��E���8អ~��;�I��I�>�^��4�$��7=�P�T&PW�X��"��h��XQ�0&�&�B�L����-wRs��3��RĐhN�`�MC�ٍ7m�@��k�Ԉ�ǳ��a.j��B��"Y��#���U���K����~:y�� �?��R���Z��bu����B ��M1�P�[�8\�!?R�鉠�����B^4�<��I��k�0��'' �l4J�0�c�w����t7�崅h��Rh�:�bm��FԲ��Dh&`?�t�@�o8>RLƇkDw�PT�.�Yy7��O�l^ �Ē�c��W��Js�zP`����B��Ѽ0�q�-�a����N}8c���`�$P�����PEm8�L���<� *�gX�%���!��N��	u��xs�x�����Y�
��	_��1����=�Hb��ytC^�� Ԯ�pi ut��k�V���tپ,�Nx�C�K�����7�ei������̇A�^�Q�͡�)Ig%8���+)�z�&�P�o�����4h�i�#�`�+��\Ȫ7�έs�3�;�, �wo�L|(vY}ۓΧ˼��Qv�U�5�P����l#����hb4���"-˜E�{m$&��QSx��)�H\D����$�	�oCL(�@��[7���O�~!�.�G�(���O8ܥF��Ts4�U��:�G�u�d׊G(�c�R��ǾA��N�\�G�Y!W�*T|].�-�={-����� (�� X<k^��m#�꼷\��n�	�vgy��ՠ��J��r�qj�/1=m�0�������5��p�����Ɩ ������ʜ�H��LBD�X�3 s��۞��Ѝ�-(��1:Z{��h)DhM��UW"�2��p���#��?��/ҩ��X����[��^Ti��7�9��J���d�q�vSW*V��%��T*�K˭����)��G@ɜ��F&��MwІh��K�r��I&��@Z��Fsc�>P�dn{�O,c\d{Bux�hp��Z�sx��{(;T.U�sH���cήS�^\Mx��4��_7�?~h��'rX����_��������������M%�P���/�U���g�B�R����L}��8}�љ��xPg��6Gj����%��\��g����W�;(&l�g�Q-&���6�����f킕L|�5��7~[2��I_ [԰ǯg[���3p� �;Q>�[<�Ɏ��̦]�XGZz5�?�nӶ-�t}	? {��`�?��)�NT@�&�㿖B�Ԗ��x�L��E���S�"P4'.�N�>,� ؽ���	.	���I4Eg�s��:�M����!���N}�ɣL���oy�؊c�j�]��:��-�e�o���C5� �FQ�଺������/O�C�t���(��n��{m�G�Bj�ޑ}�]�;]���s�G�J��Y��q�.�XE�S��k9��V1�G_̎~�LW�!�&M�(�Iݝa�����~č�� P����z�23���q��Н��F�}��#C�k���9
���K��! <��Nl�VUl+�����8���Z��#u���J/'4۞�~�1�P�!!�&1����M^z�:�VKyף��9�o=��3�2��R���dt�1���7�rE�}B�?4$S������z�����X�����D�k���,m�u�'��}�Hl�f�"n��ts:�+ ��xL���6D�T���ۯ֝^�+��+�¨�?�,K����