��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jåا{�\�u�?߷�dn@6�zf��r������;I��BJv2r%�(��c��
��*C%<u^�ZI#�j�5��e�\�u�E#*:�]L.i�+ݖ�U�D�K�t�}w�	�����`�����M�I�*�T0_Q7���g Hq�ո����X)Pz��v�� 1�����Š�`!�/�`ZfPL�ֶ�	�M�cM/�߰��0{�0���Ŕ�<��TV������aH>E��!�7���~ݛ^��;|[Ep��R���S���\ \Δ�d��/5�q�>���!����vjS;.j":2L�
��H᧨:6��q�ו��?�ֈ¼�	R�j�dΉ����H���~��q4���0LD|�n�|(6�V�(�x<���Bץ�i�Be&|���K��2��;G�6�����^9*�!P��b�}.�X�un�	����@�>З|v���o�3]��l��h��h�p��;-�އ̧���¨����!,"E��6�u|xV�0DG�|F�w��U�b$>�Q����ƃ���ǈ�R�ʬE��sH�;�h x-���pL2�����p�<�^
�<<�8	�VΝb�c��3����^3@i�IG�7�m�5b�v�Cn�(�Zw�}���XE~s���y�}���6�zZ���R1a�8=��笚��"H	���Il ���g]A`cH>@F����Cp�2>��K�.��O`��go��,����&]�P�b^��䙿a�(�j�<xdxOx���d����CtsPz�����i�#�V�6H�Z#��n�̤p�8䙎%K��o#�pV�enn��{e������V����3Pp��C^��(��-F��vO����-<��:��m������ʟ�"�e��j�H�a�s�ę�ϐC1r1:��!l�nDF�C�.N���m��+
��ʳ�8F�ڴ�π
��W��b�j��ف��a]�7�ܬq�n��q�ݳ��흽�C�MN2��Y���{n�p�̾��F�2�d��ī�zK�󩗢G۫vf���pT3w��u���Si��� �X����H	�c6+�H</3�#}��l�W��:A�m��%�N���Jao��4 qb��ZƬ���<&k� �F[��\�b�I
�+E���D�66	��Pe?p���:��`YaL �%�L�7Fml����t$J�=yDa��Ճ��#5pO��8|8\T�{�_mW}�R�/ �{r>eۮw���Z/��Pi��5��#�j�������81�~7$�H��U�d��`TB��^�k'���NN�"�۔GRF���s{�^)����e�}tϺ,PΏ��LO�y 3�E 0�use62 �eɽ�]��B=��&A]�u�I�����1=m)�<sR�2��7@��1�'�ο� ��_�rU�7%����?��uU�OF�`a�~��d��ϬV}��+aJsת���9��h�[!K"D���������n3��@<]9Pl�"p�1{����x��Jv��pô�˽zy������5#�5Fֳ�U�f�D8}R��u`"�7��	��b�H�4'��/�5�S�]�=s �|�m
��x��m_�CD�0d�d=�ڼ�B�>����,I����?#Pք4�.o������6:�f�i��$�/�oA#���;!�g4� z�K��/�v���w�:��A�)��uOx����E�5$d�oh!�<&�G��s��&T�}U�c�m����c�.s�s�y���bI{Vُ{�c�g�h���OrM�ݽ���w'�yVb@V��@�Wߒ�o� �
Bs�ٗ�I`I ��1q��林*;7]P��c��~������ϭ�qQo|�8Utxo� s�wO�R�����g|^�-Y��[%������WWo�C>e�4���bu��Lʋ9"��;�W�y#E����x�K��(���L	�.Y|Jq,����C̥A_�Ԏ����� ��cYo*H	g/��$(6MTY�H�����夸+��pPK�����AI� �]��)���qW�TS��#�A3K�Q)���S���
�����{k���ܡw�~�l&@-2�GDq���ѯ�(��� ���HA����PʩVU+󔚨�
r^�S�v�����������$#�,���r\���~i�G� 7��b� &�=�����K���1jc�+����?6{���� 2Ŭ�
1���=�/����,s�SL�^;�����򀳳����Y܌ԍ��b��(e7��2�{s�d&A�D�<�`��h���u�M:e`�
��_�'�p�5|7vM%��jxpx�
���Y����aٜ��V�K�3aa�N��O�3��֪w9���@��gG��8�iu8�^���)���Uװiv�1�xW:cU[��[<9�����v���A_��'��{��V1�ӽ5�dP���A˞��c��@��/8����4��/�oW����@�p��T�9w<����ߍ� 	���l�Eһx�j��,�,�=GT�� �	�������Mt}����ָ���	��{�ڜ�]��������5���̝����a��aO0��a�֮%����ZG//0 @�����u?#�C��e�R��k����O��@6<ـ�E���Tֻ5�˱R��e���U�[m'�J���q��0�}��բ�-|����3QԼ���:x+թ:�S���m��"�O�>�)j�X�A(䠤W��레�]��&0�H}4UBz���b�
W�e��:�2c�'fUr�&FQ ��7jw�9���]
�~��'�r�H����#��+�7fI��O��i�vb�s�@�2����nf<ݤ���x��SLI&�UA*��D();4�7����ჲ�=�:l#�[�i(��{d ^M?	��|���	���b��Uv��n��[�L��=�i�R^�kކ�V#��}���1����c$��S���[�p�|L����`U�hg��Y���E�v���?wƚ�&���Ϧ��kQ�y:�CS�FN;��H�aQ�,�p�ks�Mn�\l�(6	P_�c�5+��� ����]I�6T�y�%�#���Dp](�@��{iH��ێ�2\t�����p�GC�3��L!y�(PD�� �L������䅊4��hsF,N��8I`sK�����C����W�[Z�D h~�����OHc�<�X#��*8�UD��jf�]�)���&�Rr
oB��o��*4�]��HsXIl� V��ڂ�j�d���S�
�퍨��[S1Z|X�$w���F@nĐ3[;v�O�w76U�]y�?фGn�#�,�m�:i�)a�K����L�K��� �,�_>��c`B���3w�fY�Gs�?(��hD�|b"�T��2In J+�J���&)�)�� ¼�q"���|������Qӣ�2��8�>:!NC�(#�?��#w�N��OP$�t}ǿ��Yl�la�I^�)"������v$��v` ����M����t��ಬ_��4�kS%�{�J����џ��ᑔq<K�8�2�*
���ʠ�Nj����rhh	C�:Ъ7�A�}�D���i��dqˍ�|Ƀ�g����P��7j�L�ڰ���e�8�N�U�1f��O�{7�&j1��u��+)k=�<aU˷��������Y"��e�G_]Yz�/�R�y+Ztb�u�"���.^P�W��"�	���?Jf�T�4e���њ.�����I}>��d�����5��?ϫ�$�Q��� �
?M��A� tŬZ��ȥ�E';;��F]2�����`¯^?��#=$�7�E�Z.���j�lû��丘��4��}������v�����aE,"j�x��u�W�5(y�Bˁ�	�*YL�}�<�v<��(L�K�f�c�I��d�R���/z�(�5]C8q�{�����)����	�s�Z�Ն�ǘ!u��:;�,z�Y����x{0A����]�.�c�������WU�|�|$���O��7��&cm~&�I�w��
В�o��������l�ӍSY�5��C��2��o���Fd
R�����%ƅȐ^�����}��R�#I���.�=�͢'�%͛ѲnFlL4���"�Afj Ղ?�x;�
[���<t��A�)�����Ծ邗p�@�F�C ���σ��	�7�$r���LB�T/}���>����Ҥ�[�*�%K�կ�a*��X������;�aQz��崍r�MA$��l�ǰh�{ڼT��\O�M	h;��ê���+=����Q��]^SD��4�#a�����|��ůW/o�p�"1�.$r��k���G�|�=���<Č6g�f�ۿREα�O�����=n��#�$�����ƚ�ڃ��hɃ��kx��:P����uk_�O���$����(oɐ��y�1s&��K�_�y�{�6AaΧ���ί0���h�^�Nh/�m�q,-�p�gb�hGo|dM�g�D��t��Ck	�3���ݻ�!��~���ov�л<�`�C�x�sc��8����2��,e�@n(	���C����SD�(<Pw��B����c�w[����:Ǌ[ڢ5�玚?}CKrP6$|4�]bZo�������"�H�}�]i�tw����e(����!�R0nv�!b�b�{)���`Kֱ꟪f�� ��&����U"b�Q��S굞c�1���z��xzh� ����lo
����+��8E�o�4��ߜ���7���K���j_-
�:�q� �j%c?f�/��3 �^��K�#_e< �LG�~�.Y�1�v�i�v�"�z�����)>/�x��{���jKf�;��E�"8a�C�p�� ��x���=Le�(Q����l��
=O�q�����0�N� 3��
�C��T[����ѵz��g5��:m��^�G��0,O(2 j/cas�7M-���|��g��"��qo,0�c��zZ���\�a���><������6��e�.uX�KS���=w+D~�z.ݷ.y:���S=0}�E��>ʆn�����<y�*�����cG��AH���xX���j1��s��&��� ]���Ȟ� )QKn���Bs#��qi$kdv�7M9��c�Z֫7�#9M^�V����o]���W����up�w���0�}?o9-����g�������^'"`�����Om� z{}��MT9a# K�竲* ��{R�vu\w��^t���R
hu+ٰ��h��f�E�� QlJ�v>c��!i�=�s;$�8x�m�b$8V�a��p�}ȇk��q���73�>����s�-D�:9
��<#i0�㤂�������C[i����BƇ�Z1S
�,�,ȶ[����|����Y�����jL��cI������-U�r�Q#M:D��c�E�3��&Ę�meR���G��oѽ���[;�u1�H�1*z�"%�m�>-d;�>JYe�=��|�Ԇ8�v�>�J���M�:AC��.Dy齱?\�C�1�t;=��ŋ��	xg����mݲ��j9�C�M�E�y�J�����16p��[��B��{�ݯ���J�t�� �W�[�%&T}8
6���M��������!����*1=;s!�ر%�d�ȻcBd
�q��E<���1_>٥�j&�J���4��(�~xE��mG��W��[��2F�<�i��o� z��V�e4�eܕ:#��!]��c'�駋ua�����;2����]�� #Q�5]Y؄��_��1�Ik��DH)�ZZ�(Q��ύ��m����5��U+x��� ��VL���`��V#Hs�3j�(��K?�x��J���I}���B-谺��N?ؖ��U%M���/��~l��mH��W]�i`;��6jX�F�6��*��A��C��U�|TҀ:���@�/{�\D`� ���ueR`�-=�*�,�C��>�a�N���{�|O�`�$���O�歱:^��6�;W�&!
�J��[�D1a�ܺ���O�%��k�%�́)J�i9j ��O WP6�嶂����gY�Q��V��N�x9 z"�؉ؿ����Ѹ:"mF��F�W{�z�ϛ���{i��V�P���[o�u.f!�G/�|��>dzͰ8O�;`'�iN��!�۠��Q�g�.������SG"K�Pu�|�Nab��ļ�SU>�5l�ׇ�,�D��1pwy�т.A�չ?�Ν��4N�.?%�WbVӱn"��!�I�����e��!ޮ�h~'���x��s��h�.�)�`�g�A�щv���M3o���|���%��һ�͂h��t{�AF�z�� R�oK�"�=6S��ӳsY��sXQKqcP�u�\�熲�Ў�F�;?$S塎]z���>˿:�Qr>�y�C���~SeC�	��v�ك��D��Z�i��H昫�~�8��%��uŪv�A�����z2"9&^�5á٬���:n������m|��ʡ�uu�	�6��
��/��^<��T���A���Z�#.�g��=�Xg�\i���u����\�<vn%�X5�ӿ��:׍�0�Ĉ<qW�(���.�낞���m��Љ�<qC&�B�b��l���&��2�\h�ө����B4�B���
<V��n�ZER���٘�D#��� ��������5d�-[��?Mp���>�����.b�?��	?uo��w��{�#�t�Ѽ�?{�$�T��РG�Chd�m����D��ܮN�%��.? ]<�.�
����u���9�1{[�5pJ.Jk�c^kt�i���/�hf��/�q�!�x⅓��������ӱ[ɢ�(�U��j������2%.�٘/09�qf���]��q���8zO�߽@t��)�TX�#�vm �;�ti��Ll+2r%�l.륉��^�7}�"���P�<�x���ÃE�u�l�V���g�a��5�E!�)��Gݝ�&@��L!x�۪����#�J�ls����8���ėH���I(Y/ü�������ekK䦻���9<����6k���I��|#e���"W�>ѪGT�o��g̀M!Z���+o��Ӵ�1	��/�V��.�F�Q[תPk�A���6�����C$�:�@s��:�La4,Ņm��M���@q��xb��ɫ���W��������_M��a�^lh�`�Xg�x�1����Q�8��~�����(��9�/�s��mn��Zq�R.������8�0S䝏>�u�-GY%2���&B
��14wJ��L�ɢ�K�)�zHM �_+��'LI�Lė�H�G:=F����^,�i�����9h�p~��^Y��r{��_�y������s=RE�N��&X�<$w��S6�`�8�;�w���>�f�/I$��w�e�+hǐ��:g^���BQ�) *�"��K���r��p}R��%��SXTk�C�:�7@%�q��O"sX�X;U�On�`�cφ�I;����.^�?���Ԣ���c{��S{���<�_$:�y~��'�,3�+i���	[�ƭ���*�1%��5b�E&�Z��RI��ou]�R�x�i�a�n�kXS��ؠ z�r�\� �����y�$�Ԉ��׈�J6�[=W������{[ �;���ׇ&���o���ǖv#O(2|�������?��3��n���$X&�"\��T3���r��T.b���ԉu^���w'o���e�A���QƩw-ʕ(�*�qKm1�A�G����H�"B���U8�I�L���8�3"��/9�$'�c"���!?+:�t�����'�Nxm�nz6��n�1-�E�pbUq�� &���Z���QA�<�v�A��:�蔠ڶH�0OCl�j�>߇���;��F�`�`"�*�V������T��m�-:�
E�!�i��h�OEYA�*�l�Ipot�eG1Ʊ��tѸÿn>�*f��Q����� =;�f>~B���ar]�(�^|��Mh. ~?�'6Z"b�	3�i���*� �gQ��C�;Bo n�����M󶇴���3~$V���@2r�ѧ-�+��_e	�;�CH��Y
��n'��F��u��PV3�[�'�Mی�Fp��v�:gk�d�'�sI>�jl��G�傎�?�.�6�� �A������f�Qp$\��?�?�E�%g�IIT�TP�U�r�|�P,�Y�"x9�����:�y���Ykk�l+t"}@��l���+�w;i)j��Kk��H�KPV�KJ���%`������Z��&�LF [�"�罂E�x.���U:I�,�CY�-d0A���MoM"?���gҴ��Z��ͳ|'k����
������>��X��}����ơV�5�/r���*a:v�-�E�{�l�8 �Wj��IX�G$���K&�n?�*��Ow���O�PU���=$��w�%���qC�k��_�9c��q<�9Go28;b^���<n :a�
�מ �iYό�1��VWI�������^�kNR��?��(>Si�;��k�ѓ������6�y���E�1��a���6���2�U-:��m��1�N�{wN�f/�!>�]*�z;lH����'��D����Us�~<<YHL3��r1 *��B��,5׳�GG��rt	k^�rx���D�Q_qH�N��p��VA�dh�y`�l�`�@e]���{�;�6��8�/%����.��x���y\ݯ �en��/%����h�|�&�J����t'�� ��5S7v�6������zU|#�LjtA�uhБ����I#ъ�p�6��B숞��?�aZ��{�[<D��Mo�C�{��E���'��6j)i��z��[P����a��R$�#�� ����j�<�
���^q�U��Yx(� ��9�ݴ��'�t[ʫ��
b��참���d���61fk.���9�I�����U���M�~ӫ��Y���W��0�P(�� g�|bS����"ꀆ�(ZU��4�t�#߲�M�IǬ�m� �=D��u��=,�9їG��Ǽ��꾬���P�5��
V`J!DuhL��;�5i�eK5��^���o	�q.�kjo1\���8��|P��eJ���{!%���ǌj�a�Mj|�E�CD���64�������U��I�!az�'�4��U;��q ໆ����3��Y�rL�eP�Í�.��0lw����k|��q��l�tY< �5nL�1�����T�v��"��ˌ��\�O�]�KD���h�˜Q�n�@^��h�D\�㦽�g�>2#
p��ǩt�W�c���QhOt�!�>�"�S�2m_o$7}�r���~� ^�zNr��v�;oȟ�;h9���W�f��KZCʏ$�+(Mi�5
���S�����X�{��ư /I���r��ܭ2n���䖎5m�߽/I��`l�� �v� G��ू�D�Z�I�U��-�v�Č�ab �v[�̴�D�I��Iް�2�ث&UM̲6ՄFz�����{��>�?s�����0��4�2 �K��}Z^��Hf�#ѻ�����иGp�@���Ι�����`���gA���˭�3���D��B�y�I'�D��j1�:��
y�S�}N�[����ˏ�iٵpU��]rҤ�wӎS�����؛�ɈVz���;π��jdd?)��5����~*l�Qxg��@acd9�$�������scO��
�e�2��Y�������>�=Ҝead�<���� �{�����V^�٘,U�G�_~�w+ ������w#bGNT��|�!/�c�-{�roɦ`���ߘOμ�l>�V��-���v0U���H ��qd�����ډp��2�
R���|!c��Լ� fU�+zya�B,�wYL����t��;�J���0�c*�l��kݞ/lMI&�$\��\M��ܻ�e��7���w.}�ʢ�!�-�"s#�^���Szb2���j�X�Đ�^�7Z�����N]w7����Kԩ���_��O����������,T\#8��:qgY��j�R��WFl2�ISRx��`G��kƘ!�}2s�Q�/)O��g,Ms/1���aL��B*���Ӻ<2���rv�GًS$��Z�Z�d^�����o3%R�@О��%*x�I�#��D������ؑj��^��x�!xIB���s xg̐�C�� ���l���H�0���'���\s�xԌ�Y���09�eon��1��q2�,��¥sƄ2;���`c�cS��0}i�zĠ�J�R�kaO�x+�0l�V%z�-/��"�0����MC�DR!k��%H��-�y`2= E�M�D����ݐ�Cs?�zo̯��$P�����-^MalGke�C�����GT��/��_e���2ѳ$\:��6�BY�8�Xb����;�5��&�Ḭ'�0=V�Xf����e��EQ�[d����Q�$��2ܛK͓��iEM�:�X<���0��L�D����_Dv��?���������l		0	�f�}�
����yԏh�&]�;u���n�o��b֕4�Xo������(/���O>]m��ӫ�� Ό�/�cR�I�WB���j��jvZf&��j�z��_䟫4'Ӱ������~O�}���_/�ㇹ�4�����,�[d�	�u]U�2��)p!���L�T��u_w���H�Cj`�yN���N�Q�,'��%{��������Y�kE���T�QMa�?�^��0G��_)-�t����{�Tr\�9��ό8�������O���u5+�I��ْGܻ�0o���Hof���޲k��f�)���5OJ3{��ҟq�B�г��Zc,�>�=�`R�t[&Xg��(�����E�}���̭�Q?�I��Y@0����_5 m�[	�W%��L��W$�r�~/���ds���YK��C�}�nؼrm�1u�gp$�1�"�EV"a��q���5�>L�a�J �`\-����μ^��=X�ZF۽u�X��a/��[�V-|(����OZ.d�#p~VF&Z[PU��X��������A�-~m���	a�W�E����u@�R�~��i'���u���@�$��=�}YA�2�S��'��(7G[�MT*��3����g[#�Ku���\�mw>�a�Ms�~ ��e��GA�:D�7�@���НS'U�Ɠ�x�s�R�6�1���%Ϙ@`	adŋv1�t�J/h:Y���7�3�	����Tڹi�_X3��-���B[+nń�����;FegT^�'��$J�=����-3�5'���A�0����wrN�H1��6���No�	�d���c[�D�B����tP���4�s~�]�H?�[`��._��+K��=c_Lő�)�\&N�1R:>_��%�����R�k昗�Hڂ[,K� �Ǟ�v����Q�nX݌Fbs�ۑ���W'P�։n)�����)'/��"P\���Q)�����#i˩�6�QC�m��p��_���F��s�u�w����NXF&����7���_�U_a �%y� xf�M�$�8%̔�q�X��e'�H��h�aZ��R�G�{O��@�m���ڣPc��UC����k��p��Dy�n�V�q$w=�&�7 �l�m>	�K��z�����?�Yǎi $%<��5��=^�gt/!�s