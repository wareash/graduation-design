��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e����d���f{��@����S��>���4{��ת�AO�Q{���Ya�uɨ92!�}�TS��� �5&���5B;����tB���z�7q/��1=�5?���J��"�۝qp���Է�E8(
��$�v���c�˟&�A�[OJðd>떍� {qw`��J?���P�6���}�%�;az��n<��6�����T��7�8E���娗�c����x�;�x]P��ĳ�s��\��^9ȻZ!���d�&��/p����QY��7��P>WN�a}�p�W�&y�g�B���~�B']T
�q7¼vR�RZ��R�J�n����¥T�ѿ��4Y|R��J�`�Eԍ�#����yv%
=�e���
}��B�eһ�	;�U�p�B�P>o����=z���/�g�����4<+���(�/�NW+��cζȬ?S�"p k�2����aFyȯYl����������D���E��I`��WXa���	�nP�X�8�W���GeV�1���y�h��]ݝ���ay}�C���XB;���ឭ�z.�^��0CUVJ@�TH��F��#��2��%�W�]b�R�*�"ó%}����j 
_�����OM��E��F"k7ϩ8�r��t�8���=Th������(Q� ��KG��{�~���u���ۨ�.9�����:�]��ߐgB)�k=�$�v>|ʓ�Gs;�O��F�nYb�d�"ԉ._���Ȫ���(Zd�����KZ��ox��*Q`���:tU���:�*W�(�sX�Us�I��l���:|�;��z���^���'�ȋ�����]��<�l|\U���v&�Y�JFW��&o�<��
���^�G�{SdJ�'������kxs���f�\X_M"c��0��U�����r��в<̢D�E�<N�y-*j��K�v��Ɉ�s�e�x�>l��*����@� d�!��q�ѨP4 O�J�|%�]��%iM�M�]/��%;+�+��3�'�#��b9��i;j0H87l��]�\ё"-pD"���:1o���0�&��B�
���>7�B��z��e�ca�!w����W��ACYFH��P�"Vn �{8�۞���ʰ�%kJ�Ӄ��"M��$p#^���l@�	e鱯�g�>�>�%���[%3�8��+��s]�� o!>g\z��9�N^�S�_C �C2݄B�E�"��Ǌ���?���RV@
�v��O̬�IIk��N��(z��"�U1"�8��Q��7���KM ���QPG���e4�}�Qi�����#EA�yK���z�Q#v���|L�M0����#7Ѽ-
�}��~�Ad���c��j�ab<��K�,@�l��l�	N�C�_�b��*��Lv'/!Zn����Ń�2�h�_b6���+ʗw���cӺc&k7�Q��}J���ܬ�7��DB��Zu��]��qcڦ��wbO<�{�����NDݗZ�h\ �� 5I�0=A|��כ���|�{�:+��P^QIJ�P	����ƀ��v���<A�`p������Z�#��xu��	��n�L���G����r提��ʆ�a�!��+��~g�s�}���>>�u�z��;J3?�3��XF�i�:��&0N���$��]8DJrHK��ŬSZ$^b�P,�{�}B�d��gy�����Szs�hipc�_�$���i��hߘ5�WJ5��=^8���ȑ�g��(#�$�9IU�%�[)*�Ys���^�k�m��:ܒ׾b��@�>�*nt�k�I7ϴz9�y��$K�j��V�N�\�M`�ME��W8��H܋��6Oj�g�������L�nn���]g:���d��:�Bm b	�v-x�S5]OB>�Q��훽i�p�(֛���.t�g=����~Je����Wl>ٔ�	aͿ(T4���p��	R+��Ŗ�@��4��)�~��M%��,�^G^�m�<��k�~�d�R���G����F����]�#�Ԝ���-�A��6Ϛ��z2S��u�&b�8q��Ÿ�
-�-�`�=H�r��O�)\_W��Q|^������j��n	���Un��/7�D��(�W�+���1���	��͙��M3#sLN_�D# B����B������JgϘ���#C���\6�hޗ3O,{�D̪c��.+J�,�&(]�m*�A��%�֙S����o��hE�=E�>]���p�\���y'j%�J~{J0�}�ز��m�ty�]M=k��`�����Z6)_��E�'��"W?��p|$���^�߸e���ej�c	)�:�r\�&�=A�d��HS��s�E'}\���Y)B/�����vd�7�n[ޢ#��~V��ըC�%��Xb�Y1����HX��c+�M쵬g�ne\�(U`.*�����':+�J���r����ǎL���zy��g9At���M���3���[$��G&!��ƍD��RD���F��=_�S\���KU�"�X{����.B0&�~�`K�!�䩁������ ��y��W�@��Lb3C�Y�@"T��>�'2��F�?K�#EExQ6F�lg�w�ݡf�wD�7���)
u�o�/'�i�O
�O��L+i�R� lL@��6RyXjc�iV"���a�˖[2��eG-,�<��vys@{�X5-�[����{D�Wq�3�E��焧��jO�#5_�֘il�|�Qu�F�I��Q�'���~���O`4x��al�$�E?�SW��Ȭ�Y�(P��''採 ��p� ?q�	*�b�cnuf��Ҭx�2F���!����HղC?&�`J�B»��������{���(�[L��1�����������[^7&I�|�0�b��ë�B-Wa��<%��|�K���9��;R�7�A�v{��l��nH:_���;��ɁC;3���6�P��U�9��5������5��2�{4��)�y~Ct��ғP�����P�(�q�q[���o��S���鶄�pIo�t6�c�Pg;���癞RQ�`�\�Y�.t���O�}kHmQ�r��v���UL��W\�R�%��"�@����4g���u��B�{@����jW���@��2�)�/� ��"��3H2�|�B���܉Ў:a7�}�2�寫���&��[y�W��ċ-���͆�%��*,�cL�h� �G�P#�yR�L{�hb�.���;�B�O��d����
AV#0�k��[D˔@���K�?����f�g5�,�������L\����ѓ�5G3���N��:�I�4��>!u�'d��rJ+Ǚr�ɱ�����!��Qa��q'
�`�dw��uW�$��=��0�u~�O�ڐu3W��FB꒵?C��y���8EX�'0�ފ������]�m�c_�&
EFv�uU�u��Ь�?@�m�/�E��Z��}���<@8.j�x�?��i.gy�LH䟂�wH)ч��9�qM���T�l��Q	��
P~{�����%�R�N��3��`忸���(5�� �)TUfE *�dHN�^Ȧ���P���]�ZIs�Oj�@M�I-8GR�Q���N�OѨLu[�f,��6�}=];l9�ӵG^��Ç�v�GZ^�{d{���e��k`�Eһw�U�X��=)��v������i�/xa��o���m:,��pq� Ū��c�rL>��,�u�Z�e��	)��X��|3��p�+!� �˖̩⥣�<��:�m�B���r����Z>�� ��� ��ڌ��o,�'�O̙�2kG���F�V4��J?g9X��0�4������?��P��h��$�N,�QKFE"*���3�䷮�{���UK{M9B��h��K\�'4.-��W(��x�n�d2I�9!b��]��b��O�o2	��Qz��?:o0^����IH�b
ؚ����!"�IF�Uo~�iM�Um��ۘǭ�s<K��[xp T�Z�:X���.|��\��\��CA�Ջ?�����m�<f�pN�������������a���E����o
��~��$W��Z)�*Ɇof0�TK8t{Z+cy����pV�cDh;���4�ci�7Yj�y�� ���Ɠ^F����2Y	k�~��������\sU�:EG"�n Ҙ3��+6l�5�V[��	+T���5�tF��7���?P'�>�����w�(ui3^ޜC�ŏ5i?�ZA j$S�M���B�~���m#��h�"�^E�3�]�s��ѝP��]2~��W��qxxj���d��vr�'����I�}5源P�����%Ϻ�s�?^y�i(T��ZƔ�|v���(�&㏋�>:�pm�k��n�]��~�5V��
���/�إ��:	�K����Z0 �R;�0�@I��F[�1�U�Yj�J�ɜ/Y*��)���,H8/nU���{�1��:�"��+>�ἲʹ|����m�߄�?�:	�Y�m��d^����C@��𹠜�3��F��iҔ�N�G���B���`` �<x��y�m��B�q�b�Oܞb��t*L���V:��^��Bܔ�o��U�1�}�*�A��������]=[�u�]Ƞ�4 ������+,�P�x.�}�y~ ˯�l��jF��Ouu8L5A���0�Σ���g���TP8�6��r�$�3��^�Q2����V7����c��B�.���w3"��6�-{g����UPr&��B�`#�l�Lk����v�v-v��홏�D*e:

�rk�}(�"a��1ו�9}��z�d��AGݘ;8p�@��A&�?��*2���ȫ�& j���y��ن��ĝ넥��0��E;ӧ@D3�];�O���[�jT��2�8�Cl��p�%��u�a�q�E3�lԦ��T��~�=��D�%Z������3뮪L�(3Z������ɶ|��́��[hy6�;�䇫���������� N���䞮y|��,�k�e�<��D��4(y�:{Yћ�:���Ew(7�ˌ0��]TK]Ӏ�OH��4"��$�-�Ҋe� �;���&���%�.qv���$}idFX���dP��>�M�'�+d]|�0ꚲ�d�}?eX������
��(%����묵Z���ݡ��ޠ��������C,N�}bA˰�^�s(bN��3R���y��x��Lޚ�/Y��Oe� �[�乚"��e��9�)����?����h$1[ʛ��e��A�V�rs|�&'<�U�e{�g�J�9�,:.v��5J6����O	ϋo�+q�`tJ	ٮ������f� �YꙀ�`��t��L�U�DYLGȜ�kL8Ũ�z��_$���fvp����C�7hX	��7HO��#��\�9��nf0$qJ{�J��Pr��_p�}L@8�*���$ƁO��Nxqi�3�*��$��? ���"�2��|� Q�^�[��.5J�$ʱ�k؍�$k^��~�d�ǇKI�gA�LXN���T�t(�0w%��_(\�i�͹@Cn琋9��7N�J�Z��m�%�袘��\��CL�I����wK�V��=pu
a
�ݨ��{@���a��=q���<P�[������O�xu,��3���A��US�L
f ?GFV�����V{wCh�ޯ�K��2Uc�U9�M�j6W���]���'�����G���Ӆ�����,WuL6��D$s�^��4��A6�!�`�Y ������}ӠF��%�SA�]���(��ybL�r�� �����˟�T@3��
����j��p-����L��zQx��
�z���_�R��֬�@�]����&��=!ъ����;*S%DH�l�P�]���B�MV u^!���Zo���8�R1�( �ߩ|��� ��pb���H�׀�T�yФW�h��<�[VB����ctqZF��#IQ�f��Y$��:��J[��p��������{�����mg�[�xr��!������P�W��&(�hڮ��SݏJB�o�=P��(�˘1|�q ���Ju��1�r �]DZ���y�Շɶ���]蓧߬���k3�zc3�x=��/�������.ϴ7��c�6�}Q�����a�%�}�Ii�+?\!nT���5p�.��8��M8בu��q�L��~��Ш&-�MX���Rĵ4W��]+��s
��G=�;G<��7