��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jåا{�\�u�?߷�dn@6�zf��r������;�&��0"�*hT~�79�{�7zlC��ኡ>�(N��4�?5�#�M䞧|��G�[>�H��y���W�3�+���`n��pܐ�1�s�A�r��y�K`
�.����U��?(�GO�����Xl\�s!Ԭ�0��6W��8�u�2���L�D/d�句��X�#:�z6r}br��0���#~�%O�+z_&'���/UT����Y��bc���j���8Xz%��r�LLH��'��̃lx4M��J�d�q�qa��	K�7�嫐�à&���̕n}�bm��Vܣt�2t;Д�5����Ux��X���%���e��g��u�B(�\R���
�9��*I��[��{�2����|p���f��5���}�H�d�/�C��h����mcd�����d�ʒom�ȳ�m�a��<��#�П�_�,����8/ş�A��=�Z�a����\�V�z|�
֧?��Q1��H�>^Qf���H(���T��8x�K{6C(N���V�ɖz�en��6�u��R��c�����|Ot�c\���R!����m�Ϡ���Y��5ӿF�� P\����B�Y�׳e�|6\q$�҅ID���b�Y���łY�11�a[�4�c�8p��Bݴ�ǲT���k�l.6���p�.]� �x��vh�̂)�5%Dnlù$��[�ځ;�)x���`7!��%�(�<��Y�r���5��й�[HY��L���=�1D䡤b}?����ST�.E�k��龜�zh$r9�^��� ø�ݚ�yxI����6>��l^)dhj�v�dDΠ��d�ж�m��s���1XJ�_ǽ�D�a+c���;NS�Q���
���Bz����8��U13Dj>��E9�/a���i���Q W����Ň���eg$��^��Uj P"�F�f,��:ޖ�24pk�Y�<�����i�鯕�WH�GY����:; �b�o���Ǔ��9���Rƹ!�
Ue�6�&Q��߈/����Jb4���a6�|��Εn�iW��&q��B&���������Ʃ���L�}K�@KkJ")��&2��\�D�2���ޣ���z{�m����n��0Z*q���H������?��+�C	ɱ`�\v�'���D�mc�TP6�{��$����X�,n��
���?���Qv
{r��l�#WhKT0�Z��0�G투���*%�L�Sx����Y��,��vK��E$�Yl�e�/���Cad~�m�gD�	hr<��w鸕@��F��:Kt�-�]:JP���оV�E�Y���3���2W���{���1_H��7�ԓVx���N�9�i���b��L�J�!�8�z���?�f3QJd���M$E/��Dy���v���($~
=�4�Y�с�޶�r,�8%~R�:m*��8~J�;�Eo��y�=5�_F,{��|�b�rzZ4�.N4TG�ȹ_�{|��և 	+uì���x�l���]���(GY�dm@I�[�TB��gVu�<�z-US�m����K(�� -)��g��!��]F>��d���;&bb����h�ה����U)�����|g�@3A6��JqX���i<z�)��l��$vu��!jђ����-̙#�!|j$f��<�f�{?�kڊ�Ȱ|�[U�� r:��X:؈�Y���wvgP^ٽan��g���)秊��"Y ۸��7PJ�d�Ԗ(�z���l�՟����zM\鍼ox����+�0�����VH(�3�x���]�U?����E��<�;z�X�[��LYe��/��5��E鴕�w���0�u�a�ޯ3q;�/���2m���tX�������,�sC��!pgW�#+�b����8y����/��2g�Q�Y����W���|6�k��8"�o�����pjD9�J!��)=3�񺟲�r7:�G����/���* #W6Ѯ�N���7͎EК��/Ik"6u�O������Ӣ�+�ɂ� M<��"��͝���7��.{m�9��!�m�M��@`ቹ�M��B��N�ʓ�jS�l؇�\7�q�~^q,��ްҩ�  }F���.�H(����m��y._�)}�ىSla��bE��ˮ
�T�\�K{�<�9"��Z�	N�Si;"B&�O���<t/�wP 0@|
��{e���o/�'�7o+C�v��T��a�
�����U70�\ΰ����wj;�HQ��(�g�g`H�v����z��~pl|'�OC��rC*��XO�ފ1�Ձb�B�i�Q��UǴ������2� �4����_��P�`�����O�>Te>�Nj�C̷�S��+�����L�/6����F㔮��,DV#�)B�ʇ����ț�9�B� ��eFT#��ƳP�� �|�;�o����啊7�$I�j��I���̐�r�"7�gH�uc6�WmY096��19��et�g~V�pC��K�*uOr�~q������ȳ��حV���k��1n%�9�$ҟ�r4�R�#+u1fR�I�aO{-	�E�Tf7*N�+��C�:��
��r*7Ey�C�J���Rv�76�%���Rc��Q�\�S壉ɚLܡ�9���ٞ�b".E�V�Lk44j#��%���<p�Y��>&Y���(�/Q'��Y����&o��D:�l1��.��$驿ʨ7˰���c��E���Q$Y9Ǧ��O"V�0)�vD3T1hݤ'��i_�@�L;ǵ-���c�U���NS*Q�5v�#�����%y�$ó�&����Kn��n�o˯�Y�,�W���:᡼�!��oCv�1W�zĨKx����o��:��f/U^�iw=��Y�j�tAi�A�Om1��ʕ8چ;�Dk��Y���
���;J���
m:5ߡNM�5�����N|��A��9-����j�W��ZAa����H�Jw��v�0��X:��-��Hۦ���C����rGk8�1�v���z��A���W�l(��\���k��oL��Uק�)���(pf� Q�N��j;/������9,1K���Z����n���9�Mg9���W�T��M��!�r��	���G��]�V�}�I:K�/�ڎ����fҁ�d�0E��F���wd�5"����ñ`yH�]۞Q�X\�^�W����m#��\4˰�ʌ)�Q�x.��+ �JX�b�X��z��/&<zt�yg\�2w�m�%��Ռ�?��0���Ű�
���Xf�R�͋�>�ǂ���+3���#��dZ8�_��|R iڨֱ��&�����Z��I�����ż@���J�����N�}���O#��f�~l�+��s�����|������QRY\h�a���[�I�>~�)�ؾ�׳w�[;ș��+��7�&c�P�\��� }�ބ�YF�6�w:�Y?2�rxYW�����>&*��bX����^�$V���G�����(��Q��Nt�%�Cbef�!2��֙�&K-�ew��l����>�tI����p�e� ��@.3���E�C���g�/~��;ۼ�U�.x��ڷ�93a�ǰ�+ɂ��f���I���Jx�G�Yp��`����zB�oKg&v-��-�� �͟TV�ۢ�V�X�F�/�[��Yx����/�sr�g�Nv�ţ�ܚL��*4����Ũ�&��I��h�Ī�x�� ��')�p/���ȡ���6��(!f�LE�kƕ�|�1ݢ^���6?���/k� u��9/`Uʭ�+rt��4ƫe��T^˷rQ� ̞�x�ϴTO�_����+�S���E*��'W&���rD,O�S�CG^��⏻z���� {7�Ŝ�l�	u����>vٚ�*4sO|�����������Fs����s'��;���Dބ#7�횩4�&��R #�)��q�5+�����~	X�Vt��hsj�sOܡ��(�V	V�C��}�7�y��f�ΕP��+�@�I&�<��3Dm_�8ƻ̰�I,җ��Mx���Ƃ\��H�̚��*!��"����y���k�؆{�?��f(!>XN�)oL��zև\���L�h=�����Ibl�;I���6��[?ꞛ+x'��[�����j��u����C�U��T҅,��n�YI�$�Ʋ�{�3��D���4ʞ�o�FǾ���e7�T�x��[3�}}�-w/�_��P��[����;�\���9�(�d7�c|��d���Ai��zV#-���VXG��Z�-�0��F���t���f�l�m����>/w�E�ױ�<�79�	nR����	������\'%��"Ȟ3 �m�>p0kw��Pq܋�1�.��b��J��Op�(�)kK�ĞQ��L�ڲ��ݍ+9*�:f��K�S/��٩vG��~đ�\��
�?5��vK�<�<�����7KyE�|x�m�a,$����LJ����m��[]�;|>}MPu��Y����0�_�T܎��[��$������D��m�o7#M긲�w�biq�v�e�%~�/�</�>4�[mLĺ��^/���j"9����ZmR46tv~a�(���&覀j��5�b��tݐ/�7T�!��ʝ|۾����u����8��XhV�$�	���*Y?j�B�my����Օd���.��&����|�S�\�5D�2�s����Y<틎a�E��7��k�o�)&��@^R�6�	I�ޗ��%�F��O������*�	�t���s �U�Y�	�����Z�8�˅*������R��.j=�XZ:J�([(�ex�U|���!�:�M�%��
|Y��#^7O3t_��D�k��w��u��IN���s\�,��x��}���}:v���Z��|#��/�f'�\[]��VW�8�66/�v9xgHD8��p�<D�o��Q���Y^�>��ɥ\
}L���!
X	`l1ĶަΙ�Y3���`��3�F��Wz��2����8���4�W�.Z�P[W(���Zj�<y�=���+Gu�6�l_@U0L����uɶl)��[`��3����DɍuIȃu�j��)[�hj|%�G�2z�H�����B��|�z�2�K���=\DK�����4j�Y]���i=[�ؤ�3�3��ݸ���k<�!J�&�؞�U�û����$(�r+�|���Z�u��s�<ډ���+¶>�2��S��uFfb$��<m�w�l&D��,�"՟1A�9�)3"�^!j���zM�@2!��o��X��;�(�D\�����#��!�<'�27�/��][Alo��pg)3��r+K��#��u]�Ϝ�=ś#�W�9ǿ*���i����ʇ��8����.��ӻ��	��Dӱ����W+{�L�HNT5�p���]䲲��5��>�H-\�6RF���7����]�]Z�p�)�jg��F�$��ʰ���TDv	�]�>�H���hVS@������=��j5�*�ewd���#�/�\�h�z����7.��Mc���R=vx���N�@֍x�H�x�1��
���7ԭv��%-�	g��*Y�p� ;m{�'jޢn�a1���cv���dK�w�ϰA�3h}�5W�YF�����/�lKh�<G�y��Y2���5�"�!���X&
�����A: �G5n �j2�U����� )�H��i/�N����q��Ԏ�3s=y��<C:���Aus�Ţ&H�<܍^��&I�?&����6'Da�-Uiʚ*�י]3������i��[����q�4�j����ӻ�0��f� �J�������I���%{�� �:�(�@���T-+�f�?Ԣ�K=�^ewatx%�g%���5���/��S��e9�^O��������h�!)��7`�6e�����saE5�J�!�Se_Ԃ�)�g-wX��� (�����L��s"����e��Vf��΅���&�:�kLr!���6�46IHWX��#L�|�C'	��}]������%i�M�4E�~F{�=�Gv��VZ�i�)�n9�cbV.��������k;��Rzt�Ʉ�N�y/V}���u23ڝ��9��1�D�ac�t��'1:�,RYt0ٖnvIu�Jc���H���{�����5�AL(t�YR�7u��OHV�=�?���"PI��/�� X���R�L���@ QIz*�%�!�����7��_f2����$�4\�v��6?<B�ZkXlԣs���CL�b��-m�'���M#QϮu�;�w�&6`�z%+�IG`^��޷w�Z�R}?[a������u�8>S��h����c_ܩ��Wy����ɾVTm 3Q#�Wwf\� �K׶�Y6$�(2�1+�3{>:R�c'!��SMNs�s{~SA(�!���F5�Wq}���Z�	�S_�@��iW��I�[`gw�DR^��ֲ4���P�,�����W3�.�z�3�ZEq7̙�\L������P������*
B=v{o>��w�B����/��a��i��A�ʪ:W���*biO�G����DX|S|���iY��z3��v؂�l���݅�86��N��������� ��>�C֬Ը^����[�m��)]ܓ��_X��r-:/1}�؟T�@(T�j��F$�����׷b!�� =�3@���0��xm:�J��Y�dej�GV&}�9d@�[��ͧ�x{ ��)����v8�V=P���ϝ"3�
ͺSt.�[���~��U�	8���;sy?4��w���B�XEV:'�����<��Và16�l��gDKd���Tz�6v�ѐ��C�,�r��jb{X`����?�7�N����?��B�׳��h����P��ͱ��(O�O�M�����.�p����\�S�-�{�w�e�f����=��A
O��r�Da��BriIҬx���
�Ri�^�o�È%��\���\ĺ�I(��r+�z6y�GcP��� �!�?��,p�'f"5Ϥ��4Z������R�с��&����,x�\��u�FAE��<�-,�A�o[y��R�'���{����`�Z����b�8c�^qƋ|s�ǠZ�LJ��a��f�W馤/�Z<LH`D�\TW��U�h���B�4O'�nDTG>�������/�\�*�v�ھ*�:���vG=��<4�#B�ZNM_{?�VJ��g��?a> r�<p���QCs���k�L澍�ӗ�e�x�^a�.�t�Rr�F�b��O��	�$y�,ME��}c$"�# ^�^%˭��?����[����,#�������*��e6�	d�F&�wV�&�伿��Vs����'�nZZ�n�R��c�����Rϲ���6nV�U��`��.B��y�.��?���Or~�w�����25�@k������&�p�X���{�l0�@��e��A��4�o.:��:+��ш6p�Y�Zi��ϖ֣�cһ%j����_�jޜP�~��T�/�����:�{Ŏr�DEE�2S��S38Z�����Qju���:��R�8^9N�#E�%]W&����3������B�B٣xA������D�IH�&��G��-���6�wm�0��r�I1)b��>���������o�Ѫ5�����w,d�$mʣ(�(�V���o��1�STS�Kiޤ�������ݠ��I9r���e#��<%7w��� �A�U?�O�kڈ@t%�+\1�4��ͨ�ô	oc��F5�j1�>%G�|��$��*8#��x��pށ�'p9~~C?y��Ч3��NUj����)��-.�&�߿�¾A70l$�^7�f���$V#a�_n�<���0�0{˨����#���m�n�-��U�!
�X�(�=�a���Gf�ZjX���{�X��ݮ��� Hzu���o�Z���&/�%�Oʣ�����+B_*�]6�]��'LN�!5��@�P�An���uz�O�6C�sz�DXf�+���eڞ�K=h�r/�`�ÀIr��	��\ω��.\�CD�,x�p�=('xlꗝ�e�G� ��8ة�h�t�~�ɼ��\�o�?�:��L�*م�:?_Y����5��5��9�	8>ʠ�c~fC����!�6��v\�Z�4$M&b�"sd}�86�؍�>R/l�F�N`���nMuˁ<,�+��#���#"�+�9�5��
x%�:��8ڍ�v�z�Ǿ�w�DJ��tO���3:�5 ?Ug��d�U���m����h^�f��l�|�+j�J��;���g��!�rq��~��ǻ��I�>�d�3�ks�o�
}a=8&�?�<F���S�d;��;ƾH�����&u?Gܤ�"�=_�[V -�����?��������O�4�&]'�C<�O�kIX�7���������T_�ۯk��8x~X{t��<kG3u�]��.��P��AW��ÛHK���P�l}>=�;oK��s�Dt���>IL:�z�Z�;�"*��9��*�������i#pΦ���Q�����E:�v1K��AfLJ´���|a�Ֆ��Ae@�a5a]y���p��.o���z8*��M{Z=D�}�>[����2�G���cv �-�2�����5�{bQ:��A�1!=�Y��#����?W@��d���]M����]6;���>�}��k��8���u��o(h?�/O���Kt
E*�X���4%}�qK�0�\R�����'�4��y���|�ld�7� 5���z~�or��cL��/|o�tL�Kh�oP ����$H�qrܵ�[	"p����}�(�N.p*#&�y]WP�xQ!�큝z�'M�j��*m��� ���P!d��_������*��^��)�s��˪�(�H{(=F�F��jx��.C��#ƪ��l��#�Gn0����Z�'�b���n��������H�c�O�0��3�h�d��������w��>���O�Hf�®G�BsT�cv�80CLL�XR7��8�@$�T]�ю_��3'�m�c�� G�c}�(�Z�=��$o�*�����EӒ���K������>{3�|s;����z���[��[��m��K��h@޿��)�������jφY^��<��D��6��d�O�*�����(�-i��vѰJ��-J�&LȀ�?w=v*p�d#
~17��mHqR�P\nK}Pl���	�X�߱��y06����/D��X�L]g��N��:�,����������)؂�������־s	S��k�82�Zp�y(�T�C`�&[���ထ����sX��dK��_=��w9脚fI���F¯�.-��k^�;��XU���,F�^�R޵Ө����'��Vw���������g"�R���-8��϶*��Fe���xǄ
�#��q(�_�q�1[)��� }87���`�1'�v�>�+J��P��s��b���f#������8Įu�?ci��`k:����S栕���5���g�{�o�y�	oi��:U�4`wPZy��A/���	`?�t8�z~pCf�)�+�m�ܳ|�^;O��8���h��;��Ma����kL�,�W<���Ŀ&Fe)O����\U[/�4��H���2��Gw�5��>�<���Ę��\L2H��G�{@���:qb&z�Q����9,�ȐWA����S
O��L~�Z=(�Q�i��|�U���Ո@䳁���^�!Ǵ��Fϕ�kS�m��?���Q�[�4�}.��iz�:��/z�\�~;a-������^X�L��:�ѧ|�\$^qc�fm��S�w;V�q��%<FHy4���F�����l*������oz��c��������+֥��dF-�'�M�T_��p��Ã�yv����P*�͹�*z��'����$2�v���t�M�K9"�?ʤ���].R��ً�fM�#Eg&�bQ@d�V"��,�t�����j�7q�ꤜ�q��_����-�b�@�Z0��'(=����	ba�3��AL�c��{pd�a���Gk���b�=6�N�L�R�a.l�Ov�^�� ���FcF�z�-��&�ӕNB�˩i� ��Y���ҕ�S�P⽦�
��|�z�$,�⻂b��r�8�S�e��w��-/�q�ä���$~�q��㠔7��y�b�Sv��d��h�j�\ܞ�m�}�gz����ss����w*�*}�e���A���S䅼���O��x��z�$f97Y�w�M���������0
j�*y50����V8��zzq3�FJ���]�|�wr/�{���\\ѝ@�:V�>�&���m:|��5�H���1�m2�1�&�hUD�)cJh�E4���Z�7z���`����P��I,e���ͅя3!*e��S��K�<���+B.�ڐ��=@ڶ�x�p�޳k�����"1��T?~��Q)�[�se�WQ2��F��������L�B�"���!�$�E�I��<ؕ�{[����cV_�/V�^��-L������߽��۶�K7�g�\@j.<]<8����Txcxw��y~�$������ă�g	�G����B;g��ow?V��L�w�
�S*Ո�
`m
h��]�P7�5x,�A�Z�:�7B�f��$G]^�\�����We��ژ�=�L���ҩ��~���a{RQu��<^TnpQx��kIb�Tf���K��a��#��|�<ٙ%��}>C'u�*}��n�m�=��Nak$ȊX�N	�׸ ���bA� ��4��q���q���]�!�ae�n-2�����y��$z���G����P���-���6-f�w2{�����,gr7�j���bOC�`>��m����G�����L<��3@�� ��s�X�&�΂�\$biʒt�@��PH�� C��0\{z�6?�)D�ԉM�*N������,�c���.�P�E8�:�7��>.g%6��a@��oH�V���X�7�J+�� �8�(u���G�i������V�:�$ov�U]�:�H�wBq4;�?E�y3�A�Cm�61F���P��s��ʗ�����'x���˅	v��?P"/-�?=��<���J�s��� d[p�r�}]�~D⨷����9K�bŖU�so��z�҄���
]ݾQR�� RI�]�5�︓��}��J9��7�yh�����[6O��!\8\��a�2�����\����1&Τ�#x���* -��@�]��n����[q#p��އk�s=֒ꤸ�m�,ņ��/�pނ���s����`&�X��6m��X.p�F�PI�$��z�������\ބ1�mn�"��(�b��&}��d���-7	����\�����8U͹@� ��oJ���[�w��ҐsڋX
挶�B�NGfM�;���̈́/�F�Sx����@��ڍ�&5��
�;�F�q�����jT���b�43�u3�N8G�;����k0$#�� |L9�H�u�}��g9v�9��I����3U��.K���`U�:Dإ��f=I���j��yҢ�[�g�-
���]��Zx�{��"�|��%6R��Fs3��j�4'�Í8��-�#Յ�V';�4"�0h=�`
���()�,'�!����+�o�ʻe*�X:4
j��@����
�ZVS���5�7J׷o>�9�ś2�D��L@�N�;A[�����^RqvC�$���wP�Ǆ�3�4a+�!7x����I�'#J�V��[ܻ$y�{v����l�[�4�e�:ݝ��詃`�@�0=C�?rAǔ�����Nw�$.QS�E��srsV��:X?f�r��F	�+��L�����O�f�b��z�RK.[���N�#1�&�s�tJ��X�ml3+�X�K8����R�d5i��zP~H�}i�֯Z�oPoJ	����&��x��Ct��ޗ��iO��,K���KN�0�����3� �W�.�[��B�ϣ����@�C��k���|Fy�Q,�ꮬ}	�HM�6�4������<*62�����rU2��zWT%�g a���33�KG�]V��}�7��"U�^dwObĒ�s~k�1�� Y9�7^8�|��I���!�hJ:�ϵfn�c��;��B�aS��U�<.hwE쪰���&���N�Q �&�XV��Y��P�[�S�}7y���v��I���-%�&�J�R�$�[ ��bJ��@ZP�G� ��s�}� �ye���c~�nC���N?(���5�%�t���̓V��"8��f���&����\�I>9�k�,�2�{��J���g �"�4*�;�nr��[j��Z?�d�,{*I�����\��b � J3]���+_�*$�6�by�'2l�2��yr;H������Oю����pO9}��\FS���+[�X��a���`=��ŕ>I����k�3���0F}���B��{FY�.H w`&���L� �8g��8d�b|����`W����Z��拜����������%8�)p!X��7���f�W9�ͻ��V�JM�)�Rr�1��wb�sݤ��@_L/�4Ugx«��lOP��5ђǼH��N���m'��%�W��N��O:���B��X��)2s�d��x�/�$>��͇o��b1L��X��#&}���-r{1�܉#��zT)���뵏�X�/���'�����ݼb_�����ujY�](�x�lM�I]��Go�M#c��3 ��=�7�nm�Y��6�S������ګ0/
|��f��$"�ȗ�!�j���>䩩����`s������U�_,c/[ڒ��/75�M��qe����e�D��������cZ�e�tc���<���
 ��T��,�}].�ŀ���� t�Sr�7|��[�-��+C����-��bRXz�b���Ϝ,i��]�Hyg@���)�x����A=%��G
t��"
)�R�ԜP��8hv��2�E��vP�E�)SŊ�m������nҥ��}[@
* �R]��jb��m[��s��Z�!�fo�U%�g�_^ߚu�� ��*����-�grwc�遢\�6y쑸_xyx�r��N=g���{�U���֍0̎%�䝂��'�\�7�Sr�7�9������K�~�!rjQ��m�v���K�q`�V��z0�4N����W�L͋�]���h�m ��������)� �ձF�3���[i�Xb��|~� ��[�_��{%���	K?��w���Ƶ~�G�1��Ax�L��ח�嗼>�_P��~/�%��2��=�M�f�̀�Y�{ɷ>Ao����
Ge�nʉ��96�Q��(�0�ˢ.ɋFu����5k��VI�����x�����%�{W���s5���b�ue�ʘ�g����3���@_��p¬m!����Z�ꊲ�+s�3�֌�Ġ�9SG�$ab�-b6s{{u.ꪭx-S��l��=�JQ3j��z?�t7��=�N7���T5��O
 ~W�}\�!Q剃��;�$������'R��H�U����\�b�?z����X�B�;�*j�8��j���?��	�DY������~/�ˬ(ݧ��"XW�}]v��TMl��%cV��=���1����A{� �\�@�$0����}���.�	38O�_����}�Q�b� ��R)�ׅ���q�2t��%.�l_�9*go!"�����5��❪w�P5A@�>�>o�Y��Z��D������
���Z'�����y:�*���x�_�$�m�Q?����9�!,�����#��H�T�pz�"SK��^���*�$���ף�z-O��
ycqMɢ��U7Bv[�1>�~���GMJv";�`7�@���'���V� Ѯ�(����	#.<�퐱��Hh]����Yb���{���II�>�Ӑuq��}���@;�&�oӟ�0w�񥸜�m{� /��h,�n]���-������Ȅ��z�P b�������4/z"%V����Ϙ��C��35�A�_�}}BO���n������ɩ�9����j�Z�7�&�I�۬4`��$���8��%�ʏz�6���ݞ�����{:��2f�7x�1�Q��p������>�M0Y��7Y w�*
I��[�֬��u�����%������A����� ���#b(�B\�\��is�/��.l`��ZK����]-�P]W�����8�k��Z�
���A�IU��B+e�X��|��^�Uݨ�zL��@5ˁQ���x{U�z���?�~��?�2w��]��u��Z��Ɉ�g�������bn�J����B�Ĕ��z@��[.'�֗��f52�R�h�g�wȖr�j�`�`OB���(�a�G��X)P��9�LR�����)M5���r�)a��A �5�*��[��荿,L.G(��|�Ŭ�0�bsi����T>#!�T��ʀ@��ѬLA�o��'W8~����n�D{���	�:�;$h�@8��l\��=�#gT���{U���G�->���$��*?��!j�#�t�'� _�mRen5
�+�[��e�^��mGUĳ��9��/@��Ss&��[̔_��S&)�)�"�S0|dkL��A	�A�l����	�$����O����Z��q%��N������x�\CK�JWȜvU�� [˧�C����1��с�������T&v���]�t6�ӆ���i��ٿ���~+t�3���)x&J����}�&��n���P��F�&�-��hn݃��p��-���Ke�H�f���{�N�μ��}�'���� �2�}���$6�����}�24(|H��j������.qg#���p�}b_ }����q*���^~v.���l�3����њ���A�)@ҳ����X����XL���T�ڱ��|v�	_f=0'�|:��-Z���o 2ݣu臇��+a"�+�*z�]����T�쓕 2��2�nD��v�7�:d'W'u�2�<�Yѳ5$�ȶ+x���ҝ�+��`'�*���E����]i�\C���4����m� w5(a�<xw� jʓ+��6j�)�6`�:N�4�{忈�;t�����`D�i>��f�J<��#�&���6�w�T�]Ȝ I��,����Ӏk��{�_�Q�"��s�L_kA�����k��,e���@��=�v	IL���E����J��-��P�Њx��I2�k��WX�qncJ��Ӊ�0_Ҵ��U��kbC���o��`����mBpc�����L�a���e�xa_���J_�/]�˕��o��H��Au��y���l��0�_�����qo��һ¼��Zc�-%�\p$a�����^��g���'A���] q;��૾����rE��r~�V����O�F��G�Ӊ����Rȇ������`|}��n6�⦧�}�D�T�B��X95`@���R.���)�u���j�䊍8;���yfƁ�N�,�nLÑȠ���-�m��\C?���/>����o�  b�
`�Nr�G�C�ݰu�O='�n��:��a2��-W�,��3_�Ӽ���Z���i$��b�׹�h�k��g�^	U6��Zn).�7U�_�}fp9�^,ػR���65z5<6�kT2���鮌�_��ū�a�$�3��&L�HF/X
�J��9f%�Sjq�{g̊Ćg��f�@�eDc$�2�[������pH%ll���?�y���~K/���X�1~
�ð���D+�����@��x����X��("�J��?P7v��ɚm��C�|�0s\��Y���6��6���J�ѭ�S�!C3�x줤y���Ui�G��R�w���t�6�j�)ң���9���#Յ��h�C�M�1�����x��x!z1&��=xB�k#��RA����ԻE��WQK@jm��Mw�*��u!WK���{s��e�o���p	��}�LΊA����:%u����})��^r"N]!��Lon�����Ԃ�ƅ�`4�@zs3&�3��Z��hz�ḑ�&<�"��������_)eBh�0c�>��	=|��]���}ܥ`^A�A���+�lJ>�c��.qnA�����i�	"�X�����E3�W/��ΜĠ��<��<�۩�B���(�-#"?����epQ��-�<"a
�]!X����O�v�$5����!}�jJ&U����\�����o�>'�LW6�����)�e�b�F��T��l�k;:yˋ.�G�l'|�K ��*�C��d�����N8�MI���A���i���iݥ.���(񞠖��Q�.x�� ����?�z?o~�8����O�p@u�F�hB�ǯ��Q��/ �?��Q�մ>�^rL���?� �=�``9w�>�"*���� �A�-Gj��d�,��1#�=�[����%�z��&��xH�����E���E�����D
����au
1̪O���2�XBHF��5y��x��ߊ��D��b��t��1�ā zXB V��<{cn?����A����R�@WHf��6���������TM�jq>}\��`�B���+b���0��pp�<��H��3=���4�۝2�>���wf�$֘oբ����'�8�+v��oͬ��%�Ge���;|�;Qt�@*�?�]�5r�i�~&�9�|8Ů[F�p�����|�ld`њ$r6_��#Y����������bRN��e������]D�a۩Y%�V��Ғ��;]RFsv�1�k=��b�u"��;A�	��s���Ѷ���I�I=9�W���� �R#��ܾL��;c�G�C��8L6���}e���r�&��=<�֤%��2УêL/艣]��jx���Ĳ��.�	x��cn~ա��Kp3�R3��)n�$s�ؿ��y���bq�ؗ�I�ԯ}�"ʉ1����a�I�1�o�U�궑{W��M=��C�O	a`�Ѱ๎��-«E ��&���YRai���8yU��}f���9�P�?��n������~VC�s#깟C��4���Yo�S#�][pp΋t��J~Z.�f)�Hp���X��h����/��y�<�X����	L�J���>����Kt<[ÇG�zh�IR��\�X��X;O��4�ߒ��4@��	g��q�u-q�2�XƧ��?��	�9LG`
���J�R�mB�3�]��duz;
 ���1p�o����֛���uI�'�Ɗ,�Jہ��x��~�f���"����v��/�>n=�VK�BEq�D(�#�d:���L!���*	 ������@��'�\�.��,zc��0�br��	l�t
�>��Wh>�.,���'�k�K|�b(U:�4|c�4A�4���Í��F��=��rB�R19��=�"˾n���K_����'b��b��`!m�ӕ��{nN?kE�]8a��Ny�@g������VG���t��W@F�#35t@ͯN>�Tnw<%��D�x��56n>D�o��>#�i%rc��E�V�-�e����
����O!P��m�/���}�rT�(ւ�k�pk�4�����z0ˣ漓D4r{n�_�����yM���n0� �� ��e���؂�i�!�E�2rb+`~:�0�]����0L���<����J�	D�S!ZOi���_rg�bF:�~��0ۓG4�6�ؿ�(���EXR�su��(;�#��yL�e�~�¼w �+G���lر�5_1�5���wDI�a�U����ݸJ7�3�Z��R���FA�q�l���|V���ad�wX6�W��'���q^�k/��-���s�G�W �
��/a��秎�S����H�K
�6+��+��CSԞϸ{��E�7��3��_��� �'�q���eK�ߡ��֐�^��#L!i�����qq�t��q��Ðf�1��غ�J��m2" �C���׵l!�)��B�� ���{�m�k�
\��~(��p�j_�q�M��tu}���vzH|]
<��� h�m�1u��P�ȝc8���-�5��-\�Ύ.�`
�7�`�t��+�g��}07Tw���ăvL^�������0��	��H^G��>P��M\rǹ^����6\���ǀ���G���2�H{����/$��t҇��}V?�n��
��ϧ�ʸ����fD ��_Ee`���OZ.l��S�X2r�m.��3���>L��C.��Q�`L-.��E�B����1��j%Q.|���Q�j��H/~��d��R-*��'���@���U��
�΋�X��0�!iA{��JN���f�fM��f�#�|�l������~�� k҅>śC���\�/B�w�r��.����d����� +!���?d���R�*��b��9<I�dp�0�ɻ�F\��K�i�f� "��Q��q��WF�7�T�c�׳M9�� &SN�������`�m�+GK�,r���r�ն�9�_�xN�Gх�