��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|�L��58b�Y��uޒd��G�!�N�;&� �#)�q����C�k���$e�+�Uy~�D�ݛ�7��oP��Bԛ���Ȱy���ҢƁ#WI��3��2� �<��հ#硞�LqyhG�U��1�DN������[��'�?#�Ct愠�L�t�T՟"p4B�T�}�DD�����։@@����8���D��y��)c�:�4��k���^M�n�Brs�:���5�]���e}nG��O�T	��l8<u��;D�����I��=ȩ� �M�`�6`���%!���U"Nb�Bp��I�5d/e��YLp�v��z�d1bq�9�quz�d ��H-�!�b���Q�#�/pPgF���|#;��R$�AnXHA��0���G�IvJ
�Q�;�%mv��D@�Xe^�t���x�]g��Gw��O>auk���ο��V�kE�A�`tJ���~��r"�ֵ"�1���XS��\�c�;�b/�N���7���d$�觺��U��a�?�w�Q3���.à@RLW�o����B��ʓ˛p,@J�n�uɟ���dல�y?�5�
T�A&�\o;P���w0��Uґf��^X6B+1J��D/f-P�5��s�L� 7��S�}�Zp�V0�>�ȑ7�d
X���v}Pe�~�ð��,�v>�7�K�Lm�B��a4A����}|�a��x1�k�|�KS�����Z>�ְt'���X}�C��hp�{ܖ�D.�G_�iI���(.J��"�)�vd��hcj�J�^X�3Rt�GS0�l
���k�Y9��Q��|#l����}��|���reդ�	k���ӹ���,CP� �4-y�,���y��%�Js���D��.Ru��;I����w�a�Zw��W��u҄iv@��� 4��U/w�n}��҆!"��.��NH���M7�t7�,y~�e�Q�1i��2��r�RA�Lh1>= ��XD����$��n�JJ�,���'_Sf�sm���yIaÝ���vZwy����]�U0����dҮ���yT�G7�/Y���B`������)�~kd�'�N��>i{�n[�
���@�)�"{"Z��n݋9��M�ew@F�cC�4 ��y%P9B�kA_��]=�]����=�:6	�-�뒕*���'�Ql0kdh9w`d���>ݝ���y
��R�4SHa>��#NI+���t&Q����S�/"�u:e� ��Ef����<a�v�´�)�!��}=���r�1����M���zař�ܿ��U�HOW8t�)���C2�����$�2��l�(��%�~���Sę��qMϓ%4�L���-��%���?[�!�J8�u�b*�!L��D?Eg�[�n��͠Zi]x�~!���V��C1R�Q����W�����ń\�~��EQ�������0��F��<���('6�+u|.�[.��u�t��ۣ�~�(�|8�²?U3���,���b���aI���Q�'��%.k#��a�����b�G<1�s���z���S����q5˻�>�LK�����u!6�q���!�7��{}���}[[�|.�=���/����Me#�o��,OG��R�d�韀�A����o5;*2���>��ie}?�׈X��Z���SS/��a�5ݒuB��������Y��6~e$+�*�ZJ���::���* Ƕ���>?߽Ÿ	+��%���n�R�B��S��~��Z	���??�a���u��"ڄ��t�1Ru����������?�ny��Z�0'��Q��So���t�}H~�:�	i-L���w�Lĸ���M/��"G��
jͮB��c���Ce^ |چ��<�w�����K��_�%Jzъ�4��^;��8�H�c�$pd��V��CD���OY�0�8��$����l��w��Ԓ> �uιƮ&]#�7���ԣ�ڻĮ�|��b�D:��
eh'��Q��к�k�P�iU�H'ɿ�q�Vt����)[N����aCZ���a^;C�G��틠̰0���.���F@����6�t�.�@�=��8��Lc4�2*�J�����U��wc�"����9GFRf\�`�����!Bu��˩���:70~֡&FY��ҝc;h�C����ᴆInz����wO��k7�E�dg-�ê"�A�t���ڕ�;�|<t�_��6�[� 'w�j�x�@٬���a�헫�����5W�D_�ˢ���]uMG�(Jn�s]�x0��Np5 s��+{/��h���FOz��A��_x��T�"O��ɗ#9#�m�'��`�SfX����Q^���4p�9P�\(R�)�xX�" ���r�� �uCt_��'1�j���MŮ!���V���
���b���Zzk4��z:� ��I� u�黗4n�M��+��}Z&���&�3�re(g�^'�	���6��.?_e��݈�{��B�(�1|y&���{?0��1�RI�4��) ��̍�۶j����,]��v��Ѫ�ĤKU����� ���G^<
^)\�_�Z�z��B�n���^�{�04�aP��������Q݉�>@J�D��5/��k#�%�*ګ1���0��d��`����E
��ap.�i��`.\�ab�	���l/�_F���uz^�]�S���+>M����9?\���1�����|����AHG�c�Mj����V�Q�S�rX�EՐ�vџ�G��Դ�|�ED��+;?V��>v���c{���H%�+�=__QKp��"�`xj��z��?O�x�9a�B�T%����Z��p1�Q~��op�Voں���d�����@+Ul2�A���L��~�jтj��95T�tH�X����h���#��g�݅��Rl�DW`�\JQ�B���R��2K������s�]��}hZ�[�����:q=V]�]����?dp��(�:���9��P'l�^��s��HH�_L7����bU
s�Y&�v�>0�݂"��ߣ���4��_�/���5�
GM)�{�E��A٨X]�����I����Ay�U�07b��KXi%�崢����\�v�ɹ��"��`\0k9�?�I�T3O������4���e��nH��z==��;3�X~D�L��O~~��4a��Q�����5��)CaD�������蝺QH�{��0y�>?�ǣϟY@�,�ۙ�Ng��9^��T��>o�(7��ȯ��+����"֪�x�W]{ʁ\��c�:��E����Q�9��-@)8�����@�bZsTw�oy�����Zp�Q�6��C�}����$6��\}���(AtM"ɇM�e'��/t���0� 9�>oT&!6:8�G�`���5���ohY�Ș́IXizk��2�%VK����}�$�[�	�B�C��