��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� ��)sZtYzѦ�#����������^{���f����@,�B���ul@k�"T�z-��0��{�oQU�<cM i��CV��Ǣ���j*��>3���B��1����ݿGi�b�2g��8��H�2m��@�}
�G%�p���.�x�T$X�v
��;�b$C����f$����D�j����+���DM�#��k/��|�S��p�k�ҘMw�����t���3��	�ΆLww���LG�\��*B/qR�n�d�"O��
���<�[�ٮ<��?^�+�#�����\`2Y�Ϗ�cR�W�G���	@oU�z%�� �˗�#�fŪx��>��1=��&��mErc��ϿY>g#d����WQ��Q��h�.�8� {J��=}�17=E-�挴ە&0�3HFq���F�W]E:ń�{�B:�(��=Y��َ�o5qxE�~�4 %te���s�6cܮu_�b+�K�s�_H��м����-�]�Ô9s���f�Y�5@�(�:Fl���t�����"���s,*�D|�ޝ�'/J���v5�������n���4��>� W����� ��驣�֢�7]�DÚ�\�y-DӢr�X��5����}'�E3c�j��6�۫�����0D>��Tf�G3�>�~�0e� ��d'ɔl�GP�j0d�S�T@|�;�'���t�C����K�j������E��n1�$b9��z��!��o��1V��%��xh�Xy�����B"�u����hk-)���7�b�ψ�V�*�㿓M�}0K���.��"����6�4�yjᔌ �a�o��������6�1s���S��.��j9��;�;��|K��Z�n�>bl�+�8
��+S���������TI��:b���i<<�� Z	?+Ƿ!.7��o��$.'����Z��`T��<�����,�9�����UV�"�մ�U�
��z��f��K�Pi>K�z|c'Ne�4�p𺜀���r���%O����d
��d��ӧ�h�A��������M���F���}��Æ�`�����슅|�o�ɖG���� ƔY�JvS�Q�Z���پwE�7�0F��}��<aI�F%�oxq�}�o�X������o�����V�|���T��b{�#�4�~(����@�8VK��!�>�I8/SƇ:'�(}�v�ɨ���%|zߘj��-Z��S�A׽y.��6�?wu�l��O�;�O�_�!`�<�E�Dn��nfߧ���@�cM8�@	ä�-��NG�p��(=�ȕ�:�X� ��n�������}wM�A���\�勉���~�'�B�>-z�Υ�(p�%m�u����+�[��N����j���>t�ʪ�a`��OC<mg��K�+}	n`ĳ��EK1P��ѵ�G.^����,ɭ���݇�]ˇ�N5km�/?����2�l\��D��[�h��I�����j�O_�_3�,�Te��,Y0�P�Ұx��P�/g��Be��F�ӽkmh
|����:�v���H>G�q� P�ߛ�L���R�ug�;j&��;�`��ug�+V�
ͺ�n7PH1����tm�p��B9�0d���:X��c!� ]������+���mS�hIU��t�=�����U�\zD�5׮�����[DV���=���`�-�n�7pk �t	W�G��	 G~^M^�O�{TW�V�3���z���Uȑ �t�q�&y���̄��	eX@
��t���=
��^}"��vy�#��'L�cP�Lf���N���7�"3�5��� 3���Bq�U~(�G��A��(�������<��큰�篪Ow'W+�{�n�^ܺf�Zδ{��=A�w803����@��'�����~�W7�(���#>�I��Ʌ��x�9W�:-=vn=C�p�|�"8sj��&M���т��͍@��� ������=I��X!ȯgC������M�����=3?D|\4/p�����2���m�,GE�&x��O�FT�NSMrl`�;���M�E)-Ng��o�C_��O�7��3u8��0�/i��:KcIvs��v\�����E|�2��q�yK�0��9T�E�)�)Y�����zB��P���SL0�7��4'��I��J���T�+�ӗ,�F�Amv؋j�*�w-^6ޞ��`]LN��u7�3I �'���B�)@�Т�D�1v���F�+�r��@��0oY�=�\hc�m@j
R�r�~٥j�դ�c��{^�Yd
�@%͂�W�FjZ���b�89�ME�xq���	>���9�E=���Hv�z�2�Z,��#����}x��<:��&Ŭ��O��t������[i;hr�d���v�q�e��礊:�v1�1�"��R)3nkü
6���, 
ML2Uh<��M�e�<wO�뤰���2Ig�[z�^\ҧ^]�t���z�Z(�U��:ņ��p�W���=����[�Q�����Vz���]� ��yi\D��ZB6���r��U��3�"0���zf�(vɣ8"!�!�N�R�@�d?��k�8�^0������G2�yf�NC�*�f04g�Jۈ&(_�	�a�����5�R�L�Wϻ�yo";�� ���*�|="�^�g�<A�_�d("W���i*z�����A����/�'g�|^��L�䑽��-	Y�D�Į����:�7�r?ib!m�!g���l���[��+�0{&ؤ��(�:���~��|%$B�r��o���3O�sM� �#��D�����ݡ�*���4���i����+\X��-,�U�~�h'p�u�p<ܳ&���숇��ݐ&�?�O CfAq%Xw�U+��5R���?��h�ύyyM�T#��Ԙ���C�=K9���-�Hd7�SP�	�L%�3�x��C�����O����T����ʌ�	ﵼ9�N_o��P� Pi�� �T�=�s.�	0�8ݟ�l��\#�v��%�9Z��:�fm�p��*�����Zx�'[��]��hԠD��#hW6]�^�0Z�bgZ�z^�҈�"�+cr��-;�Әh�Z|�v&L����Ӆ�z�R�$1@Ҟ��>j�["�sUG�/4�zm�M��zk���Vl�OD <�����������$��uj憒�m�D�EB�bO�ثu��	8u��ϳN��~�-
���f�HM\�����98��m��	��9�;Js���w@�	d��o�ht�K]�a=T��\H�=�	�Z2oN�<�%FT,��"$7��ߨ_xA�6�ц�G�@�X���a�y���X��)��x"cX�QT���TO@*wm���o��]z�Ri�7>s�r�b�g� x���� H�� "X�$�b�XmN�:�h����������������%����?ݑ������lyO��?��*T�Ah� ���@��J�-��.���~1����7�>�I�;cC6H�M�U7v>M(Ux,pZ{���"���/��s�nFst��`zv_(P����r�[�����}u<�6O����"�<Ǥ������������w��M,�5 !ee4���j8�Ft�z��(�BQ��4E|b��'=D?�������N�|�|�й(�a�><�(�z�F#$Ok�v�!�>=��	e��B�qg���a�cm��ou�$���k4���6-�Dh�!l��/G&JsN���������Tɳ���