��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,G��U�	�oJZ�@�z�����>*Q�p��~!}8~��m��sDmN��3\��\�A,��y��,�y'Zs9|�v�G��Z��J;����`��"��t�������UnRt��8WP�Z#+ϙ���\���~��/M���jы�IFA�O��L��oш�eՉJ�	1�h����s�7I��e�x�F(�1?�~�e�)�	��� O�%g��\��G@ tG]��L3k���w�_!�W����僊�> �w���$�%h��gZv+�o`�0d oq�O��+ަ0;D/���PL�?���o�T����n>f/��2k��ђ7|#7��V��⢻�U��hb�y��NU�cͩw�3��@,��#Ѷ֜"���t[�imA\wS��
 �4��vCեĔ�з"�r��%����s�'�������\�ߜ)�p{�&�$��:,㸱�և�R+}ߐ�<�7��c�݃��&�{\�J/��^�U�s�Kj9���î=��I?䁋�	A�-�M��ޢ�sP5��Gd!��?t|�(Vĕ,�|���y�����6J/�?�q35cR�0��M�,�/k�r"���s�|��{�L�������4kPLM,m��y_nzS���9G4\�~m�����%��?�P`�J��"|��E����|�3�(D"��4�ѕ@ֿ�ɹ��@�7W1�c�/PX4�4��|u��."�߃Ve�R�&��ujFD��㰊һ�.6�]�=r.=����J�qл`�54���܇�=f)pA�/�n2}�{Kc6h!L�C>�������Le��4\LK�5���gꊷO4�:ZGz&���޶3�~�$�;��)�N7�����:���$�L~�]���;�i�X�G+P�a��Y"����Za��a���6�t4�K��(��l�<��(X�5;ٲΈ���ʣL�l�2��t;N)0���+q�45&�Ad����=:�t��K�����:o���()�L3���L���nu�f&�����������o��� qI�V�tb[�}�g��adp��mT��R*̻W���{f+N��juG �L�$wPidĽ�|�5<G�>�꾭%	"$�䎁�|����;h*�mlɶݯyW���]��X�RT���H��h��}e�a�4�#+��l�����R(��b� �Zq�d����� ���������)���s��<�2����r2��98������SQ4ߠ���W�bvX(������6���̥������B�o����`L�OJ��2l�����h5|
���%�G���(06�� ]a�s#��O1i����лgT�h���m{�+Z8f?�躀g׏`W���Z�XΕ�I/W�B�6·��}�����m��d�x��c�B5m���Ӂ���8����$��wA��o@��9�3���d�4<.#��C�Ժ+��[W��1
���Z����CƆ���rBJ�α@jDKzj���Q�A�����K^����������7~���_�P�a�}����!Ǣ�]�����ZX��n^����-6d��!e)o���"t6�J14�=���`�����|6��
�w:πed���#���f c�H���M����Z�������9tP9�`�P�m/��Ӷ����U)�p�4\Î�N�u�;���+P^�����V.8���5���r��Yw�D��	>��I0�����#66by�_��&'��C��-��p/e�$
�잕A�cZ&�U���-�?_�_u낈�7]$`+���ks�C�U�ҡ�{F�����/_l��l
��>_�%��%i�!�%ذ�ܒor�8vM@10`�
�����Y |É��B��Yq�� �Va�O��P�V����x�@T�kf �Xz�]�m.�C��g��s�u�S��-�fQ@��D�E+�6��k��4�6~7���b|^,6gT|�M)�;\c��ǟ]��Qs���J��16�K�w���&4F
aTm�j%�t�,ȷ �c{�rt�0"F�*��?�y׷� �k"r��{��̘��3�R;8�w�O����=����l�=I'{3���{��q
ä �Dt�F���=A/ģ#&Z*FM�:)!��f[:���^nY3��f�g	��Aż7;�-���(�ޞ�'{�]�6�躶I��U�=��Wɥ�w슟����Ҩ�	��k�c��^�������´��4TױF0&�o;=�:�$GY�K/S@��Z�u��c�
Q3����� ˏ��T*�~l�<�x��N�`6�M���܆x��Xv���+$F���_�e[+ۂz�#@�cn=����T�����@��(vK�6��)�����$N��$ĕ�(��z�{�#x��U�sb�E����C���w/�
�n�o���7���	�p,-L��.4o��� ���]:�_A%������ �œ;̎Z�]sʿ���T:���)���%D#�
>���#�AN~x�49�"�λt��\j() �JR�M��Gz��=�B��I�5��w*�ԙz�&G�8eR$�t#O~8V*��t]㦹s��dr�A�N��Do㞛jeO�re��x�I��K����YQ���U�=W4��6_���(�����!����v����N�5��މ���pY��lH{��XU,">��e�w@ݮ�/�8~6 1� "G;}�N`��r��А��n�:fsr/���Q�A��=�r��kG �m�v�zF�\��g,�g�c����h9�v�[e�"���ʂ"J�j42�m�yLpS��4�󳓲�O���O�c'�Ef��:��VNE�<W�8/W_������.J�B�:�ȱ.�T�QS<�b�}[�g�h�;��@'��ީ���M�8=]����������Fk�E��Đ'b�.i ��t�Yyy�9`����'�a$�b��g��z�`��rq�nm݌� ��ܖ��.阻m���xw�/�*U��T^d�C���Gl�t2z� 5?e�@WW� *.�Ն�+��$!�ed��F]�+�Y6x��{y����*=�f��SՍ�����{3䅣���c�Z*�)]$���X#��ύd_��*/����+\XԞL_M�?�_h&�L�Ui�5�=�m���S>��s���>-�q������$���>�rw���G�'�m2.��D"�]8�5OQ���q֝@��#9T2��v�䛾gL5�ҍ씏K���i9�zV��Ms�vv�6cb�K;$� �8>~�D\P���j�s��J[X�$;���;�O��P���z��*����}[� �@R�L%lwʟ@I�d�RK0�ݕp���r4��$���f�>��2Nι��5���$��)�*8ӸT�,!3�M�Ͽ����H�/����G�o�((��ֆ8�#��XMg�m$�nq��@����_)I83'd$��s?<�y�U %}/+�if`��b�jɣ�&����/������Ť�b8��f:e��������1x_��o��dI��׽��78�u=��u���m����F�3IR��,}�Td�t�ub4`��d���b/� m
&n=m�d�t��KҰ�#Tm� ��כ��1�C/���٦b��u���6���/�r�����շ_����w	śJ������^���q$������yÅ�.h\gP��9������a�L�F�M@�	K+��Awϩ�����;�P�r����"q&��v�A�>�:��zڊ������N6!y��zo����ֹ�t�4dP�x��:�Ƽ�YZ���:�
���Dw�g�,mz��S�޵ۡ��m��v����]f�7| ��şk�*�#���U(k���0Ǒ�Cy	�D�E4F�&�;S�W�9B�<9�?��vtx���n���K{Ms�+`�3�����^�we���Na���+���^�5)]��'0R1d���L4c�:q�-b�`[�>*����P?Z�U���������Ғ�\��^�n��.<�V��V?K�u�#qȆ\�H�$�K��Q`ݬ��Y�3A7]���ε	&}f��OܫuPb�ϩ�.1���e��c�G_|���P@R��|��D�g��/fe=��al�W�S�B�k��y�ٯk�l���k�#W8��ѣ�vk��K��A�S��J<�l3ywG�56���p�T��b���/����� EAp��{2}e�t։�(U@F'�p?=���ū�{��������A�x�_����"%�{���c�u���`���p)��*�!��ľ�ܚЖ�(���d=8P��59���9ٹ�sV7<��+7\����v�z���;z5�Pbh�1�YM�ʘI���xnϮ��H��lJ�mp�9C���e����.I��ڋ�ik��l����ã@4���wDH�����m�-�#��1>r/T��@�I|p7�<V��>���aAu���R��b�JV��~��졀�A(;������R`��)GD6	�=��&L{�����^^/D'ɏ����q�����pE���7#� &k��bɌ�`��0�oH�q�d4�3���'*�>�_�D��\A�r��[�e���R���P2γ��B�NQ/�>b�dA��'��N}M��W�:�5�h�(��T�!~�O+p��n�D�$�a�d�&�7L�;��k�w�R��C:k���r��7�̟��F��^�q�
=�,���N�&�M�|7Ō덞��S5% J*R/��]@h5�HK���C`���/v^���l@\a���9T�X���D�G����+����ba�7���Z1"
Ӥ�vf����I]{�6��N��J��%���yd|f�ߒM���?%*~���PS�ǲXe~�|)L�ͻ���ީ�)/��CX�� z91}Z�����DǕ��wy��!�6��fd�6|&��te_�g�v
��|/&h6,�E2ܼ����uvk�K���E�m���2/ݭP����$�pBS��v� A��$�S��tTã1,����Ys��t$֬��7&F+0Y�:�q��5�[AT}�"iɈ�TH���׼X�T�D����tW��o�^�����hU9��W0��8�ؒ�=�,��,qp٬��CԬ݆%>H&� uIzOd��s���u��)W�LOl��7="�bW����t��u�WV�.T���w��UZ;���<�滄j��x�Zz����~z�4���n�Xic �&u0*,ǭB(}�X��vYߩ��Ι���f1Ԓ)�d�ܹ���}tS�KIgP祮�{�R4��U�Q/{��w��^y,��
K�'񴠗+pQ`��y��RN	���a���#6r9�gl��H��ڿ��_��������F�pL��rh):�@�������|�ș�#+���	`���������{�"���>���%�
*�#~-i��
8�܂@��3�Es��*P��ؾ�'z���P��Y�0�&���O�F�k�QJ\be�[ ��:'{/.�cĉW�z��]� �i�~�HSi��w�B�(�!�sy��E�pw�i��ē��j���T �� ���qfu��*�ss��Ue�E���5 ���-4��<�Rxc�I}�f�m��h"c�m�z�Z���]�	�w�*���j�9���Aǻ־�`����0�:�P���^ӣ{�t��qu?Ei%�sm��u��Ϻ��$�jxH�Ö�Q�=]�S.al'%ȅ�ݢM�������̠O��
@X�"l�X�������G�܊��K!w�a�H"6U ��'���y*�H���������(G�㔹�4-"�-7�>�xS;��ľ�
�hk!S�=�Mqp���{IJ���V���! }�p�!C%;��Ȼ���_A,�K��K�v��g5�����I��$��F=�ƿ��1
Ҷ�܎z�\�[�2��u;�;9���K��ז1�FC=��b��ҫ}�*���讶��Jd��=�7�[�;�`/՜e�:R�Laȏb��u��
�l{%۪-d��wCR78}�Ti� (�r��@j	�D��K>8��h+D��i��6��#����G8 �����y�C��r֪�N��s���B�ONŨɛ]��8��Lhڮ�2�$.��>�o�>�%A���ٳ�KQ�tK�����Zn	 ����Pn�6��АE�W ���ƊgkEB���2{�&�(��4ڢD5`iID���?j��PK^̪�Ǯ��S