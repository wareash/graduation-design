��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�k�۸�m�i(b[�{�㇌�]�i�5'�`;Etg
<������H�W޵α���N-�`��6����ݾ�FF��eF4��_}<�ےA�[,�|{�?r+-��]n?���A'xin�XO�v⨺��sZA�R4��g�psXdm"�d��Q� N���ُ�(���o�&M枯���aO�1f��m�6:�aX�zj��h+��� O����CG�Zo&�g#�$�fa�')J"Y�p�kÅbA'�(�aMa}��;|��c(��y�O��U�� �<��`�� p&z��煛.�"�BI`�1\����LW�����N_�y��F��������v!K��i[��)?��,�Ƈ���0p�b!l�����,kWF?��4!H1�,cSP���j�ɚ�'��\�r�K���{9kmȡ���D���(Ê 4��G��5ΰ���l$5°�[�k�pA0F�ǨI�r��J�z�fGEbb���`�����!c_��?j���f�W(iJ'Ō�O�H{V&�,n��P�=��~�m5�т��{[�S���l�uj2f��>c����:(�]�u�[���K¡=�0��;���Kc\�#�2N,�V�y��`m���u?��#7%����.5Rq�4��e0�2�����i�����☬D�5�cP�O���O��FM�5z�U&�n�T�Ba��-g���_6���ƚ���ߚ��k�e�0�;��;n�I��8��
ੜ�h��Z���pq�A����U�����;��Ջ�D_��=]�~P]Рb���
~�����V�F�2E�F\޽�;�S$e~��?�wܢ[tx����&�ے�a[�Jt�ZP#!'�_��E�lS&�C��V�@oڠ^ �َP+�xH��&��K'N��>�!pe⸇=�% ��w�1{� h7`-��l���k���8�:��E�E����LE��Sã�&&n8���I7�%�k���ղ�<�4�Q�A�1��X:P���(����X�u=��M���o��d�"r�J���P����`ġ1)!��0���>�ݠO�۽�b���`�G�.�y"�6��f�Kp�F�f5��L� {M4)%��T�Ӳ��H�l2^)_��Hmؤ.1-�6�>��c�WȈ`�0���39bȹv�ZE�2�8;�)�d��Z���:{"���6\�q{��#҉�!i����H��u�Ai+�9w��O�@��u���]-�����{���>X���kG���ʳ��|��t�[�6��׻�r��4d?Ƥ��h-1�^�����4� �F�%��	ݐ��$�a���{{�=ϳ]Ӂ@�w�r��&>*2�Ɲ�fC�g��DB"A�>��ڕ� շ�#�L2F��q�d�����b�����f��QLO#d��<������6Ľh΀�Ѧ��C����H��b۹Oh��IXNr�[R��=���������ĐcLij��e��
ɿ'�ӧ�``CX��
+�K�j��F4�c,���*8�o0��)}LxE�D�E{?��U�mBF{�"���@a�ˋJ���zW�@}��T���;v�X�� �x!�DCx,y��6	���|pv����`�{:G�t�+񚮁�p�U��%�����ϕ��7)�5r��� -��Ayv=�*"����%��c�z��S02�#�hX�3�d��