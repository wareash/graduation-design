��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jåا{�\�u�?߷�dn@6�zf��r������;�&��0"�*hT~�72�nS�B�0n!�n�굑�5���ta�� ���:��=�_sy��6Q��\�)Σ��r�����+>�Ȣ�%z���nIӊ��	��W���q��=��n�j�_�1*n8����T%Qa�k���g��[�rX��3�[^��&2͝�$�}K�*�%j�P�H��B��XY��%�*p��rSx{8
�h�'0�>� l"�{���!�̀�j�9<�� �����߶w�@^w��6��I��q���e<<>�g�j����T�g!�5K�u8ŀ�b�SB��$IiX�!.��SNFH�a2�5��M,MP�1�*��x�+kq�e�ȝ��=�q�{�6����^*?2�*Sl�L��ע�Rf�M�!�_�=��X���Io�R7����9�a#s�0�^��@�[�w���V�b�2��T�a����QU7\<�N�(��7�%�?v4ݶQ"o�;�9.�n�"��l���ǜ]���B�����ڽ��+2v��N��ց��7�T�|�1���3qd'e��#e^%��F5Y�g��Y|�F$�ʯ7����ݙ.\'�S�(�c�!c���3R�y4�ڼ��E3�djXc��+�!�D��T�
"�;�]ղ]���.�i�=R!9�|Y�S�]�Bq��º�$ؐ�^�ev�a�;�	��X٬(m�[�M�l��H'�/��v�����0�Py<U�D�䒮0Q��U���(L�I[�
�ڄ=��s��!R�5&w�d��*w�"�&��J�VXBKbdH6.0V4����������1~�
uK9��i�<埚��m�}Qdy�W��^�m�+$"UkrI G�{<F��X�yݯ��'��&�0��$�ތ����Ԡ�J�p�4�+?��E��*�(�T���h�Ȓ�PK�q�ˈ�u�HSY��z b�(;��Ԗ�����'~e������h����;uX�_�Y���B�o�ּ�.�"����b��e�X�1����n]�f'e�Ono�L�E��Vm��5D��Mp�w��nj�Fx��yZ[�[���O]�B�!��Һ�8�����7^5�$B%#j_R^�_���	���$�Ԯ�D*����nded�GXP�����p\Ĺ�_^M��'8-f*ƛ%���V�Boj�A��c7��	���h=�EN�@�sN�����o�b2
�F�#v�Q2
�xŤcY��h�'�^җ��y�DN�Z`��ʨ��td�+h76D?��{�,Ȏ� ��fF'�J���sr�H|=L16'?1qA���ǝ�6��ص� (�
�̬z��<�M��m�w�����b>�`u��胨�f�p[��E�_�MkRP�䘂۞�>���K���<���C��P�|��XC�*ǐ>aj�<�X.�*�F��R�n�O���+`��y�ȡ,NĬ��ߛ��_�=6��J����Iqu��Mfq���ҩ�AW��4�M��_G@{�"xG�v^W���l*o�M��=���2���ׂ�<o��{aj)#w������O��ھx��R��g���-��U���2�����q ҋ���LҲ4	��B���s�E�+=W�2�`��;D$�0���,<#��+�"y�E�\	s�C�_J�H�?��$Ż$a��X�롆.�?w�L
I���phj�)�v�r��3)t�c��78T^Զ��pc��洣�v K�T7,�-�F
,/���f}?]�n�}טf��(����KX�	B`�6� �θ5>�2�I<y싖�%��:��/��^��q�P%#���^����J�<	��B�;RX&����J�"����sU��:�����X'����͊ff��6 m�6��.���,ܚ�?����X+R��h_�Q��������<O�Q>�ʛw(�I�S=O���r�o��fz /�7�NF��5�.N��j�;D�5�~�ܠ6k|q��|�~Q�����9�Ɂ�:�{�a8�l�=�J@gx�z7~�
󒑎���G���hx`c��pJ���4ם�-ρN�+E��6�O��"feƈ�Om���a>��7�V�	\/�3վv@�M�e�R���R�y۳������E��+|�����(�X8��5�I*��s���)R�{IA��t�n	r�ߎ���`{�[�p�B6����H��9fÛ��kX���P��SPe8.��:�q#�t�� ���=�;m=z"X�[3A=�D��ȷ�ϩ�o��f�g>hY(�u��&|+��ȓ|a� ���ϓ���Yg|D.�
�韑ag@rO�"
�$A���xT܈�kKD6W�21��QKC�RVg�Eo��VM��"!�����=qJ0�j���h����v���7-�
��OiN��d���_��3�t�����O�if_m?��!h\e�PR�`_կ��e�P
&�6I4��n�"*��3H�J0�� �.)|���\�� $d�T���^�|G%���}T˚Jf �n3��h	�!8��`*�w���L��&��o�ጟ���%��xM���79A���j�F!V�����L��@���֯z��c�_��تA
��Kk²HpT��%��# ��O8�4�ux���)��|BFc+��P� �󉶬��cޓ���~���|��n�|����B5{7�H=LL��5��꩑�~Ն(Жi[���e��P���y����{R���I�3������������4y?����T��˴��� �e�����?4\���V�"�)��#���`6%ཱ�?����~�ɳ�?�~���9`H~�2X���V�=�-p�^o�]bq��{N�b�t*N >����)�qĶ	����"�>p+X�X��b�'
���)�̅��>�&�
�԰G�!,,�?��1W��ϒ��p���5��%�=o��g��A�R��Y��R�VOK���j�b��z��c]��! �g��d0��+��ʍ7�\�0�+�\������E��:�
a��U���A�dr��q����5���9����fw��_L5�����TF�Y3u�@�n�L��w��%����M�ʽ��D}�p�Υ.y�ˉ��j`�U���%"��)�x�xtfY�6)��@8[ >a����Q�LQ�8T���ڇ*�u�>�����{�'��>4*�e���zL�c�ko�6h>��Tf�o��/��Ix;1�P�����C�Jmm@�f�-=}��(��Tq&�=g�cCt�d�x.�|�y���X�枱����E݀6z�f;���s�#c�8����	�ۭ�-Ap.��w|��y�_r��U�}�� �yiV�^E��Y��,�|>�}��X,�Q��ZT��9������Z�4����x��P�a{B�s��]L��B]�1sK��z= ����GGϞ1��G}Zj%e�s0�7Ì�qV�{)K��Z
	�DBB�}�.��ש�5�`UY>������Me��XTs�����,%�i}I5ʛF����߯s�P��<��BW̷��
7-	Mf8r�c���"C��d�s_�c�i\�5�O��Jl�H���,����Ѩ���{i'���+����c��N�wG�GEaC�Ut�ɜ�!�_���\Z�s���#�F�+\����u��e�/	$T�v�O;�[ĈBk{���0��=��3>���?';�T��"ӣ��l��Y�.����8���
�/��R&H?�a����k�{���IC�N���.�RN��&�嵖��D)|^E�"�l���-���Nq�޳g�h^�˨�M j�d2jn�!�ôo5�_>��8��[ֶ��w�rm�F��p͒u3��V�������'�Zf��E��#n#XlC�v���z�Ð�j\�>vN
�r}�ۭ^�f^k�������l�FL�_r9��-�h�9^�M@uL 덬�i��Q-b���i�Բ��*�P����J�9�eNJ>s����	����I��zS}�
 ��6Ԩn� ��3�x��.��Ga�ۗ:/��� w9��G@��O��Qg��R�T�%��?=��"�b��9��s��Z��m��lWjr�E��v�DTP
Gg������N�%��r������A��?���=�"#������y��"1�P�e���yI�cOq{щ�[�^�d���$7���<WC�a@�<�D���!d�r?\Օq�B�T�w�R���(+~�8^m���3����6ؚ���n��Q���%�S<�~!9�`�P-.����A��N� 6��&|2?j�!q� ��;�&"��x�4�To����Ǌ3���Yi�&M�=! �nI���;�p�8�]ی��L&=�r����N�q"���ɕ��Z�6�Xy��ŗt�?�e�ð'��v]ރ�+������q���x�i+8�������@'J�dًa�����/J��&B������q�ĥ���HD�٫���ɀ-�іNS��fn���]�Qrg�֕i�z��B �[���/֡�I:d7U"�ȍ%�q���mt��Rq��t/Mt�%!�2[d= ���^&c���22�=M1(-d۞KKt)���S�Ox��R(�r�^�������k�&��k�\�\O}����.2IL:�{����9����!��M"�Pܡ¾���(�/�+���*Q9{W��^j��Y�J��FO%�4XD���#fcw���Y[�x�zD��g��1iG-xw�|?�-m�3|]1t}��^�iE��T�4ɑ~]-H~7��5�0�6
���MGHa:��u���6���&6��^�됽]��\�(��>:w�4�T�i��4IhDg+�ed�="�0���>���I����A���ꔏà}��W���1���dVY��Ń�b�S��O�eM.�*m�����nlAL��'�b&LĜb�Af���9�O�F!��Ma1�������1q�����x=: ��*�{�)���l��A&<d��|9��A�E9���;u�o��:�� k�������7��Mn݃
[��n:J%�~�m-��=k�H����2�/��oiqˬ�6W�t!����Zm���"��E,�/��V��g9p���Δ��!�Y5�O�,8#h�꜓�uI�9��W������r5s�tԮ_��N�$��!u�V�u�!_躛q��"�]\�N�۱x����σmqs4ʮƗ��
Զ��㟂x�:n�t��֕#x�!�4F�����qB��blp�^�,Qİ���"|��ʹ�@eM�$�Ĝ���/M�- � �4t.D�Ibۄ�=lMȅ���5�آ˩�'sϷ�^3"�bE���t0�MW�,����A�3:fG��8=��z)^f�� nIQ�F���$��n!oc�)� o�Ӱ?mz���P/�_=���0{l��`:�v����K��xz��&��E���/U��lD��+|fύ8�r�(�1�%�w:m
��
j^T����:=�H"��fVlL����IK.�k�/�����ڥ&���/���-�|��=� ����S�^��ŏ2���ԧ}�Ei�u11�dߪe��)�����~�K^��LBx�ecl8}G���N�n���#U*����A��B��+o:fGʊi�H:�w��#wj�X�'H��lh��*~0|��9�JgZH�A��G�>��#D\�k�4ut���Ӻ�^�.�d�si_EwK�PL�~�F+��<FR4EJ���N�_4o����C�g��k�#C��0U�h(3�T7��<���Ý���4�)5�?�\&uAFO�:��s�#i���0�3��[�B��z����:���vc�)>��I���mgtSK�,DB���u�ɖ�+����q1U�3���z3�5�l\_~28�j&ߍ����:���Oܾ�ƣ �ȗ�lh�]�PɶJ��֧6ǍV �P����b�?ݐǴ<�wة;�0��tex��Ԗ4�I�)Y#�D�h��O�[�v�m:����q�;n�k]�,�N_����' �ïә1BD�&0�#��T���������A�( �:��M(#��m�������Km��A�5���V� ��^c��6Ib���{bz�����u`
P�����#+�����m������i��i(3rf��Ҵgxlp���ꗸ���=�+� �����fh�'AE�%��$�`\�s=��	`8&��0xG�$�	FEc�nl�s�0Lg�<��{�����G|��:Vc�QG(��7L��id��]=Q��dm�*�\1
W;S-��1Ǧ��a���'
�h�M��/�����Mަ�pq�Z��	��N��O�i5����O��y4��@�G�C�I��
2㓨,�'W]�2�B�8&���M���BhB��љ^U�B��22�߀ь%�&8��b�t���
�ՙ�D`'ǁ%Ҋ��c`/���]�w�2�,|� ���f�?�h-AA���|�o�o^2��;)�0���XniG<����!�C�U��q�bP֢;��xa�<ck�C*�哊�a%A-CL���|u����o�8{ ���~���~qK�ꨢ�w����^c�� n�Td�{�O�&ה� ���i�md�]Sf��5���$��������i���I������|C#��@ Vl>�E���HL�,]?�����
�<^4�2�㬆�g���vє=����{�/���Ϊ��'P�����!&���x�Mi}�V���g����1e�+p@��܂D�����'�����t$-e8w�����^�	��� �3�G�Tz�sES���L�J�y{:P5�����Wr��[4L�{s��@600���*}ۄ�B��(���d8�5�٨^E�ڛ��J�D�}��Յ�*������}�N~)dvV��$�t���\(��%w��u{�{�00g��O _���qoL܏>g��jTCs��
�;��p��mc�lh�s�͆-JwGR��F)S��g�.�CS<f�-y�Qx�k�P�)��	��w��Cқ��F�c3�����;�*�v� ��l��N����=�ܨ_�3���>!%�;f���}ɲ"<y��ϲ2�����֍d�Bݪ�&�O��qo���N��[97I�6��J*=��=���ʁ��W��~�J��9:�`5��އ}7}�ow%�~��B%<
�P��ZM��aǯ�"�	�j�#�M��4�ި���@�
��0��x���v�R��y���|�"	���Q�0�I��P���1k��G�����Q��m�����)�#P,�^�"�ɝ�h��=pю��:��$OuO*m��M�N�
,�p��%����_�$<f��v�B;�}2�2�
��*pa����e��������Zr�8>:�0��k�+�G�D�T���r7>��7���AV&�k�>�2W �2f�e�9��43�p�͂�q�	��udG��;�1������BnJ��B�w�ފd����-��̪A����jM@��U���@
f:2*���Je.*/��ׯϘ�L���A������1�R{T�ߗ���V��ţ�=+Hi�.T���ᴊ��R�1K�]R�����v�m�CT�gl͞���細(F���x|���/�(>sv���NYDӷ6�O����VD�G��A�H2����]�c���Ca�G;x�ۭì2��4o���a���Q���J�̌X��e:�g �䅫n8(`��	��p>��K�ʎoV7�����(���[C�0&b�$�z��C�Q�9̘f(�>���U�Y@�w&����<�%�#�wjO#l*P��rqU.�o��;�����bO=f���}~4�����]U`�p�r�mx�\vU�x��.������}�����d��>�_�#�U�f��LS��g�D^� �޾7UL�7���]3��f�������g�Kr!֠gUG��K���` P�Nwɏ�Cm��}e��K,}2X9��_lA�4U�&�9D�lA�&qj�X;>
5�6d�14cQ�ݤ� :��]���*j��ހ�қB��?��1d[U.�+��NN�N�M�v��>���)��-N��%5��0�ti>�uW�uv�x��imgP��#���j_��n��
@X��/i�Ooj�<y�y�f�%���vQ&z���L3����@�N�u�MZ����JW�9���9�X;.~@L���Q�֝��w��"E�Ga�n�'u��bǒ���JfUp�v��r�[��c��]�:
��}8�e��Omz�������-*��6ikɊB�a��y�? !q�GN�x��褐X�V�b�G�V%=�ޑ�s�����hA�tX�O����T���N,K>�`�{�c6\��P�P�~�ԁ�E�k¤��!��6ɬ|=XD���rh3�P�K ��K
4`y#T~��Jǝ��)V��ld�p��������SIś&h�m�|"w�wb��
g��n�T��b�g��(�2�1u�kK@��Ҷ\��y߹��+F�D��R#�-��8�jaE��/�v���+aTr����2����4��<T\�J�y)��q'm���0GL��2��d��W��L%���?���u��ʦ�F�HD�ꞟ*Ӫi?��=����_88��LUj�Iq�m��� }�	B��A��t���k�! �(�;}ʕc@X��c�R�d�F5HU���{��&�y��\f<����S� 1Ne3bQ�&[ic�A3#��+cs�]ӝZ��;�F���^��[Q���D;b��_E��}�I�@��͓��ī��8B��^���di���v'Υ3u�"�.'���8�N�ڧ���@y|_�N��p%ܾ�I*��<1���dQ$��
<9�ˋ�/W��� \U�c���ɠr�����fa��}pP޼d�e>�fU,�k����N%�»��{�y�6gj�ZYC���Q�N\�AX���&���.��H�.���M�Du�Dz�q�������p�2�h'謏�H���'���AWK/sy�WX� ev�X���y[�1w(��Z���bB�
	���:��X�g��[����7"��!̜�X�t��]^%R�V����Ā�xsf����9V�'O2��FՂ�g<�]��H�iZU��Z����		k/j���iG��ZE�<%��P��$X��eS4�7��.w�\�}X��e9�s.���*|i�{�˘�4�#��b���/���X�-���n3�Yc����R�"1�m/�;k�L�X��`\���]ȼ�8� ����8�޾��"�҆ATY
)�H��8��R�s���I��$��=�YhT��JA�t����}gFO���+�[м���0���_��%���V���s�����wӴ�n�f��'��*8�W�+u�b�{ǩ����d�_�^v�p�=���G[Kۗ���h�m�k)���f6	�f&e�8)�,��$ �?g��/��z����e9 �ped�hy{g�~]*
�;��-����P��.�)����;�����劋�M�H�2m:bEd>3MF��+Z(�V&(5�L>�&��:��qf��LZ�Y�K�]��rJ�j����A)� ��l۬"����ī��4��kh^�j�$R�����;�Td�z�U�ej)Ă�������g�@����z���u��i�"��ӭ<Ә�t��-,)3��W�R�J���Ҩ0Ϻ�x"����4�Z���~B�ۇ�h|w�V��}��`.�. �*�"�^�L�t�屮x
p���,�߫C��\,�6���L�2�4pl+����²�z�q��n������!�<&57S*n�����7�@u?����̸S�g���>�iR `���CV����Ȋ\[��k�j�ׇ���S[|���UQzC+�N��l�%A�@,҉u�͏�sl$�]����ʚ�
�z;���!.ġ#����.���J\��Zg�����(������ ��1����=�s�|�}��@{�o����������)�"�����@^��h.�	 ���W�|������Ϥʢ�8'kV�)�%9	�
�.�cs�;Ң��L��jFO��,�+v�2<,૳��j�ɱ/QN�6���$grn�3a��'\D���(s%@_95c��O�	N��&���p�v�h,��;sgE���I���-r/U9.���zc���2�c']?�����i�f �(@�b8���G-�]�K�&������ғ&��-�2��`���Ӭ��~����K;x_E0Ƶ�ɹ��h
pma��)�k�#cJ<O>鰯W�
^�H�MN׶���,���s�Ύ5�䬸=�Ui�E�QJ�Ǩ�Z�#�y��&�z�mQ�ŧ��̥f��?ـ�Qہܸ� �?�}%Q�9���\���p���r�H��n��>B�h�L:��蟴e�Y�IȽ|�<�NMo��(a`�z�1u�im�C)l�Kqf��Ĳ�ڶ�-��^}�M�w8#��I���*ګ=����"�����g�qj��4Yخ����jF �ԙI w������l�.��+��"�
�ө��R�lqa2�)���U��R��u���>��Kqi�V�#M��4?�D�f����$F��ӭW;�jA�0�~������C�y�g����&Z�X��IQ����G/A$4Mg���i�Ν�2�C�o�7}7��4�����]�]�k6�?_t�K��ro@~P���W�9|+���O�	���5���o������XbΨ�^��2�dO�#��;9,���
���N��� ��BB!EM��Ju�ݧ�D��Oȋ��t�/��qB@��8��Љ��9#Pr�=rE�R�S�$*���O#IҶo�uF����L��_$��88����=��p9���&���6ݕ$!wwB(@�y)[�3|eb	��9wЎ�G}�?�س
ME�JN�B���,���:8�]�g����d�Q"H)ŏ�`�����s�8��+������m�|���e�5�T�f���ܦnS��R7f֌Z���3�,_�u#F��;�i�0���O:<3g���#&��n��d�G��"�ݎsT?��t��!��! �q/(��V.,��$�Ћ�G�y)�N�)T�J�8p�BO̻�.�3ְ1�b