��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1h,�mwG�� ��q�
dh������n�5ӫ�2
�e?4�K�����ps�/)k޼��������a?SrL-j7%�"�1�z忄Q���͗��2��B; �/^R[����wd��\���
A3W���w2�;�uhs�SE�%�i�6H� �P�6��v挻g��Z2
�*UO?���d0�0B5(5��������\��B8�I�~ˀax�b�R`�)��lȆ,nUoR����p2����vm�˦\+Dq9������;�����fg��nUVO0��+=�����o`�3�ŏ���/�rGm8�W=Y)Jٻ�W:�29�5r�i��~���tH� *>�m`��m�$���A�Q�d6\{���-��o�b�5	�D��~���"�De�T�.%���_v�bnƢ��^i�z�Bs9����%t��S٫3x^4�?92��Յ��A���#Ik*H�V�������V�R��x�;7�-�(2�L)V���E���.�K��>�ο/e~��	�K ��71�y�!���~�7?t5�R�Oe&>��'��=gX��"�~Z��߁�<�P��U:aY�*��r+=�U��󾘉�Ju� ͏S��8�� ����Al�+��`�*?�:BI!gE�80��!� � �wdG�����2|3��&����=p��[ݽ��d*�g����B	��s��4|Uvm��D�ce&OQ9?�ꇈ�ЭX�@oon0�y��@�&}�aj�SOL�Od��. )�;��W"���F�4����XR�$� Ab\��A���hc{]���3��J��*=����V�.p�ӹ|o��w#&��������8��U�D�I|�h<��+t���_5�B����ٕ�OJ�]�:��	�D(c\� X�y�Y�ѡ��{�o�@y1�tB��Z�ʞ݅��"�!���sU)�8$��cO�a���D�]�`�p���ݲ�}îQC�ִ�z3�PaA���iC
�lv=X�� ;��.IL�ǵ�Ƹ���+S:C%�s���J@��^Z�dئ:��C�0�WsIP��ѥ��7����y+4����)�m����Cg���?ϞK]C��r�s�t��e�$����wG�^�xq��-؛��H��!�>=�`yaG����\��С�+�]A�����JY�R$�� ��a��ʙ��M��;r�q�]}=߀{^�ZH8a���fK1E���V�8!x7�Ts��.��R��]	'��vHef���T3�n8�Y*|���*���rV�K;�IB����-Y��> 0t3Hf��c�9{�b!�� ���[Hɹ�H�<O�v���6�X���w�u�&܁����jB4E�[��f�6�D(9��Z�ҝ�r��dϺz�0�e�hq.e�b/�,�p�D��J�#�3�_��M�9���0X����y�u�T?i!;oS/�E;r )g���Rܤ��ٳĞ)�>g�A1�Ԩ��=]M��۞��ѿ�+v'm�n�#;��yp��s%�H1�����;ۖsoz�KQ��L�D�뾎��_�&'�u�9���WORE�o�w�X�t$Z�����6(�U�����<�T��ɂOY���y��w��j�r��zq~mڧ��_���_#�(:�
��S_謝#�)C�����*��n=�F�;B�����E�O@H���a/��l҃�*fZG�*��;E�0��RSXI�p��|�qN>X����V�'(6&3�G|C�'-j_��	i ǖ���r�u=�6`���1ڴ��
й�8�η�%��Y8��V/���D e�$5U��W��Q�r�rno҇��;]e��T�8OG2�a���IDc�@��T��A�)� ��%x���TJ3o"�=�R��4���Y跔� ��=)K,l�?E+����&�Ȥ�Qf������s���X�y$��i��u���&
΃�Gm���i��	�n��s��ª���R^��Z��Q��ݎw��s�
�.����xly��*g���z���B͘�:d��|��};��s�ʏ7�B\?�a��=�2�i��q�x�ha�^F���崦���0ΚD`E��9P�B�Y]N���?������hA�q��Z�n-h]�&�L2�z1���h���W6��x6�pY1�_yZ��Jm��ƚad��z��t�������տWh���`v蛔����M��Ea�v��*oX�6:3���R�G��͋Ot����zKd\��%�NvQ�K���ML�>��}-�⥆�c	��+A� �����%�;�t^��x'B���K']�.'���ؔ��ږT$�c���'�&j^��Z�:��R���M�V�x��o�	��65YA��ӣ�y�R�$¥�I���s��X���G�F`,�>TT�a\vl�����z8Yy�Ci�f�s<�>ck�d+N�Tť��4�t�`�I��~eB���HM�_�W��B*����K�� wv2{�b�	|e�TH����y��Zs~�|�M���²l*����_��޲�k��c/]?�y�݁����o���Ej`�Q��p�+����D5��R�2�=�)��s��[}�����r_�GG�OFo���v�s���������9��N����⼈`�_c���
�ֻ���.A�V��Ʋa�et.q���U�5��/S�f��&e�7$�\��HY���iB*���(�O��rڱ�̣��y�&�3*fX?�@�7��܁{?���E��.�!�.�\%~�՚�+�F���h�$/kK���%Bq���]��a�+Ũ��zR� 8}f���:aI�<�c$�Q��j��]bN�|2�&Υd�wv��r/��X���Q�Þ�#�*��bg�d�"@�oFY��	���@��o���|&CL�WhCj�Jbl��r��vh2��L�G�UU"�sed�?��i����	4�0����!x�j{z�OFW*r ��l�JG��^�~~�g�%�Q7z��;�・��vP6��^�6&�4�)@q �H��J��7 ;�z�07,ͤ�y��I�_v|��\�w!���l���ܙ��o�h�1v(��0�m��2��w��?��qȇj2��a���A$B�t@�H~mV2�(d��5�,�pJ"q�=-��l�9F(�K��٫k[J�#c�}f{fX�x�v0P1�d��+%��v[|��a�Q�5z����J���/w�H��c9�D�/��W�p������?q� �16�{�<{C��!�,�V���Fn���4>���7����f窸�`�W�����4����yu��C-����9m��9�;�d��2�c�s�Z\�51i|�x�KR�Us������h�$>�1X� ��A_h��G;As�>�jC2�\��9���H�"�)�A�L�*���|hU_	#�w�x����h���þ^7U���)
jDC�[ʁ���٘�r��CW��'�Y��pr���$hr��+�F�9M��7�j�\5G�`���)�mO����te����B�BM� <�G�y�!��w~���Q9=J��|���l4	J% ��>�Ϫ���ض�0�Eo@p���̣N
J�tY�>u�c�b��zi�C-� �I�L�X������ZӼP�
�%���Lk.��|k��6cۀ#k��o7�fҳh.����^V^����)�d��Y2����!����U�r�|N�Ŕ�/�⪀皓��N�wT�T^W<� 7�c�eO���b|p�!)h��"%����y��9����"�o�/��Ybҥ���A���do�x	cΎ�$T!EhMz�r���vv�d�B�ߔ@�T���|ܚ:�f��kfԥP$��F?����wp�6��L `$d^��VB)d�BSP����fuyj��d�Yٌ����}���6�c�><��]^���^�,�Џ�g���,R��P����_��j	H_-x�敭�Ε���S(/E�yb��f��"^�	m�9돫����K,l��ZJ�l���sgl>y[��s�7�6/g�S��hd� ����+��������TE�~L��CI<��ōU+`�;�qn�O@��|��8TU=���J���
�Jo[aQ␢�z���כ�]p��N��T�=������ ��
=���8_�peJܸ�*���c�	�al�^��O��l���]��դ�0X����\>m%v���coJA/�B�~���~�K~�:?�d���A�"%�گ�g�
+TJ�ɺ���%�<�u���ݔ�!W�PU&����6�L�N���p�5���a�uϵ��c8�Q �J��A�t=|��*�+���m�Z�#��,�/���)��?[�8T�,K).��v��cz:�`l˸g�����Z�e�f ڐ.��m��
;�>%D����oy>$�� \o���YK�C�.�*������Q�`G�*���u���(k��)����&9��kxp߭Jv��}�]�uj9�n;>��"2���ЭHƥ�R{�1V���5(oS�t���.����<!S�B�G�/����w�G׸6O�e��E/V,a*Ɉ-� �W�=�������JɱW�n�W� �eR��Q�J��Ly�����k@�����ñڙ?.b��u:J���W�h�	��"X����{��U��n
I�Qk��^�xS۲�`e͘��c)�_0"h��I 5`8��	
�ԇ��m�0\.�Xh�7T��(��g�Uēb'@�ڂI�ԉ����Q(�x�[����O�	�����9�x��)����P�=Y��8�ʨ��?!���R�VL�c�J����B����������]���P���۾pѵ︧L����<,��2���\ �b_4�N{���?ײ�!��T!���2�7JӗvoB���%S�	�=ft9[u�s}X9�n;R��l�i"f��-��ޗD����s;b�f=f�G?అRt�7G���Ӡ�*���]W����d�
l�ey���wH�sԑ��#�� �̄ͥ�纫������J�`�tr�(�hʝ33{�x+�x��2�gs��\z5�5+��<��7��9ئ�EݭA��r��_�Z�<���*~���!o�s���4>�G��)ǁG�
��7D���\=5n0"	Q?��C'�
���C�?lSg֜3��1Z�BRJB;��Ӿ�^���Zهq��5���h<vT���T"t�h��zc�!�"!V%"�P����=���E����}�������n�G���K���9��s��I���P����t.�P�z�nM�O�N��f��\/]f`���,��m�����Ke���	)^˘����]y���)�H��k�*�kt�~�o����WuN2�*�=?rnc���8}�����8*�;T
��lgv�n��ad	�d[s	�@�U��C�f�������G1�&�3����ڵ��k�_H��҆��Kv���[o,�����SY=g����٘�:�cxi�5���븪fyT���gGV��H�q,/�V��E����6Y0��#7�ޥ�����D�|��ǘ�jVn�VK>�����pd"n?_%���.�z��3�����̈́q������M�"�A t����,�+����c�	�>u��9k��`}2��b=��5���-�=��8�!��}*�.��/�Q��>�����`#u�x��Sxdxߔ�oX��C@6����!�;��!r�5�[
]�Q��6&ȩ���0R����ĦSuv%^�AaYN���n�"3h��ZY4�v
>��c�=�����+�K�WDz�[�/�J��]��i7�p�a �޳����;DF_v&�<=�>��� g��F����˧�)��n��<����m������g�����Kf\�i2U��B�����x�d���r�T���"����Ъ��$��7�Z tzČ��E`�Em�09E��.V�t+'o!���egO�7�YAX�����]��`�{�^I�� F�r�6�����X�B���E~�O�{(O*ɬ@x�fN�9zL�N�+yK�EWVi��L��k��K�^����oF��l�S� �]�5�ߴϣu��E�p@��>ܷ_�0J�h��O�Ls#��.	�E�hlM�k�6�(%�s]"{5�V���7Y�7pm����W�����I4��	�o�]^c�R=���	�|��{\�*�K����O��:xLi�����a 0����$�I�MR��aF��,�{3�j�/jؖE�N����M�-���!>gPU�8�H���K�e[G7�T{׌H���2RG���i����RPs�����A}�ӿ���2|7�ZY��ځ��c�/�~q�Mk����V��*F�Xg�/3����%L�w��ݽYgbHV�5P#!�һ�(�'��,]���]N�ֈ ��J#{a�r�Z�h���I�Y��zw�LD�$Km!!{Q���;�����[U��	z�v~��&�_�T�����!�M{������� fݨ�Y�̎�2deY��D�e��p$��uKޜ��I(�YO�_���_M��&Q-SN;gɽ�5��v���i�[{k	`1@F�U���[�˞z��ׯd�����R�C}��[�����|v�����=�I#��ZPt�Z9Ê���eW;sve���OcDtL,i�m����q<SEt/��!i��+Lx˃U�2N}2��k�!�\<}u5�Įq0h-�M��-����
j[IH �Δ�������J�]��a��v���%�E�Օz#�i#	!���xU��Eo��/���pr-\��Ft6��;E�E��G�-�ɞ��A��V��c"���o<����ʹ���#gW/�=$SB��;f�E�m)�nB�Q
�|�3H��n��8�j�}�j%0q������?S��#]E_�L����1�F�����CtSю��4g��|Wef�����E�=�5=�r��(��N+�3]����h�uz�+�٣�wv����5�Mk+�8��!�_d�/�]��c�����#*�xZ��LQY����X5{���r��Q����t)���~�Y,�#�	`lʰ��ŕ�3ww>���0$6��+jԕ`�x�GK�$@ɮ��1��/[���s=�ʜ�:����)A�n��
�# vA��w� a���Eѳ"0�xXE�g�����Z����2���Ud"c��#��A��?�����{u�h�P]�$X��>,�=�$����U����t���:�V���fuh��eߝ��CW��
�>��o�r?}�,`Q�ٟ4��b��JC.TH�M���^��{C�𣍵��.��1U�S��U64�s�`W���[d��H�pmA4ӛ��7��L�s������{YrI��ףBkӢ�g]ݐ����
dW�Ĭ���iL��+��>VQD;�z�Lq�y�9굛�l�G�Ba���W��J��E�������.qx 4�5 �K��5/ ]	}?)"�������� pZ	���&��9�~;}]25���X�(��
y~(��f�$�H�����'̼��Jn�ybQ=��G��~QX��m��6=y4�Հ	
n���)�X2��dGZ��"ǿ`K�8�ȦR�Ec��=~W�G��ȅqW/Ӄ��p�7�[~U=G� ��3���ve5��R>�>0Ox��Z�<5bض��~�x'����������k)r��8,�J����b^��k�&��\�	YH���)������IhlMHS��;Fo� �lf�H+@�U�	puO��>e��*g�/�'PCN��s��k ��nE*�ĵ��\=�a*�n1�~�J��Y�G����?���l�,�[��L]?�VY�}�S�b"\8�����d�kH�=���Щ��`��s���6��!���^�VJ��cu����5:�i���]dn�:���/��j�������B����B#��b�,AL<���l���7r����A�*�5f`���4�E-}�������V�,f-Ӻ ���Zq�;e�I�b3H����*��H(-�2�S�N��xu�K��q�<���<�����\7=