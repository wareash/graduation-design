��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf\�|Vv �q��PNc~�eEث[�r�ٶzsg8BWF��te ng��;���NșW�	��5�M8\��ʋt��«]!��f"EfL�"�j�W���"oE z�S�vӍ�cx�Ϟi�'��Pu�!AY`��Z<x�w�[����O�:���Z�����rk��z���j�2�������Њ��tcp�h�N�-���i&*����i�>4JK�=,)�>?�����Q�Q�S,��}'�δ)�`z�Xn7V�à���+=�3J���K5H�b��g�x���˹�fS#�ꅨ�w���eL������2̍d�"�C4O��-\9�6�^W�m���AI����1�?{�`��:�׈�ra.2�Y��Mܝk�b�?C�V�	4\�2vc����A��@�?�N��h��,U��D��&6�	��ぷ��py8�#�-�~�Ԣ����}3�tԬCl�SG�ـ_����4��_h�V�c�b�y�|w�T,x��, ��*S�GfΠ�(�Jr��w�9�CW�f[�\�����i��_�/#�r��m�Fn���&N��:������ &9?=�A�[�	��1��Q�m�q����I�K����L�����s���{��o�c!�Q]�:O��X���CC����7�+k��M�_���Tj�L>�0��AD�N��A>f@����߮�ϰy����'9��>ٺ�B�Q�U��n�x�g�������b �������S�����C�.�W��t�ũ��a���: �t���q��wS��_'�e44\��`gf���Z�4��+��:�������v�%��=��w��>7���t����M����I�rt���A����r��p�2���%V��ZFr����_��p��jD�sӀ���O=^����)�j��U��[���z�h����B��<��)G�HS�ƙk�`��{��D�Y�F���2��%XB�a�!@)���@p�`�\��c/F�ؖ���v@*g�\��Y��@3h��2֕nd���h�X�)���JU�d�4e�r>gV���vЕi\~�Xv���ȼ��<�!�z���щ�݀�#��NB�_s& �S��z���A�P��<Xs��"U�������d�GQ�uE,��-@�V��B�f���}W����x�B���L'~
$G�˟ݔ������M���0�Tb���{�Я���?&�ǫ��(�R�l��w�R�M�3�X�.C���Qҗ(n�ywf�Ck���OazX*!��gW�0^%e��c�S�0�af(��&ՒF}�WF9C�]����0�\���D�J����8���$�J�H(�,��#H��þ��K��lO'�M��6�2{�9�c�S߳8�~�s�֑<U3���/|�&�Y{YX��.����v=��ɼ�-�e����?�*��Ɛ50w "���^�!�W���5����|/�Bbs���>�9_<b6��cǐ"?#丐�k�<גOF��vf���Z1g�\��1-繌�)6=��؎���-enLL�����%���\����mNJo2(6��qJ�U��#]&r�ww���I-��M,�K�>H�5߽��*ҳ�|��7&��(k���+����@I�����V�� �:���4�����:��>�դ��M|���T?e��}�ځ���Pz���q��d�M W���P�%����cy����-3�Vц��Śl.*-�����?���&1T�ْMm�6p����O4��0^i�T�E�>p�cZ�җ�����Sg�a4~�ه����a�������C�-kr΅P6$�������T.*�f?��y�6����g�[G+*����t�Sp�ū�/3Uf�aSH$�6�
�s�J�#�ad�f�lI���x�I?-���wÜ!���u����ȤW�yH���\*���,��0��j�L��E�!k��̈���%�ޥ,�'�	�]�A�?-D��es��֭�KҴ�U����m��M��^B����yR{+E�a����<��q��ll=#��D�Ԃ�*@	��^�lU���~rZ�$��@XǵI���"�{�(ۑ�N�@�jVQn`�t#s�I�C%�0G"抽�{	�-5(�k�h�+��p$E� 6\n�QX{���W��ֆA��U���ʍ��V�jߐz��w���Xљ���E���cw�dNV�a�����s��^,;��f�Q��#�K����h7�D���2C|j���'Ƽ�LM0
�Rp����r�����g��VW�=9Fy�k�n|ÕҪ6�����N�E��y�k���K�v�\����~*��Q��d_Bh�9���Z��c7=K`�RR����ȥ�-��L"1��iI��a���||�F��+������Q��Qa�p��B*�bV�U���<�T����b�Cu`bM����0��=�u��B:���Q~(#]�x\	�k_��G���|w?�AVs�V���(���s2ꌭ����ݴ�`��Pmo�k�Ϸ-�"1�k�	���	9e�󒿏g��+>�)��	����3�I�V_;�߮���xe��8��^�ĀE������!��"ܯ�%n��eO-�"E�@f+�>�X!��Ԡ0�cJ^$�$�6lc)��C��8���規��TH��wY����"]�
�F�Z�(4�Q�����ś���Ps;�5��a���}�4�a��[�s��sC/�rO~y;��Έ���dJ�Ge��u����܆.j�x�^Y�n�3q�&q��G ������z��`ĕ�j'���������:Fkv�e~�X��� �!_D@
�΁�? }��d��Zy�)���uD�w�ϵN��>��8 ;j>�Xҹ����a���~E+��5����J�x�mL�EC0g��aV>���E�C>��4N�n��v�U�a��UU�ڈ�,�t����n�Oﶎ9[dg\����cҦeߚ�ÁF�ϓj1s|kT����G�~���F�Ә���
�
�#k��f��H�F��!s%-�Z+��6�(}�[o�E�>+cf�U����mB8�׊�ycsZH����A4��z-U��E��$�/{��H����
���\i�ǾYV-���¼]׊��ޫ�M�;}A=ƈ�#�t�8����A@�pvv{3S#},�e�۾�����;���"@��ɟ�(��z�g����*��OF0V��{r~֝{��ǅ�z����� z����-��7����_Q�|�~�p�Bﺟ3��Z�7����s}��:�2J����T�LUiJ㉷N��HaQ�[�ٸ�L�|�;���&��LN�H�`�tu@L@1^X������5w7I�����Ŗ�UC��*�52��N�םF��M��eґae-k��F*���5�ô�9$�n֫cR1�^�Urx�J� L.�4���όwWӖ`�B�C�x��������	��g/�9��9I�^Qe�兌h� ���$�ؚ~m���H��ڍ�~1�U�=����2��́zr�ʨ�^��_������Vz���U����N&����R-��'��k�r��T٨s>�v8��P[���� �HU��`=>~ �_8�	�I����j'�ri��� &�C%�wI{ך;���k��0~��+�od�	3�K�� �����N�%t��q}�`����E�d����S;*����|C߄��>&{�/��AL_��:���3�`X*��":��I���c{�����#���9F���o��e��RW���{��O2�Z�Z^Pl�U{�P�l��4��)X�����AZ����=��[6�f�'L���$��q-�,c*��^�]�m4����GjJ��؃`�p��ryM�0�4���j��J@��R�g���^����Ɠu�#s�y[i�O��m�� �5����a7!ѽ ���\����.�^rν�9l�M�I+c��U�s*iP�$z+ ��m&�Q:�\���߶�� ��--��a
�j`]X>Â,� �!AeU��8{0}*+�G{���������譕ǅl�<0lX��(�XwPu�T��s���K�4�,�!�D�ftk��_��լN)���o)"kVОd�/���Q�f��\֋8@��I����;T�k�w�0�D��fv�?w^ݏ{C�!*�f9��3�K
��3[���C�}��6�8���y�%Œ5�q����EH�@�&������[ժ�w� Ǟƪ��46��u�Ě ƲO���)�,h�(�����.�`g��D�d8������[-���lەˊ�ȩ�G�z���諒�Q쑗�k\��#�v�/Éu��a9&������7�X�i��`:y��(�|��̺�z���kO���4�-�R8M�%���.��񥎅���*A���_)�I`��(�;�W����Kj_L�$�����+�"��sP'�EG��FC5v�{�8o3���,� �0�M��$Z"��߲��T�*M���K�
 ��\b�('�W+�A4.k�]̃�d
�YXK� �)LF�d¸K�M�� u\hA�5�E�.��T4�J���k��]؉Y ����A�/�?�H���O	��4�c���H�pB.�+d�H�>����\�B4+Z��ᗖ�fw���%	�]ɂ��q��"br��@���U�7��9;V$5_u.��b�qWq?��JR�ݾI&�n�.�s�,�Q0����d�O�	q�֙�È
^��b�8G+�޾f��S�)��
o~bx�!1��ǰ���yf��B���|�5o_P��e]u6�"�`���'�@���8����0R�aj'�X��Rm�*�(-"
:�\]��g���4�D&;�	 ��Y���\��(�O� j'H�b���V}iU?K��r�}%�#V\�'?ܺd7�~�s PǬ��0�zu��fVVC��"R��j�����T��Q�pu���%"h"�O��Da�h�l�R���qI�ͅt*�+�ȎU�Nz0�\�����d��;(����1HJ����U�Q��dE�a�-��� �>��_Q���3��/������������_�U�����i��Q�o!ФQ��� �����w�������[��V!�&���	���,{2��D$���*N*5
VZ�����v��j��_�z��<L���/�j*��G�'W�*�0������~
��ۇ�*HL�#�=۞�Kc�I�^4��Ȧ~O2<�����3`D!rV�����N��)�`�`: * ��"��i��'@��R��)L�_�3�O�RP���r^4�q�����U��1�K֒�%Q�����N\�*|*am"y5���q����/��6Z�#�ǹ4�ܼr�p�f�hM�$S��>pc�[$�ԞR��<	�NӜK0�b����f_����䆥�ڋ���8��yj)�}Ϝ:�:����v����0l�� Sh�\Egh�5�����]�B=ͫ���*��8�X�(�� ti�b<����f��:S��q��IS�#z����^L'�R~�}�1h	�o�+���3��|�[��soz�'F���g��sd[}P��9:q���ԛ�|�Ҡ���6�ڨ m�x�`�:�Dc�Yk�����Gq~��G�A���,$AƗ�D̑����~V�n;6%`{�����S�u]#=�h������4�.c\r6�l�:�tZ�U�Tf�����rK���/J�͢t
O� ���ա�y׮��Z��ڰ��ݫ�+z(�!qe�+�|?z	�p�F��Q�4�d����,9�h{.��� H��7�BA�G@-�n4�s��YE�=�
/��`���<EH�W��k{�7�ZB(<Eݗ����p5`y2�T_��;�K�ѕ��8����r�ֈ�'Z�|p%�u�\m+7�a��P�\s5y�#�ގ�iX�'~�D�i�t�͜�uu�ϞI2�Z��"q���!���\~a�E�P�5e����;^^
$q	d6�@1@?tIi�~s�٥���$r�O�	��E��~��tfiC"�z�!������SA�D�D��̏�#�)��&y~������`��C�T�<JC��=�	<4�B?>1��UQU1WR�!>x����^��Jq�e]V����m瞓y��j�@=p����b��f_}	e%� ����~�\�$ �/�O4�>��=2�|K�8{)�o8��e��� ��N�<���lK�)l��A5�+S臰��Dܝ�\L#eT��S�g!��4�����}5�/�(�z�F�
�Q�r�9D����R�_4w`����*H��	�=�r��®�՟�����,������ ��;7��Mqx"�]�U�8t�4���n�A9��i����1	�w@U�A_[����^s/���UH�/%8Iv5;��ަ�,�Uq�w���>�eWo-���Q(�i�7���B;z�7Z-c�,��rn�Zʛ�	��۟<v���IWֵ�e~��a�e����DY�nB��*�T"��h��dÅ ,�xp��q6ɴ�L�"�Nʶs��K＠Nմފ�Oz���O���f�t����ѓ�nE��`��N����~Z�ql��[�n���Eh���|�H�����F�[M�_i��>�3�ؒ�e��4��N-���F%�����z6M�|�a/��4�_$?n����<�&Gz�a�Bg�,K'��K</�g��{�������P���#V�E��M�,kmY�s��Өu�$�s*�ܬLv럾3�!J�43Mm�4%�N���X�X�}���_�kx��2�0��E=7")�2�B 2�PiPotp d��\��|�I�{�\�E��μ2�Wԍ#_�R�Z�%p%��S�������8FS�{��)4Ġ�;z����/�s�X)��ʑ�a�D�ۢ,7�	Dr1�I�BÚ$p!��pC{d�@Kj�y�2��-jk{N3T���!<�z�����I��k�2�{Zv�d^-%F�{Gڋ�\uʖ;��2��FKMz��L�'��i�yPԦ��	��s Q�/
2����&-��)�p���lRW�[�^���5��Fwe>S�;?h�a)KI�[��t�26��;�~~�jr���LG�
]�\<53l�D���N3�O屆ju�e<��dn�-���`���͠�}���E&�0��vAQJ*~�lَ�-�R�UDݿ��t����:1GT*�F�*�)M�J�Dɯ=���س�[���ƽ�+��dq�)��aH�*��2����&B��+�7B;�Qn�K���eS��� Ֆ�n�.�B%[]�ie�sY9�\�d�TZDʯ.B��Hm���@n�m�;}��Q�}�@�̍�d��d�)6̗�+�A�#ٱ*�H�OCv�֕�M=�hs�xα�����^�0+�f��v�5���?��W��H��!��Z$2��8�
�p��w!��i��ذ=�c]��?~�Γ�*(��&к%�l��<Pd���?�>��:�$�vC�{�x^�4���x��}�D^���H�yvPi���-s�e8e��[��R ���t� ɂhͧ� �bȪAH�-z0tfb�M��7�Tl�R�bxe�t�=��q��W(ɸ,|�7'�0w)��h:!������Ŕ^%�k��l�lv乳�{��`c����E�'��(x��GM��l��~�N� ����d
���������ic��q�=�j�6��V[����`����C�E=���o�����H�p�s��/��:1"��^����Y�*>���t�B�j��hEū��-m���]ǽ��5s8k�D�R�2�T���B�pb�
��������w��Z��y��J܂C��b�����5a��-�����U;�s�BVp:�&:v�������*W����T��c:���&cb@u�КL�΂
-~��8>K�p%�f�ϰ����Ijjw��|�(i��v� lCD��]���_�F��)�;�����)''2J����S�~z«�'�n�|6��%�������]�4�N���1\V��1p�zhY)���W��*-���0�,���ݜw��<������|Utl�@�"+�K���ʆ\�<h H���]s��O]7�0�5��v��0�
&y׼���\;�
��ƽ~�E=�ު��(������a2��Luśk�o�N��p��^����!4�/�0�m)��Rw�wQm�k$�`4;��<��b�,�F{0�FD��L���챔���WiDe���!m�:C�l0���j��¸>��( !�WC�·�(����K�"C�l����t~x��?��g�GZ����j,����l'���z�%� ;�+�b�[l�1�#p���޽���>���/�?=u7b׾Wݿ��U�FZ"�qV>��6ݡ6�-�G��8��L6�1�@ km�G��F�[��歇�[�T�L�d�W�8��r䔌����=UӴ��Aӫ�{����F�9&cYpW��������n�P�vC	���y'h7I��|��q|��ѾԲ���].9�+�nI����RZ���m挼����+C
��Y��j�����u�[�|�b���yy%u�]zDO��9h����
��ėV�AS�{�qߞ�s�=�EaC'g̙d���V�#7��(dCY������_�[�Ec[��oq_��]B?�5$,�Gr܈D֚��x�Y+��e��c�!��U�8���!e�O�{��w�(E39�ø�G�e$d�KN	�X!hI�Ǹ�fb�^�P����_���S�x��*�V��E�zA��1UK�W�K����P�"N�0�9�����[x(�T-����)�����}���B���qB�2CX* ������d��ܙi==s3F�"���{,�@��=b*��o>�,gxq�iH�J5F���#n\��%.��r�=���X'��/*e�v�g �3��j�v*��,d��¶�(�<���1l��s�:�2���s&h������/�+��Su7:���"�"N==�F�H�OY6"��0s˽��&T�����TR؝���vY4E55����՝��O�0�*S$�V��c �ɶ�^R�b4+;�拔MO������Uǌ�+r�'7�h��_���bː��6|�k��HX������CY�ӀmKl0sb�gѓ��Y%+v6�#��o��d&���f�����乜��B@�l��v�i�i��Qe�r��U>{S��x��a���Ml� të��QS�#]<��Ia������p�&I/!�����d옯3}S%,���=V��,�ҴxM	l~�7�I<�W1"���f�CD�θ��<������Q̒�wH�QY����9N>��j,�It-O��(�9�nǯY�>�T��9�EA�!Z�B�fn�.J��(o�^|*@�����۝�!�!���)�L>m<�R��N~<9�_��I˴��
)�ө9ϛ/K�dğ����ZY;Mf#�o;�My=��-.��)i ��ݲ�(��W2� �ͥ��񢖻��H���BH&��r�:�"#Z쏎�� �˟<��A�$���X���<����f�~�*x[�r�"A�	�( Պ���\�5r/O�
0� \ ��]������f���X�ۅ� ��x�/K��Dh�
L�L�����%eY�C�ab���w!)b�<�ê���ډ��)tݶɿ$�S
{��#;��*���z�rm	撄5��X
���?ɦ�%v�B�@@
Z���՘ˑ:(��r�m���ۋ-^ҚP�;wn/B7��"��dT��������=�Ċ��d{իy]������s c��6���?�yW2x�"�%�<Z�Z�UaEM0�>���^�of����p��ē|l.B������N�.�'�Uì�� �i��'�O��� �k�wn��A�����^Tx�66s�&�e ?��f�Q�����0S���	r��*P?�ժ��p���A�:5�ؒ��X$ZU3��O��%�DEfI��g@Q�L��/	�S!��y��8Mu��3��:����z�
�;a]z�@����i��q	p��V�I����*���x��yHŮ.�wcNb�,?�ۋ�4x�7�����c�YGU� l�ӥ�r���f�0�=JA~����9?��һ�b��y'�$��@*�F؄��4�T)��c-ik� =(m7����M�@=�]4�4���m>��<$�)�3MVAP%��XI=[�Q#�Cu��9�����I1�yQ��	�r�c3��V�⬐�]�����J� �΢-�����S�(�6h�vM	�����hS0��S��p�����47��uX}��qv������~��	�o�5�`�9r'=8�,8�8�~d�(焳<��::�<+D��2�I�;/�c�9Q�c�S���w��n�ZE*��!�/��ø���_a�u9��h [!#��Ȋ�R�:��{}�0TS�$��e�,<% U���,�-�,�z�n9�;dHeА#D�����#�HFۼ��K��U��'��"Z�=kcqg��3���F�M��v��ě+�+�FOO�^V�71j��*�QU����{E|޴�_�����[x�R�w�ڏ���݃�;�s�%%�g6�%����@,GzHq��J��ߪ�ٷP
�t)Ѳ���p���`��B/�b�)���b��_l�Kì�v�f0#��겗Y�F�N���Hqq�LT	&[
wݛf����N�EW��c������W�az�
>)v�����.@�����]C A����ҭ� |`%��\�0�'K� �"&_��<�8��K	�
�ꇥ����6<�(sx#[����1�_���L���!0�
�[>l�i��1b(�A&�^��]m.�j!��\2+�ij��B�̧�H�� �dJwQ�e�YkgbWT����"Ĩ�\��oR�=�P2=젛l���N��3�A�ӭl����W��n;���㬫?+܌�B���ڤ#	��l@�� ��H9���1/^�R����ipc~�ާRJ��b�����ʀ�(R_�&�䭌"�a:���@o�@"x����7�H���@"�/������Q�
��s�:fJ��ȿ���
��7N�"F�c�_��|��'��4���ɃǠ=\ͷ����Kh��S�д�`,1$���6X����kEK�`w��վF����#p�� �ɲ�z�'�V��S���ݪ4|�mԆ�-��H����/��+����cj����Q^�
7M ��P���i�-K�W��n�l�~�Ik��=h�N9���1��E��OOs�Rͷ��fa����#۞�C��qȄa�vR�5#^z�u�9�<N,H�RV�⢊$�F����wx�"���@@$��]Q[T�܆6,��YS�T�5�%cOL1�B��a�OD�Q�pLg\ƙ�1���B�22��ٗn>[$���A�e���H�n!B��̀@MThekyO�`��*g�&9>�yS'B�%�|����N!���ܿ�)�'���Sj'@x�zb��Y�@�-.f���d~37ѕ�ǟ�PZu����\��5Yj?�e���V]��#��H���bn=S�*���8�P:�Q��#ޒ���� ��B�Z�+�k4�u��Dwꃤ�u�ĉ~&�c�h%�������1�{˻����u9�.J:q��~��CD�iR����G"L���
�[�k�c�~�s��X �8��c���
F�
0gE��kZ�[��i�2�qB�� αFԎ�gls�Z���U�,�������� ��},���oF��7�A�T] ����N�ڤ.���!CE��Qv��W��r���w�����gġ*��Jּ�*F�Y����[�ݣ'��U;B�㎾n\���o�8Eb�1� Eߋ�D[�E[a�CL���߾��%t�E��� '� ��;}h,���h@(p��[ʆ2,��x[ֲߑtkgg�{�ض��>)H�5gѺ�Ǽ��ڭ/"j,�ZQ�Z�:����$�6���u_��i���ŋ�j���4z(Z��;u1�l�z�H]�'�ؼ�֑B�Ve0<V`m��u� $��=4;Rq��wq�t�z�R�d����ў(jB��]����U��(oRI@��R�=�^�n꾘z�|�;�_W�k�{�@]����bxq�&\���rb�.j�_a�0�zP�֓y�5-	{�-XB��}��W�^��h"Ǥ�.x�Y,cC	49��"��#�|߉n�5=}�;�-V�����AΡ}kc�Gtͱ��yo	���2�#����)�5z�yY?�>$���|a�u0[gH<���$(�Ǿ#[���'�/��l��UE!�v�c�nK��@���lo��?�)/W����Ib���4")`�ī)����w�£�+��*!�����Jv\@��k"G�r�G��8�����ebC�y��
���I�G��4i���E�YQ�[�T���Ę2�4����
m,�=u&N�^Jٝ����f��s$�Ǟ����3'���&	u
�:\{�ꏪ��'f�*7���w˴*�]C�>�'�Jt�U�+�<�H��G������M��^�PV�U�W�f�KE�x�����1-�H���P�ҰJV�l�nD���2��"���K��}�ˁ��>�B~J����b�c�z�ۃ��Q�Rq�s�1�y�&���
�z�f�rȁȔ���9�� �A�_pL���ťG�0�z#2���wx���׼��	N��ޘ�|q��P��gc��u�O��p	��R��������_=��R�Q����<`�{>�.�-�10��� <j�<`m�`�$2<�B�&�	�E�o�}�D	���'���BF�`CE�+9+]��2ܡ�\��3��'5�\�����+U�^�E��)�� �YApo�cg��F$���^x�mذ�Q��$��Jjc3�u�����H�{�jA#ek�hN?p?��N��I �@�6�7���Ng�`��ܙW��#TK����Ř\]��F��C)3�'�sSE��iX�ZeœY�f4�����3E�S[PA���dI�t��cH�I\�j���F�@���5��n/ ��+�9�>�X��dlD��DU`{�/�օ��8{A[]X�Yb�ڟȧ����=MHX�ʃT����>j�Y�u�5���d�u�����Md�)$� �i}#���8�N��rh��!u8Zq�r�U�Ð�}��ѐD�9C�)6ꮜK�]�hbTK3�!=�-�f4؟OW�q[}O�q3���p���N���������x*�4��,l͸���}��C��Q��T�{�C��K}|�p�,��a4k��ʎΘyY�A�	�V�,#=�N�ؼ��l��^���g�\���y���o�L�!�{���0������.
Ss����zb5:n	�E�d���n(��ׂ���
G�1r�=��1 Vr<�馥�!���=)�����]�# @�M>p��M�����$T!�L\����o��tٰ��T�7O�@�I�X�S�3�l���F@<�)WboX���AEl
�iWp������6�;������=���t�����5�[�v�����c4��"x=�S��?�I�RS��=��N�z�o����H	�P��
 �e���C��{N�9֭���!���9�h�w���,���:y�2BG%�a���!x~AǓ��I!��n���O��tCVHjD=��0DI�+��Uu��K	��<O0w^�vm������&pz�S�|S���<���R��hZ<�,cVS�4�񊽨�8���"��q�V�jnQ;�M+M'�T3D�˞������3`ʘ�i��)��kzt��d�1{yC�_�b\l�۵^��SA���T��H��1�ca�$P<IN�I�|�_ m��W�8�'v=�������3����!���xA`ǡtH����#����	/�f��p~���}}�A����@5�-{�C����`N� ۓ�֫�+D g�!�e�	�q
�hÚBq�uo�R�|<s�iY���2�"�L����f�>�˥׷���!��1,����z�!XK"\� J��]�A{ޫS�Z �+��)��_�	�;x"R{���uЭH�dg\��Xed(7i���Mhya>�JPD�0�M�V��d��K ��Eg77�@M�Km�q/^+	�}��Y�~�K���K�N�Sm�;��c��w{%9���{TS��M����`� +hO/a�я�6������7L��0'Vm��B���
γɩ�)�5d������� �Β������IJ��,�o�	�6����V*��6~����s��Ҏꖫ�M�0t�I�=�QHZ[lx����	��`J�3C�� �(C"������L�F�z+�zw����3�@�D��TW4j=��b`fP��m]N-��IAm
5�$ٸ���������&�l[���<0�0ܱc\��3Bh\�:��d0����k��6j���`��:E��]s�hkF�Ѳ�Y]gJ�^T��\Q��c���t���Qq�I��&��À.��c��%�$�X*Y+�ğ�pg��J��__��۾��p�U�;�����3L/�׈��JV�\)�~DoR�-�7J�4B1r~��⁃Ʊ���D����͞�n{@�1�T�*go�-j��HpL�!T��3�uŎ���e?E���e"i�%�ڡ��-�/;O$��u�C'�&��*���;��y���{HKb���Ks)�vy�e��*7g��ڪ#GF��{����e�"�,eO�$6A=0|�x���_r�|����E_-{�%�?i$��`.#��I^$�z��4��&ƶ��=PVv�������t�PI�?]���[���e�[�8�3Fũ��ˮ	ئ���[��?���7��;��S@�h���"p4�'ˀQ�ʛR�dKz��ZZ=L�my)��H�TX�����>�U?���S���e���[��rOP��� ޑpKY
}�gz�o"�YM c�:t���)L�tR�Wq��MB��	�̵A��u`���Z�\�ӣ�<�Ⲥ�`�NͿB���NI�rz�gI(�#<�l� ���TvI���󙒝�*�c��9������ʃ�6͞��$��ˡ����M�1�GK�f�;êPɔ�����D��W����čC&����Z��>@����ز>F"�#(� �����r�uVG�%i�w��Eq��ZD�k:R.s���Ö���+.X,�S���C�"�=�~�N��V~��u�$�5��s�8�Ii@V�rI��:���uZ8+�봾���
:|°В(��A��F:cX�T�$Q��}���^y� ���ȋ�01����0O�\��?B�u�p���$����`ttR�?�=�^��<+�A���~`��;"& �8���Jj��!wz�f��b~,��G��YM����e�l晱][��
�nB���H�L�W�Ӊ�)�"_�.�K9���㺏�RQӔ���)}�/l�\�=}�Ga�9��e
�U��M�)�4c����	Q�9�H��?1��2zɄ�i���o�̟߬����X#�k����ȡ�2A��}���I�2�QŖR��l�v8 Ho��T�+.�7%A�+�S��g��
ޔ~�k�r�u�z���Tm 5��=
�hJ�?�ꜽ��q6*�����:�����BF!�!,r���	l�S�����B�C��vcŊ��Ō��^���8���Ł�������u�L���0_EE�8Z�p���B6#&}� ���r����v;]���B���#�if�iE��ж~S�)#R�j-�֯*�&O.1<ZBen�������r�����ϊ\��D�>�1��8��o�ߓL���m,���Μ<�G+3m~k����V�,k֯��k�J���I2D����9N�(ЎR���W։�Xi�zN�5��(�,���z�'pkQ_qs���������\_$�.�?'��=��.�ھ;UY�7\'�5�0���D�rV���X[��
'���ѓ�A�F��5�o�#����j[O"�+@N�{}[UUq[/��ηq.��0VB�Ghr"��E`���f}��K����푱Z��'��t�n۠�)�L��?'
He��3FqV	�0����Z��9�TW|�Y�\���ׅcd�\��tH�q�q��V�a&����?ί{�"z��x'I�2�xY%���xs�._��ϒ��4O�X�ϴ����[\���L˖~��r94�ؼ�fo	6�ޅ�Ź�F1`F�).z�����%��R��@� � �Sz��� Ip�`Sq���E�P��wհ��ܴ�n[���"�{��(���S�&k�OZz0�)��Q=w���e}�+`�y��_\�T�"Pw�G��]}I�����n�� 	�Sx̦��>puSu�#O#>���^��c���D1�݅D���I��{��n=��O��|k�!O/�Rp�Ո3A$��qc;�����|�;����	ӻ�g��+���ⶻ*�5d�jԹ���m�p/RY��!��KNm�|�PD�0
�a�\���i���M��Y�F�g����,�u�1[�� Q$��|P ��J0�~�Y5C�Xi�ò��`���^��������Mr�	�;W��w5Æ�*�㛨J���iy�8-e�xr���'����(�ϓv5._6�}N	�U�o��}�́7�Tt�(O��oD�8������p8`x�	�0'z����-�u,�ɥ֊F+�.'��[�;�fN`�����aK��`�u��|�Y(3S�V��O���=<��[3�a������cI�ev�'��%� 4�PY��NyHTJ���46 ����J��JB����̅Wq�O�\�Ȝ�=����>v#o��#eg��7kP��hQ�v��ZEw.�*" �򹺖���Ap	p���<��;�� �|庁~��s��d����F�+�"�h$�������ۃ����Cy�!��x�1ʜ�*��V"�2�S��5���%M��G&;^��m�Xo�$\�v0��3(A��Ur�6}�7aY�F��q�a�b�&L�c�� \/���I�7t#�M�"��Ba9<YW�X���J0����r�r�}��_�U�}%|��@�qU���F�3x���\���:;���4&ҁ�K	��(�d�Q�H��mo:j��Ȏ��y�0y�v9��������	%:��r��q<�:^
'9��g�7���Y��`���a��vͥp�*o2��t�P���6@���YF^BOȬ�x׿�9.��~N����5C}7R��V��6'�ͅ>[f(��y�"���>A��,�үV��3ԅ�$���U\��)1؞��h�N�i�mE��$F���_2f�BN�sH�"?�t.)�����PB��9��H��1�B��F--��-[��.o�f�R���yٯ8%+țF�}6�H��?����M��t>����|�C���UG�o����*�e&��0%W8����[��������p�>��ft!��A�>�U�{B�� ��$�~$C(/T�>x�6p�����~�&g�f�u���8�uJ��/�O:�Y���;��N�R��?���ه9:R��/ ��sν�zK%��3�Y/W�ggP yR�x��F���u���qN�z��X¾���ٹ 1��c�b�=G��R�5N�g2E��G�G�"�&ڜ
Ѥ�i�7�*Ԅb���3��+��J-�Ӛd�<��ּ��V9����:-4��
T �D��nɲT�2�z��|7ҳ���<Xԙ&jc����a:H�ܭ�`Y�@VZ��t���i�H��{k���������V�#�(�\��[Ӓ��9ᆎ���#��"kd�~T�nx86���$��R�Lˢ�k2߼�J��!?�2�qH����'o?eN�說e�g�Y��\�\�OOr�4���ߺz#���B���l0�C�#�M�����e�[kZ`Cd{���G�l���W��{Lsm]FqPJSP@��^�i�����G��Ti#��b�z�������GTK�R�I�HT�b��2�"�Kc��wi�!ː�Z0����e�lD����_�]0�ٕ�;�O��
�z��Vy|%����u�2x/��k���Cq7R�k3�1&����=��<�&�����R�+'"�Xjml���2 ѯ*�Q2�+ntG��D_@g�ϰѪ��l6�JL3NM��n�XS�B�j��e��T�fVU�>
���U���.��<���J�4j�L�s!em.̀Jݱ� �G!����;,���^-C<ExQ3J������o(DL��ٗ�����3��o6���G�P�OR����T�q�4*Hg��Z"}h!�b5`MK,��{��~J�ЈP�m��W#K�]����]�<z���t�Aضg���67�1��ܚ7Ǖ�����6��`Ʒ�B�ہA?����d��a��1hS��k�o�?�24��J���Cwp��W.Ϣ|E��Z�hi�<JǧqX����
{@�k�21!�����7�xaD@X�a�70P�	%|��l"��jp�5�A��tW��"N-K?Һ�O4�����c�V��|�������"��b��k>`1e��1\鉞C�\)s��9Z3��s�"4�����u�l*J�s�E�1�N��c Q�[e�����G /F<�R���o�^+���������Ge�5�4ymkG��81e��;;9��)d%���T�S�}	g��iE�
��(�ɛ|z��v���03'��s*��_r��YőBޞ�8��\������@�lDU��9��'^���``B}�.���[NHXM����W|~ߢ�e6�c頍rn�l�N*M�����9��|WAsDm�-O�µޘjC|@7�`"���,1��ڶ�� �]"%��"y6V��N��Ǘ��31�v�ݫI�w1���&`?CTq1��Ԓ��X<B��|{�(a�G�%������(�W�Ոғ)P� ~,���٬'�?S�:�J��A����_�=WHn	�z ���C<�;���$�l����=ǞZ� :ˏ�Րu���e���\��X�s��]?���u��@�R^�36���w'�MՆ�zC������y17��W�P����mڸ�"Oe�?�M�"X���㫳'Bjʦ�|�m�`L�J�X'�U��^����7�K#ղ�G�]_)�}lP-<՜��͌�w�m�j`��9߂��X����iB��BC��F-�`��˨����`�AtP�S�i��d�1�[�^�2��Wl�U� �(�[eɨ�
�^�N c���{cܧ��ܿD<H:^���J_�Y�Q6f�B�
%�~)@�E�U�31�{�D~,+�k��'�Eƻ��
�'pv�CR�4+O�ǽ+E�sΉ4�J.�y���T��m��@�N|�� >:8�P#.�y�I�eHG�Mʝ&%��N_x)g?C�����n%�I�A���*F~���f��w�n���Q`\R/�O�(��숰�2b�SxA��귽���|Bt�X[iIB�%�R�%x��^;CۄZ�6/���E^���	d���e�I:�*��ɵ-;/f��k̪��	�����G�Y��Nt�ie�bv-b�fUS*�m�{��9��{��ւ ,Q�^>�����mA�+��-<����4�cF�G_�-X��U"{��P!���]�1����t]	��Ǧ��,U{�Ӄ��7+P>jɊT����Z�yjz��ZG?8�{���R��j��&y�j��9�M����`�;��&�%�b��e�s��������!T����$��HN��t�����H�ܕ^J��Б�MA�1o����T�����Oi�!MT��鿄|2pU~��Ѭ�������%�@�WX����y:?��SI�XY�껤1��_�a�ۊ�^���f�ϊ�o3g����6��F&��>�O����Ab.��}�F��8ѻ��	@�}�\-5�ث�mKÍZ|��g��T�'yn�(=���v�1��A���0Ǒ��rՂj�~�Y�)�,s	}i�$-��J\�pS�t�.�[��Ű~����MzNw�x�����FG�����R�#YL3�
j��>�#��V�ȼ�w׶t����r���d�lb�;t���N�Q���� f$8�ӟ�|�/�Ǩ���!V.���Io�k�J���ɑ��]������ �l� v��a����DI��������KMd��8B��W޿FTy�|���ye�6r��\آçA��Ԇ��iEZ@*��(�F-��(����Ḱ]��\ӓH$%�*�ďX٤ +L��t.B��(H��j��ȥ�?w��=��e#ۭ�C�k�����d�l���`��hz��n��'�}�H��/��<����
���yR�QZ}����na�����1�h2�\m{_��L��J����=T6�
���$�n3���޽��y���f]���;�~ϪWK��f����~���F;fr|7��C���5�[�'�~��=��d�����1��P��'��]=!l��-�~�	/6
�PY��$cU����h֦N���R��W�k�$%;Sv��X�X��	) Z
�E���^��H~9�. ����\��]�z�#�Q�.�po�e�͋�P�� !ե��b@��������&/��MϨ�"��)5��#$�pZ�|吸���Q��qq���R��Ti��!��	���C�~���g��t������Ή�HL�O���}�M5��Z����=rЇ�~C�3�m�2q^9�.�w'������)�e�N�����ߛ�5��A}���׫�J��$��T%�C
0�x���{>9C���̼j���M=�?�2���8�� ˂WƸ�46��wF�s���o�c�F�p�] $��|n3��C���i���I,��`-�k*�����Q��L�n� ��>t/NRJ�"7�qRs"|���p��o.��/q�68����Zэ��[)�OhU�Q:�o�7��}��XbA���O��:��6��8���{����մP�|>���V�.�Rs�zx��?�%���~�L��,�0�E$��O��r_�ذϑ#�d@�-e���hwt���-J��̬���h:a���iw��ID^|����OM���\��-
:�3w��~��������Ũ+ۀ.��bszX�wj���ױBx�_/�H�2��U�)���AN0����s�.����_��s�WoM���ֻ��E.����xcwQݠ$Ŗp%�"����U;���Ì�M�2�n����H�#G�8r�{*W�Q��s0��zȍ:�9���[�⤣7@�_�� ��S�(s��6���\ˌS�}�(B�i5�qh��0"pQF0��?IG=c�[����7ǭ�.x�d@�&-,2kL�����D��f
���ǎ(V끅4Q	J�9���kM�)�j��Dq̬��u�I�lm�\��Z�͢K�3����ܘ�/Zբ��%�+/jĦ��*]��a
g�%��Z� 0d�'�A+��?zT���t�~`r�Y��aZᓆ#�Qjq��;��y���K�i���7���E�;Z*X���@6�T[g67㮽�7/�}��dhoAd��F�(4oh#�����V���C��
�J��� Сs,g/�!���8����;���cK�쮐���:5�6c��2Љӵ���(�@՗4���'�p	�����1C�r$�@�+�e�8�Y�
�/��uu#l ,~p�Mg�cz�j]�>����|.o7 �o$J�=<~U��19k�G�;I�mc����׆��x�xN�,��z�OW�Ύ�dJʀ81�Cy���l�.�s����)=����$Q��!͗�_~���t#x%�����NUS	]��pH��+b���a�,�w/�_��1M���S�Ho3]�9)��ޥ����I��%T�$���9�׏�>�����W{�}�)iǶX
��O�m$QI9�t�$+rB?�d:�IlI愱(_B� }��Rap��A�;� r��^�W�ͦ��R����@���0�>�&-�c�l�/�t���ت�]�P���s�iT��('�D��0�I��t	N�h�ۋ��W�í���7�R���$!�3I���c�8�ord���9�2�֡ờk����p��5Xʅ��"5�2���r��(��5[4%9,ЕR���6h�_���$��|��N�WEƆ���* W�n0��r�p�M|�"X�O}[ŗ�BY�=)������P���H�^`�c�S�-�{w3��;m���%4����� QV� NH���=�s�'��߼�ۗ��+
�5�$,�琇�_�F�w�3�N�x�*آmD@D�'�=R�I(�䆥���ܼ��9��Jq��J_�����N�gY��\�QC�JrE�:-��kie�c�w#�����ӄ��xnn��>�kE5�p���`7�7�KO͏�Ǵ��+��y���xHcҕ��I�a�W�i���/jp�s�Ht����FK�'������G{w�����K�X��\];n�*[�Ќ��V·��\