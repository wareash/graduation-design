��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�tڐ�!��Q�����xZ�H��V�� �]d��� ��h�hQ�/���o�~�կ>?�5�z�+|��"D�[�!#��.J �SJ�Ҕ�5�Y7�0�f[秡3ڕ4�O�~�	����u�Q�Q�H��)*��V�o���}m�'_z�8�y�@� K$E�R�5^R�Ԇk2�vv�#�80����I��JI,3)e�TN	�W�� M#d�*�������.m�Po��jR���R-�A�������#��Y���j��ȯ }�RUۋ��M��fS^���	@nYB��<�21B5c�EKw���2�(i��C���Ԛ4@AY9�a��i�Yp�Z��V��5u{��W����U1�*��Yom�n����{7)�&�^�fȘ�&c[�������1ɦ�\����;}}D�����[��LN?ű�F;Q�
����\�05rp~ @*5��Ʋ,��˱�b8�E	�����+=��z���V7�i=����l�x��}Հ~������O�ω1�B'�}�!����?h$L�󳁵�a�Ld�+5�rY�R|ߧdu��wh�1}, ��apH�!_�(�_�q51[?s�x+����3q�߶�vG�SCUz�)�6P��^����4�0��r�A4egH��$�pʎ$<�+4Mӹ�pC����8�c{����!ie��e���2�����P��:�����B�*��(�� /�eU�8@��o��,E��]�9A�Z�'í����&�I6n�z�H�ڿ�'�xy���C�F���bRy �Bz�r������H�V��m�'�c�U��A���uU|7��he�Z<�%����5�D��}� �W����HM(���\��b�j�`h�H����; �M2T9CU�~�4���a�b�&j$�����Ls��5�fAq�������hr�]��×2��	���
�4 ��ޟ�><B�H�Ϟ9����}Uc�<F�U�n�}v���z��4ی46����>K������3>aOitհ��x�л�q�[�i;�ƻ2��hL�Ɔs`��1��TnO�:SF�0�ߏQ����aY��۷�j��j��%�w+����uV�؇9
�"�)�K��5��_2)7uE[|e�1�B�kI�c���7�?!ļ�#I@9k�M(rW2��Ό؋��b�Mn���}�J��9�jX	��j�1�/'�\K�m�2�_?�a�Y#Ƞ���Fȡ`�&:P��̎j�n<��"��Y؝�CͿ�_?��h|�����Z���T�'V�����W�낈H�6�
�)�{u�i�!2^��%/���'�J �;��;���q�A��8T���D̗�Y�E�j�M�.�L4�-��M��Nr ��wudr8r�U���U����0WS`��|�>$�1B>:&g�{8<{�n��f`�7O�������xڙLw�����m�9�h6��*���.��	ā[c_�M��l.O.n��e�����e�2�x<tU�%ϗs�Q�H���H�n�o+_�:�t�wA���5[�}�
���>�o��P���K��5n�r�j}���u�p�_�w2��f��+җTXl���6p�"�4󈂉�4���~~�/����0���sE\��(c~mW0?��ԟX@{N�_��bhjNRWJ#��4NFc_!�|ͼ�,�gn���l4���^��Wb\҂�t����9�����H7#\-�T��r��|N'�*a������Id{SK���g(RswO��#�/�q��'*;�.E��a� Z!�9zT
s4s0,c��H;� �W�DV⌐�We����{�����}�N��[�v����c�}�U�gJ�U���g�}�>�K=C�X�R�Z�E�,e僦sd�ꡪ[�l0��9�]�\P6�һ��_4�d�֛�u�8څ4S�α/��W�`��L�g�e ni�%�6te�x@V!Zҵ�M�dG�9՜yl�U���:o0@��S�l��.3���
Y� x�E�z�0�/��I׊G<RC W���2�Y�{��Ȥ�ﻭ,/Ҙ�es.�;8i�$7�!q���I|S¡n�	f�Q	f���$���ތKVšsB4�:X�}<�|tw� [��hWf�N�H�r�AZ�cr�S�u6�<��?� HT?2���WkRQe~��*�G�SE#�?�f8ըB���i{�䲡����/��6�&#9��2�*�z�	�ؕ�MH��`�Hm�є���P�&I^�O+GLD���_�W��q.U�m0�}�5*6d&�����#ãW���u����J��l�v��b�rn�.jZ�:d�%_�<.��ag����nn?NX�'/>^��%��{��{e;�VȠ���*Vu7F�����u�����5��'�pX��k�5�հ͟��2����D���4����b�c�g`g���7n!�M���g��R�Y�R�t
1�J��6��Z������r��G@�'\t�hm/r��~��;~��Mp�אs�����c?��UHw�� d7a~*�$W8�p>��M�|S�%�!��4�����s*Z`q�^���`e��v`�*��ڕH JA��I��f���`�794�<�������S�e&��g.�M$n��|�{��"���g��5��]f��k��P��3d�� xO�P�m�c��M_O:�
&;{�8P-M�5