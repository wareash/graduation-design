��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�k�۸�m�i(b[�{�㇌�]�i�5'�`;Etg
<������"0F��}�h'��8��<���9���-�j����,W�_/�H: 2���x���CH�^�gߦ�Y�0��:ᓕ��Ѩ��`�uiRI����p�s% 9s���uY<�W?G�y�]L�"�8g���G��{�6=��'�$QD\��S�\j禗b��JŸ[�T�Dհ��B�/�b��T���M3��6�JlY���{�`���)s{1�0�Rnx���B3��P���z�B�&�$@�#�{���.��i�4����ǵB�*� MS���1�

�*V�a���ʦ�N�Nj7Q�Ҧ#���uB\yn�rl�T2HM��_����7�4(�H� ����j9��i��)��N!�9���t����U���.E�]k�?��M�q��r����ɾ)��Sn��i H��u��h9�c�3J� Żp�V����_Rj��%>���C�U�B|��,�J@����3�'��+V$@	��g�ђA���A�\�D��IE&)|�Q��i�v���R��稭�}��l��v>/LQM"�l��z	}_<�E��W<�
yTNk�8�P�<��HM��3��^���`�{~/(���2���a�F�WWP��gu*�w0>���kA^�uŪ�Lf�9BO1j]fW-���q7�5�+�|*7L�i#R�����9�oխU�yپ�Dj�_��x��6�Z���"t'_�S������f`��tq3g.M���G�rmm�H|�)kuˢ$Du˰#�X��X�Y��-�� ��ږ�~i���]�m=/���dN�CT";���tϹY��	l1W2a����J��	�[vIi.{y^���55�z������7֕U�,o�8�cH�|��q��-8iC�7��Yd�ֹ��4�씈���Dȉ��C��XFRGa�"tW~d��S|hRS݀�xr ���^RNǍz,�a�=���~3�GSg�ЮR�?�Ab����pn�i�|Cj)ub%��4�Y���ۖ�f�Z�ݍ�S��	�A%�}3;�/���K����W]��s8���G(-c�@��ys���d��?'Յ��N̊
簰@�����]B�}X#��\�2����LQ�i@�h\��� "�%O��K4��!餩Fb��5jYb!�?Th둄n�(�&!���Ĭ̝��-� �@�\���+� s�SS�B'4����۸ա����*�xq�����g���ċ>����&keF��Ĉx+�F��/��ljD�����R_�Fj;{ו�	�#L�{eٙ�0��������D�>�H��KiD�K�Jg�W��$<�ه�3QO���.�bαo���]����K�-�|�3���p6��s�ؑ&p�t�ׂ��Y)��K�wT�� ��� [�e;NU�WS	�Zȝ O�Z9��4Jɲ�z����\8���u�4�1|g.b�?.S�!�GP�7�K$N��r��c�g����\�n׮��o��M)K�?해��#W�eC�r���++ų�T!����XD�^h�L����7Fg1���'����q0�Hj�n-�8u�B�{�V^_h�� sV��tټ��FP�(d�"y�)t\8��F`������_d�Ԃ=�Fl�+vչ&V��MڅU"��4;�eW$�0�V�G��%:v��3����;&����A���v���<|eS�O�E�}�[IGNTG*�4�K�Y��\(����Z~�a���C��&v*L[��3�tщzv7�� w����]�nip�_�/R�[=a_%��.~o2�o}K��Gb�A��p�ڱK����H�#9f:��~#@�s����3p���`��E5�Tu�M��-�ӝJ���B:5�a��;�b�E�8�B�Ɋ��p�K8C��<U�H����U�Ge��l�[�Br�V�צn�� ��o����nO.�f�*����%=�2����j����&;��:���@���Ǌ�V.!x�i�KJQ����������|p����Tv/ ��hR��=9���J��˘٫��5ŭ�b[�"ZyJm����w�n���8�]�O��d�,�G���l��˹�yTJ�M��H��J	7	w���r�"���N
K�\"��
k:`5#]?�=�z��\>GJT�˫fP��ͭ�����U�L��D�S���9�-,��d�|*�)m�X e�uj�A�L�3ſ��Sъf�Cah�nA#��VV�Ѭ�2n��� G��p��Ça�};Ö�5�Ġ�M�KZ���
��Z��f��@:\�J7��?���m��g��%y'�A�f
��5���0ϼ��Yhn*F�d)D|`߸]�7J�Jb�<���N��	�v�r
Ϥ���mظ�B'ti6��R��ȣ�w�԰��!�.�kl�X�Z�x��<�Q��ّ3�e2���/�[��̪����%�B�!Q�� �/��b��]�/[!�]@�����ӂ�|o�)�kػ�̛%'��Jť
��A\3��Z'�J������t��c����fH8O���!�A��i-���V�W�֍ѧ�ͤ���%����k��>� ]� /͈�0.�f�f<�Yz8;���q���*���i(�w;r�ݜܠ��A>�F%!���}�.T��m���P�Se�L�l,�;nf;��"�Ɵ�)�:P��s��M�dR��/MVpe�=K�GR��☣yB��{�U=C6��8�Ս<`� kQY���]���M��?�mw�r�(�����&I�vN6w���!!�'���Y,~gN�Y��05"�`+�E��ο�Bp�C���p-�����a��v^�7�h.����B�|N[.`Avv�?���KW!����R�Ĝ��G��b,>�����'��b#�0�L
m����/�.�Z�������e�fy+��y���ۉ�Y7v���i�NV���,8Hdf�R��� �E���Z�s\��Q� �u׋]�HM`f�?�b������z���kɌ�{f�����,e�C?��n=]�i���̐Dk���[���[�a2y/L�*�]�ʜL�%����tA��G�'��kH[{Q��s{����v��)�M���gx�i��_��*M�`�؅^�bQ�}BU�P��k�}�B3���k4N靜��
R�_��{�"�'�S؆^p c�!v��מ8>_����eT�ߌ���J�)+�X>;��4m}�5�@��0��]]KɆ9"�R�Ϭ"�g� ��@>@�N�kNg
P����e>���^:{�I�M�F ^�kyii\&�i@#u�j�2\c���_?���d�&�P�dD�Y�����!pH��^�rF���@\㜆�V�	pC���1T�,f�7A��7b�{�ܬ@Q9R���"�3����;eB�(�d��v}'M��C���.?�_k��T7�d���q$a�+�$�yT�-�s�����'�
�F��tdDߖ-��.5�
��+寥�_����5�:�5�҃���z<׾K��x	蔏m]3i]�]nV�c���	�!�A
�ܑ�r�)ӥŋ/�ß� ����^���|�?���_���_������������Y�,�����$�A�7!ӊ'à��W�dx}�������U͊���X;���쨫�Lc���gM�г�
����ay�v�d�I�b|�c��m�}�>�7&Zr@Q�Q٦7��gK��$�x�c���$�k����7�:+��R
/� y�s絮��]ҖL�?�ZRyLA�HO2%܏aԃ ��2�4�"�Y�������n	�y��ݛ�afZF!/ò��˜7x���B��m����H�u���^U�NU�ï͛Iر��EF'�	�e��˂�<z�Y˸"���f�I��:xw>���R�ޡ���}cu��+��������Ue�$��N˪�2ȳ��k���w^����pT�M8l�q��G@�l�X�z�j�����5p���X�^�,�5��0���6�Y�5\#U�0=TH[����P%7�����re���X�#�#w�����9��C�
J&�9�*v���Կ�zI{a�P��ף�މmVب�o���G�}.�b)ֻU��.[ �sV�������E��}n}�l"����Ks� ��Qb�`L�h;D���'�����J�mLr[�p�������M[ ��n#$�ėT9V�G��AՠC�}�� [���踉��w�,�O5����F*�%��0�zK8눯x� >z�ow|o ��G���#Ŵ5���A��'�D՜�Q�.;E��ٙy�V9K{=�~Ҳ3gkTl�-��g�o`�34R�K����N�f����K��x�P�}+R����@��9'=V��3�?П�0nJ���F�Ȁa栳��<Q,�:Ml��9�׃�n
J�=,jp��p:��
N&�����"���ƐS�0t0}�* ��c�#�*Q�,Ń	؀>��jz{�[�D�zvQZ�)g���#�p͵t��jv�!W�0�����^����-nV��5T:s����&2���IH%� �c �5�;?���%ur�ϕ+�c Ηk��ߋ��12�J�69w���F�`+��Y_v�h�[��`,jރyH�
�Шe�R�Ou��2\�7@�ҩxۚe�����w�-y��5�%�7bbt)��1uٚ�$ n�$��V�BۿN�|���I\a���D��tFJ��Z!�
0	y�	ΰq��i�6
�mk+�R2��n���]�z^����1p�a�PX-��h>�U����4�(��=�r3� :o����G�`q�*���w��%n�J������[-��F��T��������&�s.�/Q��;�a��5$KBacP
"��\&T�B�>�d���aD������?s)�v}W��*���{Fi��m=�@�n�\ ��q����=́N� �oD=~������|�9P��ڴ�\���<.uLd�����>)!��љI�|�6LQk�v�aIέ��uX挔m��@f��QM��ҾI�if���o�p9��ߣj9�]���(�,ɥ�f�H�\�)ưp��ڷق���䢵��+n�;g�q��V����ǐg��s�O���Dn(N.?��9��Y)�ߛks�n�A�$i��k�4(��z��Z#,?oP)G�x@���I!��[��=ZV��g#��ro���/�F�2��Ee����w%��+�`�´T��	�3fX��=M#ihћ��
t�E<���b>"��V�]�O��y3#�����ƕ��t���y��{Ji)	��
SM�O��-m��>�N�|{�z%[�-�e�"���꥚m��u��S�� �ޡ���n�ABbQx�	B~��42���[��`FM��!08�{Ve
N���C��,����n �{�b �.�%�i�u�́YŤ����1�rl��dt�muPN_1$ڔ6�Z�@	��É�y( �!-sֹb��w��#0l�k+Ǔ��.OK�(;�lP�C���M�Z�;�Q�����q������3J0�ۯ�fŇ<�t�����C����6	�.~7�)�יc/�
�
���69p�h�GO�(�p��
�/������Q��4�̫5��}V�hg���S)����^���)T���=_{��V�%{�ح�iT�NA�u�%����i��e����4��~�K<�W��hDx�����x�H���DsA� _�^ɥ`�f/p��k�'�[5�����5+���tH�b�84��o�I��e�"z���x�*n�t؋�'B�"��Р�F��� ���Tm�prL��~��\����4jEfW��*��o�nd�h���S:�����ڋd����0cP�<.�(�}C�Pޏ�D�M�����f�W��D������� 4��1ݣu�#�M��씝���jHTb��kJ���P�Lߩ���]�5�������Ĭw���rEjN�Y�ܳ��:�>��w�u�s5'�<n-ԴΘH����qȾ�Ԃi�;$��z��ì{�J�3�K������.��%�D�{�ݡ��c��55n�0�ò����z��'k�B�9f�����L�����dG�_M��P��ݥF��mCI���X,�c�0��6��Mg��S��j���mDƾ^�bCdu�@��i�-C";�6
1��c�ˣ��d}����= &�d9_eZȽ�#.k߇rU��<�!ή�=YA#A7��!<a�0]�re��L���-��~��-ݰ���Q�5H'6����GBl�z���]eɿ�Ο��G�h����=氚�5h.���U2"*�F�LoT�!-�N�{.h��C�b���!-�{��IO�j��i;��Q/;P�P��G3b�u�נߌi-�,o�!6\lu�7Ex�v�U���M{�uO�jǈ�V��q^�c+m�I�X\�l큝v&���cj@䅽Ϗ�u�Ľm1�H?�@漢Ad�!ux�߭ȫ� ��sq����$Z9��j��x��r���T���=�4�z��WL�p�6τz0B]�ׁ�d�5����Y�Q��+��a���ϑv?m���b$���G��U�-� �lG��d�"N�t��ݝ�??	k,�DFPYfł[�-x��ǻpf�M��Q���P` o1,�s2�Elf�U� 6���[�����_���l|������|�`�/��QT�T��h/���	�{���H��
��P�L�Ɖ��o7$�[w��y�mk�_�{�7�͝ez��0���rՈ�Nb%?���q��!�����dv���ϑO�q�KI�Yx���E��@���L(j���:���2�MVܜd&�_���̨]������<%�5�����<9h�_2yI~[�
��M�#��2F��/��� ׫O�$	4P�����[��r��_��K<��y�I����;����J� ��{�یZ�ګop�J0���,�yF';T� ��o �g����0z/���&�P�������S��U[���aL;.�FT����(t�f�RN+�@ft:��R���;�#����YP|����ON��̲�9�!b���� � -���0~y9��e����h����5磀�y��ihˬ�0i�����L?�w��	�:H���qF�8�kb��msu�HF(�r����V�?7%���lN���]�W�2g�($D��Xٳw���'�K��n��?����)+�b��	���kw�|2ٻ��B!o�@���1�k�#J	�;�5����'_�y)U4㮴����d;�}�H,W�	�ڢ�z�U��QT���UA�(�ԸF>jUDĜsMbl
f���lQ��OҐ����O,ڴ�R�T�� p�כ��,�S�|��v�y��zP��2(
5X���rȫx��Ir��OĀ�u>`u�J�Ր��D�$Xx!���y3h!��ήeA8D�o�=e<�W1��/"��x!5X�!��ZC���u^L�H~�޳�`*T�^���II�:5�C�aT�{�g����P?����&{ʉ����ǯC��6����ޡ�w��j�(���.{s�÷C�;E��b����"����Y ������6������#�#���#|A�,H��j�eT�+44�� ��I�ة�fF�[Q; ���)�����a��ׄS\�*�f%�jBsL�:#�����q�z�>$�o>9�b�M!Υ��H�m�70(u�M�g)وE�\�C���v�*��b��ʐW'����A�������R@�<�K{����q#a�`�S+����[�A;����i���G��Շ��J� P�ȧ,.�[��2ޜ����ߣm|Ԉ`
�\%6.�YHǉ<BУʢ��_�
Ҽ�f2[�� �~B0=�J ����B4m[�N�^ �WVv�|���VR�� u��@��M��ȳMZ׉2�/Vl4���>���j�8+����	xcft"0�x��ݦz�DwJ��jM��U¦�M����Ѻ-El�� ƿ��^#^��� �Z�C�$����ٵ���$២�hA��qنz
�z��:��w�^L-�8J~e>��{�.<w�w`Z^1� ��͸�9=Wu&�ضX�Q���g��p��� �o�W����'R�Y�)�. ���L�����m>��Bϼ�d�� �q�(+�J�C��n�� JO7*�0��zbn���/�LAB	�)�(g���+�q�iN��;����w���li��������GۏL6�
���Z��Dbu��6�%�߯��~��
}a�7;�E��K��Ӗ���|+?|8ܲ(N�}������6t<�M��R�h��N�H���N�Ο��'���bYJEyF��Fvϯ-��N~լO������G�h^�B7ȼ500�T���R�*
�2N�����h�a:Eģr0r�Cۃ�(f8{�b�U��h��{�h7Y���T�K)U���Ԩ�$9ȜE��[@�8��T�AQLs� �.�:�K�K�yg��K�#��P�̗�;���46n��)?��PW��t�4�fk3ԈnC~����N��KI']>��XB�,(ގjr%�V���2$m�L�����Dq�v��.��2��ySso���m��Y��E(�DC'�!�z��S�.�6@�4������3�0�x���e�-;��-1Q��u��
Od��ɟaI.��1�PܻAX9,�HB*	���'�R��D@$K�//��m����3����9���ܸQ��1���,S����L�I�qf���V�u����r�M�n+�%yaվ�A�.u���i���g�,!g�=n����^J���Z��4vd6�BPY�xʘu��q�S�Y`n�W6%�lۼj25a���>/��i�:׼�QE�ʈ	��r��S2h�Yf��x��f�^+;'D�+��=VKFZZ�2U+ e!g��.t�0 ��F�k�?ѻ��2;�Ɩ��hh'D�цr�xg��Dw��S�ޫD��hވ�������
��M!�r�ug�+Y�&�=�Z4�n���춷�	�>����F����f��du��������Ѣ�0{�H1�
��* C2�N�Ԗ	B�a���f���NYX��*5ba<�M���b����xE����~�w�Tnq5ؚq:��������42���ԃ�Z�6�u� )n��<�4�h��5x�:�	3�3���Z����(� ,�
�S��`��'չ�v~sů��
��%���zqC��/��Ė�}�)�@a��Q��;��tśc9�U^�h�x�8��j�� i걒G\��47WP,�mXN�8@��)K�ޱ{v3g�&��㦅�F<z�l�@Yd�=�|��������:��*4�(f�F��=(*�t�
�'�����a��+�$�1P�ad�jw�~�����p�>��N���C���zF
q�\a�v�ٞ>IHD竽ZR�P��V�V��`*�&���Zͺ�L�ﶩڮV���N Ф!�e.�P�:�� ���,*ZX1"�ʤ g�uh�1k���<��b6���<bo��{n�I'�>cT��^�m��aGI�t�V䩸�*����k锹�S0��J��Y:FO��m��o6�^i�ŷ����|0�FӋi:�r�� �Nh'>�B)�x�!r�7��Ŗꗨ��R�OS#���1�j�ύDX�k��j}L�����NSG1���Ag#,��6	&�P�~l���|l�;�o�|�\�tu��;�V�C#$G1�:KbW(�� ��\0S�ơA����G�y�����+�G���yoe,u��{�����X���p��0�כ�އ+3u�^�:���ǲ�%����͊��m[�<���o�Ə����l��q���I�������O[���HIL�hS7��~9uv
]��avukm�9l�dM�o{l����)��c���d���B7-�h��f�'r�VZ|S#�>��ē~U�~DP���A���������|)ڈ��gC��D�m���%�����P!�+���
�2\�Kx����b9�5tCב-G+*��MIBT����[��S��S>nn�b(]f�T�&�B�{T���I�j��p�[s���Z�U��WMv,;H`%�p �	A��D���x  �@���՘w��:ܔ�S\Ʒ||֟�X�'�`�_���ۖWX�.���S'����jVT��uR֋��k%<����D`����Z�Vs�`#�װ-jX͚�r}%3�0�B�X�a�����WP�=VY��I���g�/?+�"M�#nt��A��a���h�����m�.�)��چ#�&٭w��G���#��L��-+x19��+�a��qYw�s���~&��
�pi�k�����F}��Д9�}	�*�4�	"z%R�#�W����`�i�9��ȩ�- ,TD���IC"o�� ��Y�͆��og m�n6�-2���dt�Y�󚃷�`ؙV\���3D}Q�1)������q9k<�p�����Sٜ0B��!���1S�1��.y~��թ�i�@�&Tz��@�.����A)a�W��1������i�ݼ��:�H&�]�® �4a`�K��"�;`++\�+��H����(S����)�u[�CbH���d��T�%��:%"����$���l���	�XIbc?j�Ⲃѣ�Ǯ?q"_��}�!�x�k��V,�{�#N��Q��L&��9�lǼ�.ѻy�E���J�*� �9M�<оV}�IxxA��*�S$�^��ll8�	��HD�
���إr�����F8vJ�q��ig72rL~_=�\�?ܪv���eG'��5tW�l�p�;������Cm�m��l#�3�q�ڳn�n�͝îa��D�d��r���7eҸ��v���[��B��9gry/֓�?R9�ɣ]'{(�MR�����sZ+����En�����jQH������<�U6�Ή���D��B�J��cK�w�.�V���JpU��	�"3� ���N�b�՞pt+�Պ<�,�C����!�*`�gL_S�����C|�Ƹ�	�2xѼ~�8�2��K3���\�_��8�8C�6��Y�^C7<G���f�5ʡ B�P�P��V�џM������G�����'�$�D���70Gߣ"�N���������Ld�|��I��a1�6���?��'f �Cv� 7ۑ �N7��e�'t� �\�H[V�{� o?|,ܖ�[���kh�[�|���*?A���Ό���|���>3j:�M�����<�iG,q=�l�/����*ȗ}1Q��eÒ�*���_0��mfw����%��DFK�V=٪T@t