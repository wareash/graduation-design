��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf�&���>�m��`K��+p[�������7��5���1R�'6�2')� o�#8�*5Q�����Fi
�� [NQ�c�T��0�U)#$�4������I�����>��0�5��2C�7�_xf&��So��|�9�1��"�y}JD�[�S�3|�r#��U��U��j��$Obx<#T�$\�5%�����<Lz��l�M��#�Zt�R��Pw��1ã��x�|.�G���f�{��j|ezZ�W�������4S:���n<m`���W�)��C��������d  Ei<@�'E;0��|�0V���Nf�)�`��w�J���Z�Q`��T�)$��=������ЕWp}��75cA�E�D������`�d���* ǁ|��@tЫ�9�W��{?��
	�Vi^�6��C����YWMf�IR�{&�vW��ť�~B#���c_@���`��-���nm�M�	�BƏ�6~��--ҭU��x���s���]��d�gr��}w	���N�8��-FȬY��e��H�w{L�NB�9�}be�ـ���r�P��J�Z?�E�U��PPVX7R�K�D�i��|�q]�Ҷ�HE}ܟݒ#��@�ܹ>G?LU~�.����hy��w|�u����s�M�Z�&�֤WU���id_<�a	��X��uf)pU�y>ZXO�mH�aM�U:��8V�e��B=��>I)i���|{,��(ȣ��~��R��.��`EHj�y(�mF�D�Ա���,�"�J��<-��߷L��\�����8����>W&J,�/�w������X&'H�FQs�-�0-C�����^��7�����\n��(�9��x��
����97H쏠l��>�d�
.S��ݭ�uW�o�CN���^�JK3�� ����Y��h�p� .�K��yU���\�0�`�t�?n2%A'趉�0<o7�5
�n)�l�����0jv������f~�7�_�=UF\�l�P)ar�(�&j�0�t\�\>�Q��`m���+�N���d�� B'��ә�'}��\{y�E� �H��Q%��'�WV���zQ�ՒƂ�f3���.�($쮏6�Č�˒k5p�UԥQ� �)���O�<�4�{����:|~o��o�\�z؈"`ؽ䆾��u0��ݗ�ǆ�snl���l �u�7Ճ�膦l 	6��L�}=����X]���W�&�\_��d�ef㵜�1jd�)�f��c8�FU��J�zgw��3Oz�]����^c�~��r���,t]��ᝎ��cΐSċ��
(MV@�䘷���`�*)������$p�"eb��=��C
܏[��wg9)pւBWUa&�ۓC���~T�RqJ��s�[T�N+���^ddwL���J]�ˁ���D��#7�	�k�a�G�A_W����ogA!�r%Pӱ�h�Y��:߬2I�]m���~[��x�jO*2\����w��fO��{9��N�tt��?y��3'�`���`�PP}*����t�����Gg��{�ދ��?�#n.o,(zn�nsU�z2,&ѥl�L���.�f��Tw!8Z#~���<sz>�O�ܸS�sKf ף�c��D��~�qjh-�I��N�kx	���h�06�5V��'5�
Yv�z�c���bA��&��396ɏ=��Ɔ�x�����v�=�\y�!�`o>���oT�����"�<3��m%F8�!@�`���sI�7V4ߚ
4Ձ�[<E���N�U��}>R���G��d-*!>�`�����C����q>h~��_ԖAYzᯩ1sЄ�I��ze$\Q7y�l-(if��TS�؎���#�u�� !��h�ɉ���%C]q���^�_�����z���)vÑ�P�Vx��b�SZ�L�n!/m�Ͽ<|�,|c���S�7�i26�Ւ�N���̻��1<��
��i|ȹ s{(���Sg�G�f\[��A32�|�f��D���T��G����}j�����73.7$��aP�� �((@�W�T�\����s3�'X<ۼP���Ԧ�4 �3R�:~�X��H|:�BƤ�@��hSIj9f]50�}$��Oq1M64kF��Ey;K���
c4t�@��_�e�錛�]pd㹜�˴[Wa�� ��X��؏2���`bQ�!I<	��S��pa�c��RC���D�O}��O��£�_��t<qRo�N�P�F#����c���n�ʕw�'>�g��ߩ�$�VJ��՛j���B8��#��}��F갻� C��k��N%��d=�[�ĩ�}&�DJ����Q��МB��4�=���̧�ô׻�AӀ&��s=/L�1`$�:�~��R���^�;:�´-�����ΛMp����_��n��_��y�
C��Y	��=��5�N��._�q �'l����5'�(+�.�8��pv]����Uz�DZe�i)
�;��Ȋ-��G�@�Τ��s����B���t����;}�����/m�s��7[?��@}r���P�,8�t�8{�T�_�U	prl���B#���qbe�i��Hse�ف��0���&�"bⓞ�^EI1q�Y�d^`�ĕ�N!Wx�;��䯰����c�G��f�q��ETj)��@OJ��s��&�O�מ�Y���"��f��q��v��Ri��>�[�"r�R����i;*�c5���x��h8/�;g=�N늮9qڗ茐��VVz�L����t���ye{�����0=\��/�5�V�����4"m�ύ�S�Q���*��GFҩWNa����܌�=l$�j��F�C_Q{��n���O�Lٍ7J�Θc�n�N���e�ԂJ@��jvx�`�k�8R<P<��1Y9���ֶk�ʒ\N���.Ա�f���W<,���[�O1��,�%��(g��Ļ��M�*�uy\�C�V��l����ek�P��t)�Kk�z-"P?k��i��l��α�� k�_?Ä�k�(��r���7��)5f��$�I��y�ɋ�_)W�o����c��lo%�4fp{΁�䫲۴�x�4G%� hF�aA�7^�2��>�Q,Կ���W4	��n�i�汣����<8c�Y�L
{Бysa�1&���4�Wr���jV���Њ�bvq�]���/��X	\i�8��9jU\)r�x=5�����%���r�*#a��*���~ߊ]��&��.��)p��p�T��gQ��x�X���!DO)ƏE%�{E��U�e@�/�R�EH:�%��@��)��$�����""�:yT�[y7�=%r�;��;� �8#~���g�rp�oGm#N�en�7���4m��8�O�{���.ij����d/j��K����㿫C��{��uM��>a��ʇ���ǉ�4s4zc�+��0B"�_�A�%K���u*�3