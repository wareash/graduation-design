��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e����d���f{��@����S��>���4{��ת�AO�Q{���~�}Q_�=��3��y��դS�.��P�	�ᎡÍ7���&�5���uO�F�	�����@n��MA"���_�Ѡ�a���y�Ieo�>f����HL�y�m8/� �4���a\Bv�U]MnUf���2t$���u�IH��OAE�)�T�z("���m0�k�|nm�5;K&�����O�A��Vݖ�\j�W��k�����而7��^f�5�`�=N�0*\���*�Ȏ4T�lBHFh���_�h���<Y2-��G���mb1��(OP�_�1`�de�40ɇAW[�N�FHу���7;��YS�y&��Q��33���Nfy��Vo>��.h����"�`�g�#r�N��?��G�[{���9m{El֟ݳ}�9��&Ѥ��c'���R>=���g-T_��n��y �&�Ue�*2�SkL�|;ό�$��L��*&U!��?.�ן�������^�o��B�ޯF4�"|��^V56&#�׬O��@�捞�e7p�W�~�tw��),0���w�Ḽ��hbY���+�Q�E�O �����z���$��%g�Zk�3Y�$�#с~�ET��V����7���	<���@�ny�w��+X�M5�r��b`i?GҘU�)��h\���������_?C�S�к�7^��"�.l�29E
M��G�k�A�x�K��������^j���>��>ܚ(��-9n����/[�x� M��U��B9y���f ��h����c�}��eԇ8�1��y�=_�z��A�rw�q��������S��ޣ��#��`n� vG�S�(y?F��ݛ�OK�Ї��DJ�Z�e?M�Y�����=�p~����,��������j�RV�2rZu���u3tQ��������7�{x!���?�f�D��ɔ�T^�=%�ʢw��F�l����詞-`�ՠ����M/����fE����:%�h4�I�߮Z����%q���m�� ����aޔhUrEv1[�fї_��$��/�l� cj���\�2?�tK�i�	Ix�d�8�Kd�(W�3A�Db�Fü�f��Qk�*��e�����4D�]T(�,$-�J@̈́����>����ǪQ�K�.{ ��Wq�ܦ��9�����n<e���j��_?�sdi/��)��ai��Ls�����z��%�1�鴞�z��{��V�x��+dF��8�:Lg*�Wi��]�J̀�{q8���sk��������
 ��[�!y��Q�}�<D��ːޫ�4��>s����)@Z7��-�G1]�Uڿ[{�����_���)/�{��?oqdFE�v�VD�n�Я����z�y��s���˿�ړ���n;CxJ36�R[��9�aGI~&��qP�|�@>�0����iP� 愰?S�$��w�l�'�y���i�my���Lޤ�u���5�y��sd��A���x���\X�\��2�UNQ ��2h�s�U�&^?y�᭽�� .�D<�'~���c�z����;�k���"6I�:�t��a�[�7��_������_D'
�����HU�I�?��4Qe�,X]l7�o�޲��:�{�]?��7,�}Bu���Fb��P��mt���ͅ��U�7^��@�\El�}��2�0��ף�'n�V7�l:����CϦi��k�61b��b�C�k��܅l�A�_�w1�q_`�/%4	������y}ee����;P��~�"�4�t�w�8̋<��B�**�a{����m��?,�o�^YP
I��TF�F��0�\#��b�w�Aq,T$	�_=C�E62��6�yg�5.�ȴr����pO�X������Dx)M<Yþp�r��l"9�v4�$MVx���2��%�P�t�<̣��4cѲ�3E���%˂������:*��#�[���S��"����ǅ �3qH�t��ٕ�B�Ca�u��2�/�2i5����q�uyi����d,/����EP?�YAl�"�کK�=���h�-::��fb� 6�4�B!J<Q���녷��feZClЀo���V�DΜ}����)�^Y�x�3D�)E�*Hu��2��}�&k.��s&� �ͧ�
,<�"QN�7�Z�h�q�	�p���U�檗r=�jS(�o�X�e��W��s��H]R��?����`�4U�SB�q��9�:>��U7�S����kc��KX�_D�	�6퇖#LR����4Z��e&d��  ����ܥ�x�`-���8A�]����- 2
2��dw*�OS�ޥ�u9�i����_C=�K�U�&��dB^��ȟ>h.�l�,���}��Fa�"OAQ�H�cr��fO���hɶ`�a�#5�}���V�B3�:4�Xq�$���C4�`*1�t�C\.1��H�/�@\���ћ��B��|�ؠ��FQ�L��K����7ؼaV�y>�;�-Pi��N)�f㙖D�6��l��7a�VC��2h.���	N��G��?���M�E�>s���EF���P�n��E�����m��5S�� X�Ԟ졼	���\=�i�z����6�f�{�g�(3����:���Sn��X�2����ҡ��1���|��'h�$��ZH@)k?���� �ӆ�6N��j��_��A��Y38���E�0؁�y� ��V7�m�FS�π�6H�>wU�r�	�7�V�:Daq9K�('[��백Z��S��WR�YN� �_σ0�Ȩ0���5�%gP���|��6���s����+�[�b�i�u�|�gA�ѦJ���%�56Q&�g��҄Z�g��W@ꨮ:��,�`�F�9T���!�W�nhq�B����B�g�჻���}���;N1\T���Va
W�A��g�Z�b���7F잲�&��h�~�%4S ��C(2v���6ՎsB��!��xf��Snm�Iio�Y}l��|(|��j�\/Nf	�>	J��s�Q��xWv�Nf���7�l�L��v�:Ϙ�Y�ۋ|�Z;�{x5Z��}�� F���R�&��NS"`g�]}[�J�p.~!U��l��=��`��&I�jLfk�0�	H�3�W�����G��k�s ?��?�ϜgaăCv�G
�]Xa^[��Ai�	��k���l��T�a$\����/ޓ��\]��;9�V��l���ʪ�-2wx�M���xr�ØA��x/G�F��%��^�V��'��=�ռ!/��p�=��0+�!�D��*u\��p���;��� NKq\pL�ϫF�"+R� %E/�G0Ue�b��@�l⺻���ڂ�\p�$�K�j��'+�f	�ܖX����A0(���۹#��Ƈ�%^��3%�G:�O[�4���#�VR^��˒p��k�M��beϩ�F~�~����.<m�����
��5`m�x�p.����+�'"�_ʧ�t��x���~�9d�d���Vj�C���_���\����]�N;����f2[S�z���^h	�bee��:V�^�G��G�'���k���oG��~�������a&��T)_{�AGF;�Ww�� �97�X�B�`�a2�"{�����B��9Fl�^Ah������b�����ӷM�ʗ����#�E$T�a~ �_���I��?o�V�uF�D"����D�GD���U���a����X���"�&jR��̍w7���O�}��{���*�$X�A�IN�=�8px�%��|u!,�1nN7��.C��8;����!WF���(_�r[���SX��Ɇ
Z�̙���	�(��"P�ˣA�T�s��C��w�v�|}�;Ӡi�hv0���7��<3f|�CX�ra�7^"��&	���p�L����o�YȗQ��A���[S[���̼�s-^�h�'��n2�	H��?���L1��e��+�
����ܻY���Ģ�"QB�o�|����I|��f�n6E��^#�p�zv�f��`J�j�������`���I�Z�b�5/����"ԛ�ɌR����m�!]��o��e�+,��ĸ!�C�L��NA펥���;?�)����+����H%���Z�D& i�ؼ?�{+��ܹ��{����PP��9Ғ&w�@OW�Jb�Ԧ�{@�@Gaoz����:(�5���N��/k)x���<���p��8��OZ<�ȼvlB��&\@���6��C�m^�N��Ng�M;?�X�V�4�5�ٔ��L���7�l����q�`n�T	��� z��v�靄�;�O�Ԉ��H w���Mv=�Y��^�?f֘�d���ɉ�L��ܨ��%ۛ���8.�&o�f�^cӹD/. ts����G=ן�%F;�ڐ��#���++���I�Ȥ�ȅ�'���81Bm1�z�,�T��Vս[�����:р5jn�ݠ\�8�S���zsF�����n��EY(>T��๢��z=)<G��}Ke�� �h��ZBn_^����x|e��2N�.���>7Nw����V��0�n�Wճ��{����d����	'n��Sz4����d#D��]Y5��������l��� ��$�k�����!!�o*���P�fƛ���k�[�z�P�*�Un���%N����CȂK$h��aji�Z���`������1S��+l�,S�-��[���ަPim�q�T��G�I��ܸO��I'��]���7IL�z�5���f:[�_���K�,��}����5р�M�|����`u(Sl��`�-�;&Ǎ�������1Tis�A�g��eM&�*m�{	;U��H�~iH	w �^������3N�_|�Y�E
��Ҿ}_�B��`)U��r�9|L���q�F���B�ZPaU����=jP�`I�����g{/����++�qG�*I̢�����|����&T�v6��8�H��z#.M!�����9au���iP&�{������A6I�2v��NR��&J�m�M��b�{���'�P�YX��b�L�!�N7K��e����RL.������d����9�*H�1ѕ�#:�o�0�k�Z����av����R�O�}ړu��׽_�jWl�%��`����a2�YQSb����@�#`=Us�eB�՟y8�2�D�t��������,���a�A�%u@�Ǣ�^�fQ��rQ.�҃j�rJ��7V,Ə����~���h{��G�%^^��ꀗ�4�tA��?x�����"�V%-�b���	s<L_��Y���_km
Xp�ߑݮ����J�x2��~���;Y��Fi	���w
�Q�<�4�3B+�Ҋ&lQ�`䙜1PqV(7�͞�e�w���B77��{��b��YД.U���cO�͵���?�2��5O���,��X�x4wU]��hMǨ]�ot"2�CB �jrE��CB26�]L(��&�qv`*(e�w5�΂ФKT�{��p	��w!��N�=�%�J��ěAw��y���71{[�8��%�)B.W��o�*��W���?0"
�����Ⱦ�l�q����Sڼ�c��^�F�a�������6���o�u/v����ub�Z�sl^���# ���V)p�i��[�5;�����o��0ʎ��[�T�.ٱR D�6�iȯ���c��,�GR	�it�a:M�x�Aȉ��R!+�>j�i�����Ω7/�jm��<����(�pW�n�R5�,�2\������߰�P��h��z�g�D�0���,|�=�Z��o�R��æ]3�����ff$t6��vN��`�>��jN%Vi��;�߱Y;V	�"�E����B�1����@�3�wszk|,��߽�:����%�O��Ž�ݑBӅ���������8�d�`	�.���p�N�3�<��MDH��	Y0aKax݀��Y�W�z��A�ۮ R��v1!�X�����0�V�r"K�iL���>�.l�ٓ$���V'��j<�h��٣A�C�lB�t�	/Z�&���)oղ�F-x�.;4�U�h}�^Y1D�����m_b���$q��v���\8g�w��Q�l������%!��r��������\�m�T���e��!o��;��/���d��:�h��r^W�>Zڮ3�B��L���8}��6�pd3`ʃJ0Wj:U�d۪	�����	??�����u�b�iӤ@>�Y�?8{ɢr0��ޟ��Is�'²�&�=�0�:#�.��s���-J���D�[���tUv���MhDX��dG�.��
~��5T��d�i�!݋O���Y>�����N����k:¬�����u'm��̼�Q����ʑ��"���N�mx�/��f�1PM���;7v_Č@�p�� MT��H����=ȥ,
�ˣ���GY�%�!���^�1�QG��qJ}.�AZ���Y6�?|쨑�;l�:F��Jo�2u�Z�]ӱ�^grI�]o�>�ǂ��l� �6i=�b�m�9`u�������g�g��N|�"�B���zx)[���5{?w#?"ֶZ\@��V���7��
�m�Z2�-��vY{Zcb�Ѡ<밌�&��i4���� Eԉ��0 A��>C	�����bY������2��]�VNv���!��c��3��g�脿C���)v����|�P\�\<y�Ojǘ�������#�s����Dު����g0�Ƕd�':��9&X�cO�8�1��+�vg�ueDI��u��'*�B�L��"���؈ҿ#�.`��O��Aq���qOs�OxҬ��Y���:#"����+d8���m���F:�o�~� K�v��W9xSA�l��i���ds��r�� �^4��7Jin��R�^P1@`�m�!6]���bkG�md�p:���ɬo'}�pR��]_��ja�{�K ��H����?��r�?5�n��5����j��DڂM?h���N�e��T�B"��@�5�5%��k�J���lp��/�����q�sڼ+�����N;x��Ԣ�TC+�=����k��\���e��������
�	yv ug�0�4a��-��H�8�����я�0�Z����˘�Q�I�f��C}�<�̀��]�Gw�?ͯ�	Y���(�9Cd�m>��~f��G������ܻx	�mU�WfZ���C���ʌŏ(XR;��]�ܬ�%��:L�}�Pf�X�"E����)G�P��)F|�+=Ec�8@�3���K%X` f:��<��T�:I�v�#Gg��x�+�P�&P�_�x �*�|�C�Z;S��y��qsĂ������7�]���� �&����޷�=��>Y�bW|�湴�һ�Q­�)f���HH�ީaG"9��;S��
O\��$�kmP��ZRSߠQ�L���ˆ��yTn��W\�&b���+��r�������t�Ɵ�-h����{������2���	��	����2�'y-4D1�o�Wwv9�x������g����1A���;X ��~N�{	�V%������)Ƣd`��ig���\��4v�^%l�w�-9l��eл��nAk�`��u��-���*�`�����?[�vf��
���Q�TzDf���TEѣ���{��|���dt�:��L�C<����^�2j��F9T0�u!��v4�	�b���|�����w�5����&�.�!��GQ��*��p�����v\l0��u�XDY-��<����&L(��-�)�@�x̮���&�&����V��',H�숬��_�<#>�J)h4��%������Ž�,&�Ş��|Ϫyz�}�����Op�q�k�� ȍ'�7U��(_�����
Z��]�0>��_��sEҷ��4W��Q��2�74�>d���U?�_v	-�=;�uږ.,!�D��/��[�@��`��<������yb��M��� �!�t�0R(��:W��\�f(6��"r<΁�����7��mF�����ϫϑ�UV��2�U�S����@�՞ ]eۊa��x7�.����Ǣ�v��6��_Ĭ8>�Bx�<G��`J�vd:��wn�\����mp��yE��M���z���[��4y�j�����t������
K"\s�J�����g��Tn\��e#��fM&+%8$��2�8]܅a.�0���v�6l����uEK[�J�ĻO����
���k�z��qhc�M�u��&3^��OVe�Dqs�E4��������� �s��z�R��6V��� �ɌT��i4P9��┮���h�,s�E$�|�Sy�n����3�ea�;���D��O�ʸ<9o��������c���*#�h;�oͪ�2�Qbf��w����C�Ң���X"�\d[U��T��EK^5�i��5��\@6��I^�|� �2𭝡�T�(��u<1$�Ԟ�d�+��:���yX�<�h��U��rw��ۿߔ5H��ъ,q	���8���t��ʏ���l7�	v5<[Qkˍ5�D��䙉?����	���V�ڿߝ�oK��Y�6W�9� ��w���F��C���1��7�}ad4f�8�����*�����x��
"�9e��8�0�w,��9fi��eo�H�!���V���`��(Ln�6�>��-�)v�۫�G��;X>���Dy�t����4���'�
/oۥsa�����/�	�i.VY�nUU��	�_7&�&:��� �k�M�O4���yѶ�<[.��ega���fɓAZ<�n��1�3<K�K
�,�ka=�hw\x8'���F5Ӑc��	܈U&�m���:�����6j!���q)��sj_I���<���SZ�$Q@{�ڨ�Ff,�?Ö�8N��+*h��H�1�`67<�Vj���"|� ����|SOģ��x��\�nP�{������q7�I�l^���4�a�j�am�٢�����J��d�#n���*+��jp�{��	�ҟjL�JU����R�ɉ
���"&eh����է��ػӀg��,�g%�p׆������a6?m�$>�:m��v,���~�#�rN�"���1|@"��!
*�}=#���F����bP�2�����z�TP\SY-"�*���������c|��5�Xo��8��F'��Z0�q[�.�`�Ѹ�����7D����*<��69Sl�x�LMQ�4�ٶU�K�t���_��ү�ae^�� ���[z�+]�ob\�#s�Мp��?2��*�U�,�:i��(�������<��T�~m��$�i�n��ɏ�f
a���Rf<�}_
P�I@I�/�tE�ĺύ�a&y�U�?hf"#��������B[�QdR��d��ُ7N}���w����o�
JpU��@N��#*�t�0@�VQ�M������&�=�.��r�`����GPJ���p�e�N#d���5�ڨ���nu�0Ӑޞ�Ȓ|Đ�o�m�PjA@og�ɂ�3�dp^;��b�S��W;t�Q7Ć"�U��������r|_=Ciݤ�"c�*���Ϳ�2�ub`R�a�\��[�$�|�](+��%���+��u�:.��&�pR]�cg�w�{�g�:�(oN$#a��7�4��B���CQ=痱	�xd� �n��ǁS��lXe�&��q�7\�I_^��O���_�jz�_Ŕ���tl1Z^-����yz �@��`l�#����'��O�9�mJ>��f���M�X�2ܭ��j�	!>�$�m[�m������U���=+E����s�a�j��a4�B��?eۗ�U�/f���N��� ���l �~�4=���J�MOu��T��bK�[u��GC,��L��=�'{�;�"<$W|G���U<����K���p���Y���_�$Nk�EF���q1�f�pF�����B`�#e���D�<�,g����S̓u�Q�9LN
�d�JH
פo��B�rd�����g+!���6R~� �1֠�4$,��� ��.���n}hD�,I��ﱸ�3�
֝��c�GJ��E�pz���+i���	�@� W%S�B��-���Q�H)�Kc}d��
��L���r�Z�|�gc��sޤX�ػNT���w��J���u��a�+`Y;z���{D����ޖa /V����M^l���R�2�-e�W���>E���*�"*f+��CC*M�^�m�7�R8x�?ɛ����T�>��3N���CS�uU-w�a5�T��_�7}@�ό�~�aC�D���\XSNrv�Xj� ��;匇ٙm�S�~�g��˭�Н�+�@6~�U&~�|�f�I[��e_E������ͱ]��1�����j1���c��ߖ�0��>��d�x���||aeF^ӗ�IXX<A��g^��s�
�ւ,���̄��3��L�?��#ߡ��:�bՅ��;��L_8���u-['�㴵�R>��b���\��o��5�ԥ�~�y�y�*�ZJYnQ[�WZ��w�O'S�����������"���	���;DOM�d@�F���똊��T_���A,�&�u��6��"݈$�8���ku��NL�r�� ����'^t����d���
���#���& ���N��%IO����Qo��&\��_&#�\�Ϣ�KV�y[�~�������l�<�K�hK��/�H�UV������o�Pp $ݠ]�d?Q�'����s����
��S�� 8\iH�IH=����a���d.RnHc6E�{権��3���T�;�C3�9C輈���1����M��"n����˛��%�?�\�H����D)���Y�C��	I˿p��Ձ%XP#a{��j��d��������`�,}�D�<aosP����%V��r {���)�t8S��O��U!�����h�� =������^	�3�9�%���'�x�"��I(���iL)k@Z�y�X���ړ�zM�$;ٸ���a����;sL�#9���2i?�F._k>�Dk��%���R2��Ku�׎o	������Q���]����&l�����Z�r�G�z�Gͅ��������O�������;�!Р��ar���P�4P�ij���!�jP-�M��]�\�ۜ=�nDVQ���(Q� �]EEo��5� Ҟd�1��E��3�qZ Q�#����aw˵���%0��Չ>se9�h�A��wƹ&\y�K�ɲ��D�C@�;��ӊ����͈U���"��'/V�=��C�YBsw"G+��eG�ذ����!޲��O��#x�ub����&Ej�����K�
��{���	�,���y7������bb��"�.�ֱZq�w}����F��#�ئ�e�;�W�[d#ȶU��l5#*M�����y�%���]�V<�̷n��!f����������,oh�mwVz;���\Bi�_��[
�e��M}��)0�;�|��[��8?�6��G@Bp��U���^��_�)/�)����	������r��0	��s�n%0������DW�k�Cm:w�OEc��}�GB���<��6MeŒg��G"}�W��Q���l���)ː�G9@�1&�5��a<e¡�Qn�ɔ
L�zc��hI��P�={#��l���5��]b�<�L�#�_"�v�0��IsZ�ЪԇG#"���wWZ�v���7��i�Vm����6ޱ/!�~� !8��'���A�6�7���j�������_b;�M��a��Ob�X/�u:���3ڕ<��{�r@��9���Jܚ����%c}��c7��k�C�Gc�]c[g���ν�4Q�Bߛ�\5�E���'��:��+�l��/Gug]9��]�NS���~�yw�N��>�������d�V3����N�ln�1p9q0�F<�b)�ӻZl��t���X��2����&HwW$��̦���_F���VU:%*����xj�l�f���OX�he횋���<��'�iq���$﮶���1�63i�����G{�lj?��[��[5����m[')0(Ӻ;��-y|g���הp�֑qM�C:����/wjbk���β	���!F�ka�s{J�1��߿SC�Z�� 
�zr�znK��r��`T+�)�?rt�w��(-A�3�O�� �(��� �w"'��byd��8��a~��x�Ē2�i΂[�.�u-�:�Kc�}��"1�G�9��6����Z�S�]>��CI���d�pr�"�n�� ic~�t����k�^�U�8*՟�+QDВJ[��g-Nn�b��^(C��w��'M�))�\(xy|'p���2���+adj��6^�D��gq1`e�xls�d<���HF5��̀���A����rXR!l[~>��I�� ?ѭ�,قl*\m=���É�����x�e�D�;1;�i-@c��iq�1�*��'!��7h�NGuf�Uٷ<�$��K2��%75z���t �@������R���֪���`_��7g_�W��x[g�i��Xx�O��ڸ��sӏ\f�mj�!�F�I�0�*e�(m�t�Z��_1yVW�(YWږ�]�d�bO�1�݃�HG]Ɓ��RrG�߯cPz5~� ��#��G�J�Q��.kC��ϡ�\�s/�d��e�?�7�w��r�Q��Q:��72ޤџD���L�9�n�b��|�d�3���j�N(ng�nJ��Ni�%L�+��WQ�U[ur��ڌ�<�$�x�'��"+����r'8O�!Wh����	��)��8U�����)�
E�k��8	Y�l�Q]Ӂ%�{WG�A�tiU����5�MX���V\ ���ɚ�*��#W�:s��Rmי�/�P�s��n��r%b��@w�� /�n�ڌ{�iɱ�����-�Il�PZ��ˆ�4�i�ur�ɷ��bZ�.<�W�r#��6$�8����$\vzd�>�a��_���n��qŘ.�xFS�'|[槗	Y��CiICY�b�_t~@p��PET>��ne�祄~Z�&�4��_K���c�L��1����d���i���������婉�h���+�LG��"���-T��=P{Z%��h2���P�
)�͉ ���P��᧧�X#��|?�X�:uōM�5�.�#<�4X�5��zW(�1��hEIXa���,��#�FS,�I�\`vyɤ��BH�������{\��y��0LU��9PR7�-r��eo�&h7y2kP�&$�����t}o�r6e[�*ID�=3Ye� ��+��Y��P!ַ�7��M����gm�Z~r��bGqem������T�a��\W���z�e?c�� �W~7�z��b�)�S������I�	�u놅���/����4|(�\�m��9Q�I��e5'~�ɀB:�n?'�n\^D��@���8�T&*���z��,�tɰ\�d.{�Y�<���agc�o+�']v��Eh#���[�#A��d��I����opnW�8}Md�ʼ�W
�G&�܋@��6��F��~�iAmBāi8���Y��c�1������/!e^K�Aaݷ�y׈o�P�=4�r�;�
_��w;5]{�r�����#:�<��w75������g߳♡1��6T�t�f{�WS���1�*���v�X�Y(r�"�2Q���W����DQ���)44���E��Q��F��bAEاn�;�8ͩ:�V<Q.�<�1:%���ԣS�aǄs��p��2�<cC�I�qWfl�%v#MVg���٠z~TVC ����_�)=�v���W���@�4������7�$���5����x��w��,2*�l�`��[^@�M�	�&�PksS��^�-��vP�y���"�$�Z���]4	V[����C��S[��pȚ�gI�t�R���[������]��/=MT�Y��s�/3g�ʘ2�/���}7#�����Y/U#N�Gr���S�^(x��B[�襜:��&�>\v[Ҕ_��E�����d����L� ��ܮf����7����߶��O�~�e�W1�_﹁[�I�c��7�1·{�"6�8�<ˡ&�y�F���-|ද�]�*P��Q�h�0D'M�ڪ�~NM������ʙ�2�6��������6�-7bs�F	8,�,^|Oq%%c�~�FO���
ҫk#�����6�婾����z7�O�+�$=�6o	A߫��������X�V��f��>���%���H�ς^�ú��{�P5&�)�S���oU�2�b	��Ӫ��;���X�ьG��i����Q��V��W�q��G��t��Ľw�?����h���͋r�+d��	��<��qۊ�)1�(�*$N]@Ϧ*���M�8�C��-hf�a�$@����Υw/���Ԙ�N9�r�F���J֪�f���iQS*J�{��&��>՜�,*ڤ"��k�� ��g&7���ď��0_��%"0�۔��w�)�0D�,L�'��_}n@�g<���~[����r�ҹDtHK����O�&��w�?��{7��q��(̽�H#jȕW*�I�׼�r�?���2\�.g�z��/fV9?�m�^OR���l��@e�.��.zy��U�� �"���Ͻp�;�A��%���#h���c&ّB,hf�fG=>^)�9�g�rv-Q�Q��b����?�!/�m!^ȧ�#�:ڛ������P:��,���54˿$S�
6�2�j,�7��N!pT�ҭ�|�5d�k*"k&�,�4ǧ��W?��>��W5g� ����Z��U����F�c?���Y�|1��A��M�̲S��^Kori�
{�"!�
g��&���#����"Ii���0�9^�>��j�[^��(�v��~P�!bKi��v�1�C�WiUe 24D6��*���2�@r_��o�,��neX�`"gֆZr���>���	J�M�m�xw2����԰��Z�͹B��d�0 v�
��]+v(L�Xz�9^��F�r��a��O��&j��5|�R�
2V�\��iP��R*zI+�ALkKd,���֯$��}(ug`�w[;�J#��,0����0�TH��Х��'}Vj�*.I�(N��_�:�I��T�g�l|]w[_tÐO`��Z�
F��v�5 �ԑtY7ƌ����1��#�o�[�?�/?u/�|<�i��J�� |v������'otx[Z��\'}�"�<���W���v�����:XoԾ=��I+Gh��/�	b�q�&N��8�g���%w�M-��T8k��^����0+�e�[�;J7o�:#Ӝ"��Q_�v�e�$ǈ�C��p-��qsr?=�)���Q%9�B�4K��\1�C���M]��|)��Fg!����d0��o)��D�����G����[��X�a�b"I7%���p*F�E���hO�ƙ�t��a%(/�Y��⿪E�{ٍΣ��>�l��S�ف̃�,���5Jz��l*��
��,��E]S0)�W.@#��ʺ�ׇ�cr|��~e-��5���?�0E%60��rv���?�s���6��Ɖ�#��4�A�W�TMa����ԇ���a�b���}k󑅊i>+[��v�j'׍s'{Ά�P�.���GT�g�����_����A���>����Tk!,v��3� *�G�I��x
*���zb}`�v7�{!�)��֢&�O�${i( Tp])Mӭ�]Dc6�(�E^��D��
�M)��L����\W3�A,��$P�!�}�������d0�`@�a&\
�~�0�R�`���qA+W� GnUm!�NV�p�o[a�e"&j�ںo��G{�!�w(�ڭ��4=;>j�N�1H��H�ᅡ�&v*�:��J$��U1O�cmCw7h�⩢�"	.AS�.��(vA�x�O4��%R}���	��7��^�7 {`�Tq���U��X�����X�͹Ma�*^��ۧh�I��u��}ш�0CrSՖ� 0���?f5�v��O@������V��o�d�C�B�'1^��\�Yēa�\�0o�H�!�%��)��7O�[�d��ހ���j��~S��XK]݇X��C�Z�(1�%E:�?F��{}[ >�F�~�ŕ� |���㡜�a�Tu�/�D�f1s�Úl���J��x:��U4r$��K����ɒ|�_��Ҍ���_����B��z!b.�<r¹yA��_hZr	���O੒��h�0����Kn��\�;�^���n�9�I��n��Oh�_�rTT\5�S��J�)�|m��˥[��Gh�����0Do-5y�In+!'<|p![����b
�Ʒش3�PC�-&ɍ���<�@kC��7�,\�тs���%)�U6⍻-ڽ@A�1��~���ϝ�,oP��HG�~�Y�t���"◩�|Lx��+��<a!�J��Cd���cÔ9ҳal�,����V�����j�V���퐺#�!���1�%�"�NT�y�l�$9�߀B#>�=���b�c�څ�k�v��c���*
��%��{V(&k�Rz%��Gc��3E�ܞ}d���P�c,,��7��W~���j`|թc),�4��NY���]8�}"F���e�1�����kp|P��*x�)K�^�Y�a�����)��?�}��!��1�[�|�ٔS鵠u�=�aT��h�ڼNtZ��{��
�z4*�t����d�r�tJ�x��4)Wb�Ln�$�3�~T��oY\L��K��Z�h��AdpPa���$��������Iy�
z�n���D����6�g�2�h$9�� �d�eV��cV  =�DK�j�*K%�\�u|��'���(�9����Wu>�����@d����Dē�3oΡ}Ԉp�՘�:�s�#�@����Hs�U�`j�|){-��6��C#Z�3#LB�4��&r�a���޾!`k������g�=چ�B��o�<�~���%����.�n/(��lP>�¡q�/)���ͱ3������I�~�����3��P>�߷G��F/������0�9U*�	�F%�v��?-���̎��a�V<�9��,|�ws��2<}ꖀ�;��dA�0�T?�\>�Sج�p�~B�nq�����A%�<��� ����y�(�\ x��.X�A")���/[�x+�>~��M��(_ᰴ��C1�Ytl�O�����r��TW�;�G�w�ò{Sm7�C������q�[B5$a�d�M�9X��"el^�\�9-��RQ�������5̋�B0�1�!�Kׯ*�
W��ƥ��(W�ގ��<���_T#`yt5�*͏/�Q�d�����p��ꧧ[2���E(�X�u�+"��J[�p!\�Rb�CYl)��qH*#���FAj�
�EI�K�,���V7Z��C��T�"��[e4�}Y}WT@+�q������ïݲ&A�b>_��f����� ��c����V�tB(~u�G�K�џ��ݜ���=輴L�AC��cT����賰,ۛúw�p�"�B��Q@YX�U�o�J(]�4�JG��oЍW���4G���|}Ԣt��mPL�E�V%K�#l���~��Z7�zֱԫ�5=g!&���/��+����m��U��R��/����o��l%DY$3uMVȄ�Z~���=Ub���RbJLm�}��|_��ld<�S��I+�c�]7:s�S���Y���u��tD�o�ֽE)���0u[p���bE}�pqs��h5؅*���-)9>)���EpV��u#4��O�{O�����`�_�\��^N6cO�/B�&���LxN]�ٔ�N&��Q��T�_��_��`I��1�Mg&�\�hR~���|6���J���I{Xx�+֪���gek�%E�/�Σ
�ud�O-��u����Vb�[��4�7�t��g�8V���P�y����fn�
zd�˨�
�+F*L^�ur����s"�ݮ.�o��r^�k���^+TSِ��j��"�d״)S����e
(�̯�#�>3V;_:ǈytՌ쎽�G�d�{�ߺ�ū`�[��3Q��.H��!#��H�ڡ�ɳ���25S�K�!�j�1���z�������}P2  �r��"o7�_F��xkz��^:z/yq�G��i��J��g��+M�{�I�$��į��.�jf�$����5��3���#Ԩ=^��#0p���\�}�~/A��3�@�9����,��'�+��x�b�T6LE�c|ߋ ���R�"��x]TZZ�W֏�<��9Z1�1�TOM}�A�°G����Ā����j�6^0L|}�s.�\Up~o�9� �V]�{y��Ap�6v��P�m�7�S����i!���Yg �Ȭ�o�@l�j_�Z�X��S'�m��
9� a��OΙ���(�x�{�Y�!)oN}O$ٗ9����sE赣�,dW�0�n#��	zH��dO���I"��-/�Oށ���uL���Ǟ�3��^���I���_E��8�.�-���Qq�ɿUDS��;�M.�YXˡՇ����94�߹�N(�y��M��
�X��Ձ����4
g]��� b�ގDQY?*k$�	�G�4�f��sК�(/��^��>]��SGWe�=�ٿ��@5�H���.��˂��L�f��TL9g��H�}�"��q��-CO��3J���H���A�q���v)�ۅq�/Y9���'���z�Ӯ�L5E������}Q��|�l@����t�P(�;�I^Y���$F1Ѯ}u�Q�Q%4mܧ	��R���-2��F��:�Y�^�����;S9Sc�75^����w�z��c��um�Y+�1�hż���{��OsΩ����vO�&zOZ�)�|�$rQ$�0���]ަ�QK�t��0�2�pu���.����&'3]H;�[�_�)��p��2q��vJ���`�~�#]�X�`�\������(ػ1S�3�O��"��%���@����@���\�Il���Ŝ�o8�����o�U�l�R���m�����
*����p9���t�s9��iCx��l��P3�����-
����{\�O�^nD�`�@YPK�������\�����`d|�����/x�q�'��GH�8������sx�3��ǳ���:�}`p��JgM�Z���9Ӻ>`��
�&��:�5��7��=�6�ĶŎ�@=��Y�ۛ#�x��w�P-��}:�>�H2�\��]X���i���:�����O���1�W��^�n��O���LBp���w��ZA�c�����N��f�1 Z_������[//�ّ����d��$F�6>0J���:��k�˖v=��y�=�wKG7�� ������=�%�8��Yan"ף2Ş}hd#��# ?3����V�G�Т�'Di���oiROek�U��c8��� /li�+.�`5Ȅ�H����4|8��g��i����2���Y�pF���#���۽�{g+!�-���Q�$�F��s&4,&
4ٶ��������33��tw��EWw7�-䓫�0��*�t�T��ɕhr��H��2�GW��� fm$��x�L�I����s�h��
��U����8	�>�`;kXN7xwu���Q�mI��u^��܅���6xt:�
Re�w aL �O��.�σu�#s�*1Kp�0�9Y�e�#d�ͅE�niUz#3�, %����0S%��C�[�;�ԏ���.�ƆЭ+ ���5�{O�ޘnM#�׼��l�d�>��SBR�Я�x(���Ym%��mϰ���c�8�8��P�� ��-�/
�GRl
���[��*}��������GݖHsh��q.�ֺ�;����8k�	%�W���hΓ��W����������2�i[>|w��=uOn>�U	R~���C����˨sE�q=� Z��#��ѵ�f\�y���ߢ�u,61�i�1�dQp�P�ײ�%�RPI��s�[*I��M�g�4AR^�\�KG�����m��:Dѱ���/�����F��fN�l��1lS5��L���8�`RH�(v8�#>���㼤��ܞ���G�x�V-����3���	$r��U��>Q���$�xI��/�wjHo7b�f�d=[Q�xMxj4*&���ǯ�������q�*���!<F�+g� ���}��#C�����owyVj�H���g�jeL�ǻ����c��징��M�zKb��ꓞ�q킦9ZϺ�Xz�=p ���$�x �	���{Ș���mQ{n�S���!��1��m��b�1� �*Qe�TЫ�T^�˕cr�Ck8����U���L-atF�{i�Y�$��>\r��2<[����p�gC��fM��=����"z�7*/������T��pi�ˍ8~Q 1�w�㒸�	�!@�wM�����GaH�-|p�~���Yg��Y�P����I�g���<0Qd��R��[}����:�aFh��N#=��z�"p��%�3	�Z��t�˼���(>*P��Ē��Wt��x*qY��"�~�T4��.ģ�"ìF�#Ԟ�U��H�N*�c�G8i!����P��rZ��v}c��28�}4�����-t(IN��@_L��爣_@��=A��� KL!�$gmLd��н�H�uK�z�?D�:�6���UWށ�о,��~�`^�N����(�{RǱS�PQ3�N;�?2*@�kd�q�L�+�e��gJ�7�í 3
��l���_&y���Ζ2g[�S����	��d��XX�R�*�L5S��ʡ)�Q-�W������;��*bŁ3�]ȴ�l	J��ްz�3�Nl�(�v�oS�l��h���#�לe�Sk����5fC��__�����0M�[h J a��h���D������C��~{�������.�,��գF,1=IL�dg�7Ĕ�~ތ��)�7��U���
�*2��-�9kI������d�����,j�P#���@.�-�' x%�P,�#����e.����:�ؓ�_�Dsty}s��!V���^pnw!VR ��&���<+����4��'r��;I;��?@Y#��u�9�#���7&�K���OF�#L����/7�m�����2W��~{��u����շ�P�ŉ@v��[�8Y&�/�^���NPuU��㉳ťW${�B�5,lv����su�y�����B��Ѹkc�o�
%�����+�j�$�$�%f�(���B�?�E�J�k;F��֑C��Լ��=��?����/��|X��_�-���}����DV�4�_�^>˻�+m"4�A���!I.&xe�����Tی��c�v��魷�mG�;VM�˂u�~�R���xnG�p�	'����q2�32)B��d5�w�\�D9��c����s]<&�[�}a�v,��ij�}�3�,j��6��Rw�|�z���êxb�\i3��,�c���ޥ�=��+��{���d�n�tc�>E�h����_�M5��:��#g�Y6�k�7}!���>��7����|�0=�a������u���.XV�8Ł��@�V�sc�� h3̹�/8v������ݻ�a�+��P�L.iJ��0�؏��i��#��AB=4�chn��s������Er~H���?߷�%.3`ӆ�!َ��qV��7exE,S
I/�~T����Y�^-'}J�1�'�r'�V���&�b��>mjk�{��S�7z�>N���|GP��C��lmk�1����"��d��d�kq���.SSM��r>u�ͧ1I}/���Ųn�������(����JZwl}�Z�dCj���fp��N�(w��"�w�ZET�*����&fJW�r>���gT��O{ui&)�qc_L����(�d��':��n�Ä_����(Jگޑ����v"W����;����6IR A�`�����J��j9�(�dÓQ.�1�<j|���5=y�O�a����-=��{o���e �����tBOo��l��h���Ru���"�ñ�Ű�W�J��%����q�Ս`ϣ@{�.w��y7W
���ܰ)��f 1����J<��6[i:̡h���E�Y�Rպ��}�$����\N�Ǻ��M����:�d�f�\�����ݽ<�4'�l&q;5;%Cr���QIG���T�����:'���L8T����/J�<43�}щl��N�[K��]�����^4�l��M�4�8:4���9G�QRsQ�>o��,�3� C䝃��:.�o�>��i�wz�0�<�Et9wu�!:'x**<��tNK9cM��S���LX��e�H$��G���>`�#�]K.k���x!+��&��U����T�N������g��Bs,��ܼ>�j/����n��k8�̸�j�����|�4%�;Z4��6�f$v`�+B@�Q'��@��[A����H�v�������9ʡ>��$�ŗQ��d�s�C(�v�fh񀷼�<�XN']	��)�F��Y!˄��FhÎ.�l2���QF^�+��sK�%���
��9�q�JjS����[�����݈���4� 6P�h��Z �_
ٿ��@%�LK�i����g�P�]_�3�\��K�Z((���X�>��ԓ¿+q��5���CyPa�}��t;�#�h^gj ���=�f}�f��o��ay��"����RD��=�j�ӹA��xN�u�?�3\�6㼛��kf�난�<�{ =��%� \l�jE�����\�rO�F��0���T�V��mg��Q�'95�@`����v��2:5��0��	����@�I3������G���]��@�ζ���M��~ŏ]��}���-@T��$�����v��>��dĈ�_5g��zoem�!�������t��#��"�s�۔�Ik(!1��7���k�m��˲HJ��x�P	/�(������0Y7�A ��U��i�^;B����v�!�g�e�='�Zv_���lW��=��L����P���N_$њ��og�Qߣ�;G����"p8ˈ�Y �?=栈����«{hU�#<t��t�vB��'�#Xg9�Sfa ��� b����
�L_�	*їF�� R�#�cIʋ��n�	7Z�+�R�{�Y#},��C;Ms+r�B���e'_��ږ7(R���ë�}]���ǻe��-��HF3��+l��A2y��+�(�X��gBc���u��Nߋ jF�>��+��f�A�c����Y�9������*�A	�_�K�<k�t�͍+�*� ���,�%�X!��fؠT�wd	]������`����S�#�?���k� �Sa>���u�Uy���ad.�<S?�q܎lw��9� �\	A_����P�%^��i.�"N�s�Q�<����S|��S����J�,���>�/�g�W4�P���QԬ ������,���a3�e���'v�q!�?���F�GD�	��ב�v5sh �J��.��J�V����9 ��bC���حMJ �y;��l��1���kA?jUÚ���'-��p'���芘*�X�Ȉ,���7$[��.+:q�~1�\���=�*�鰅�&G&�h���[��A:�g��|���ȶ�cu��	�n�q�z/=k4����2d1�B����S��%� 碘v��u�'S����h�Y/:�eߵ�������$�v��<�̸J�{f�`d9�|�,�4ep�7����vȐu.�+�&�<�q~�M'��D�旾u��/�X$AW�-���9�,�߷r�ߞ�AV�-g+}����(,Y��??eΤ�O���U���jB��\�f��J��w/Mz����Tn=1����r�
o�n�<U�#:��l�!; >��=V�K�o��g�%p�9.��.Þ�Kh �.���)j
�i�s�����RRl812���>�2|R�n��z�Z���Ru�)��#���{�r�z�``o����k�4�Z��q�{�9{����Ы��_~�c�:��J����?~�@�@�yMFw�Ƅ*E�  ��ty��������gN�
`���͟M�-{NT�&�a6{�r�k��8ē ��%Q2oI�kD_3/���p��P�[�^e�ީ��l��_��!?wF�FuSKҴ;W��7������J/�j�ul��~�_��9(T���IM�I�=���Рۃ� ����|�]a�B�۹�L��Q�M�������:��Z�P�*}\�w�S�r�K�%�xa�ƴ뗈z=�@H ��B���/E���T �"�q�K��Av��4��IuB5fJʵl����t��4�ܵ ��ґ�� �{+X�Ú������D�����K�./(��h��&#l��Q%�-̀�>�zD�����ɿ%K�9.t�l'p�lsa;�N�|[�R��VWV���3�¹���=H��aKg�2Kj��a�K`T���#��/���y���[E�t�8�L,�?�###`|����kխSٔGD�`23��q۴�DP#��3,
E'a�ڣ��3����W����mߊ�O�Mj�7���8K�]�N�a}�?�~�߇�t���"���M�^n|���Ih��A�L��s��]�:R(f�*ڃl����2ک����YP��^2�z���,���3�Q`�t�%UPA���$�t�[�g>���	<��� �͈���Ɔm�Q5s�I1���B0a���������Jާ-xu꡾*Ud���Y���
�*�E��U99��{u7F��(���s�}��9M���s�s�t�&�#�V�K	^�^q�7|�a�D$���t;o(c���.26K-�c���zo�v�d*��6T�h40�<� 8p3�n;+��l�Ab�W�G�S?��0�`]F㟬H
ߔ�8�n�6���{�ע
N�0)��e'zX��':���f���
v|b;sWd�=Gݠ�*�U����;i�bO5"��N2=I�`ÇBC*�uM���
\���/A���E\Nń��������b7��L���7MrV���gO��*�\Qe��H��XW�@��SH��܊{4���˹��rm6i[�4�/Dz�2S�wح��"�wN��%M��r|&H4�ԙ�<����GRh0k�e�o�2V�ߚ����Ȥ�x|�E�Űv��M�X;%��ǣ��r�WZ"~��3Q�@��q������P��������U�2\�=�Y��6�c;���H�%%�G�=#8$����+o�k	��VJ��u  !uA�Lov��Ѽ��>�;h��k�t��7��� 4�bp&�xfހ4���{
��%�>��Ϭ��k�H��,���M�q=�7�:��r�s�K
v�q���sL�b�A��ݛE@Ya�[��]��_��ݺ>�C��m�y��Y�m��F�U�QSݔX�`���ܰ���;�&^�M�N�����,��%}CT�j�j�G>��bF�R��2�l�v��Me0��xn�z��_'����({fm69>�Ǯ��P���u�-�ŽtE�����X�����h��\,�U�tE��2����`GN��`w*�u�;j$�49��ʏ&o{�l�s%�o�S�����۹7��%}̜��'�4i�$&�?Sc���?�sg��_��{V�(51��
A��<���j_a�+�׈����	{�f�M�P�&��� ^dRA��2mHl)�P��b�\0��f�^�j�����K><�#������IɧiPx�?4��8�b��H[���+ ��0�%M�l����ˏ��ˢ$
\�e-��T�����J��.�D'C�sp�x��Śp���%K��Mo
���'T6b�)����nx̢��6�L\�nŰ�a����Vn��=�>}��D�t�.�j��b����������b�18�\����~����Rƛ��6��M�4�<��p������BP�ĵ���hOH��.�KUVP���Y�� K�ɐ�^غ��K=FY�̡�dqP�B���Uҫ��x�o�s����"v�z��f/+b��=	Qgs����ej_m0��*t'Д���$uǭ}YXbi��-?K����f
4��v�4&NQ��Ur~�5����@�2V`Xh�ƣɂ��wz�Np��v�Q�����0国�e�����{ �;�E���9�I!L�!���tz'1e�����vXj,`Ϙ� ��<zUf��۩K
�E|�b��Z���(� YX�j�O��$�k��I��a;,�4�!s%Q�ڻ�B��d��A]9���gJ�߅���Y�	�_��1�Ym�[�����,q��A��Xd��1��^�2����ħ��"D����ؘ_G�胔��n�ls���-�n-���;5�+1�d��8������$nk�D��#����*#7�HG3c!a�e!�=�_e��/ "�f�Y_D"c#e_��$�)c���i�}��:X[n/� �N��@q%�aw%öX���N�aLW�UמOk�W���tKi�pQ�Xf�/N�S#w �j~jl����k���Y	M-P�q��]۟�E-�r�\�n�2�{B�j��j'[����'���DN	�7�����@��[�z�'݃�쩼�},�Ip���~���P�����Ӟ99ɾ����{N0_W͢��9�� �8k����R	�W�>}�ꖂ<b��htu�I:d�عl��G�ߖtj>��)��¾�F�%��`!hG�����Ds�X ��msV+���a$G�Bb����tZ�l.QsE�EyV�����Y¥����h��r�~��fiGP�ٷ�&�}��Q{�
�:�#u�(OV�� �EZ��<ZŁ:�Y���y�he�\�4-gۛ��G6u��P��;VE)�>:�+%Ć�7k��`�}���ï��
���ۋͦھl�w<H�n�C��-�����6���-E8@t.��ǟ�#�7^ɜ
�!L�t�M��fh��u��������葖%��8R�o�]d��Q6&�!�줇1-$�D��z�˻�>��E��S�0*�w�h��X>���E�Lo\9�H ��P�5Z&a�5`�D�Ol{�)�'�(#m�n^ܐiI}7�&H82�I�S�p,
Yl�����Q�4�;?�n����'W�/CM�K��4��ɻω��=+7�B�2�Y(8���1����[�c"�Ǣ�0��������>����
v�iw��e�D �פB�n�y�#	�{���m����&=EA���?�p�)P-h��t1�Z��\00nhI@hW:�+�Ʉ�?aF�zV��%�����ΆBc�Ծol�O�YՅقR��f�qk�˖b��T�A۽ƣW��M�i~���^�- L�T��w���>�%!��n8[�P>��gJ�ʣټ��"Ċ�������W{�}���W�ƛ8C��l���3_����i?�z�#�ۉE[�R&�{���{w�4�[�C��a ������K��#_��T��`bE����-D�����,Yn��wu7��|[\�|S�['RZ����v�J�{B3��.I�-�t��Dt<P��:S��?%Q�s�=���9)
V	TI���9�D�8���������� Z�~�J��o�f������<�V�Ea)2Б�ܲs��p�-�D-���u�5+�x��I�Qׁ�q�9��� ��걝AU`QQ�$������Z�=M��'��ej��Go�
���ΙQ;[��u�tE5���8S��|�2EU��X�ހ0� ��O�� )�ƯK��M=]��V�z�q`���������h���Ҳ�M11rͩu�'��+
�eW���F�Q��ƪ��+H�����&�J��;��5�!�6V%��rs��S�+X��YK�;M(wk%��im�	l�&TW��3�d����)�T/��t�5�PRBTHd��Xh����Gi3Jj�kz�	�j@�&n���}~ʣ��6b��a\&%��/�p�F<�.�e�9d>�o< w�]Տ`�YO�	���G��>* {�B}I�M�2)�Y|v��f3��Y�E7�D�yf�v�[jh��d��#�:�Q)���t����oib=@�Esk�b�t�K+�r���l	c2�'��%]�=D�\
d_���Uz�����x��?���O��޶w-}�� .�Zx��"b�rYm�
,I��~����߯���o�/v�=e���*��C���i��Sp��#�V���ma=���[���cs����f+	����^|-,�?3�-��9�����_/~C'�+�k���MmI�\Ϻβ�D���f��h�=;M��.h�I�|\ў
���$�תv`]��q��؟�]Uӣpx�4�1��zٕ�2��vz,���!�*P�O1�.�e��83;U�2̰��׻x=U��\�f���0��q� V(��=�q�	�� %�1Hҹ�6RVRCcJ���	*�B�)=?tq� fˬ�������;m:��0eע��'{F
F��Ӆ�߰����"�m�EЄV�f͚��(c,U���ׄ=y=GŪR���5�+�ũj���ژ���O�I3\s����A�\i:|Q#)p��mzQ�u�r�{y�^/��ȷ��#���]���/�F�@/l��ݾ�¾=���ڃrecB9DK��"G���|��$	���r^�{���(M,*�VE˽��ue6Mp�L�RD�u3��CT�ꖒ������nr{]QЀ�� F9�B>�#�jt��>;�e�G��D3�����C1�2>��p1����f�-28Ю����������6�*�ԅɟ��Β�Ku_��d t��P�|ܕ� B\"�8c�L��,CUO��j�y�C'�������Sf��}�x�߫,�r��5�&y� 6eR	�Y<���������Z"3��Te����h(/d��cq9�����7�>����}�>�v�����>"Zs��u(U�Bۮ��!тkI}�5~���D #��Ǫ�����Zj	�槻��_�����;@��R�� �g5P>݁j�d4�$GG���Mts4���s��b���&�F�T
mZb��k��(�X��n�z<\��'I|r�p���I F=�%����:#�����fk�VwS�IF��ގ �ߓ���lK&������m_�S��,-���Ǥ��!t��h!p�=}�:��pa
�;�A���+��۷�Ơ	
9^���=�F5�U��{�K�W��IA[A�O��$O�`�C�G�Q�����Im�ɰ���=�1�	�.�x�jɔq��c���Bl��mX<�����U�@	�>4%s.M�8�I(@jn�v��t�&����6�Dy��
d�8O�����H�z���腳�Oދ��r�������D�B~0�}b���FT����v9��g��qZuCwu����"iFms�C�8̌��=m'�n�UH���OD'!*@�R��,�%O_Ukl������f<e��,N
�Xck:����/a95,닋���@��6��Y���;*�xX�zܙ#�P<���Eb�kG��;
���p= ��Q�9m_������,%H��	�D,G|���Ђ����$�b��Җ�bC���r�{i����͎��{wrJ��3	SP��D"P˕-�q!�pU��K6�!��i3��U���u�;W0�x���a��W ��������Y�C�^@4�%��CCō;�����hP�bM@U��f�-��Wr ����;�,;�fH�����ؘ&i��{$f[E�7���I�|{�G� �~ځ��!��.i"}�WOhkG�'�|�2��7�qF˹Z7�i����ԊJ8��{�t��׮C�7 �Y�\��UK��G�.\[�"��MmC��D���h.��vei�-BԦa���B�eu�?%�9_|�[V���n�h�|�`�Y�[� /��׫J��j��:+�Q�K�D���o���6�t�m����pƻV�ƪ��|P���%;T/S�����T���Մ.l�l��c�%YOî�`;�'s�	o "�b1w��#T�h��M�QZ�f���I.}ľ�(���'\�h���lCO�����	�l��I�KlȿǕ���Ϥ&r��~4u|�ks\R�o'b��:ח������@���24#�e�U�_�c�V�X�ط��7�51��gh(aǐ�o4��Aաw�T� �A�0�-�	rj�?�bſk�W8�'�G�w�ʖn���@��kS�>l�=CH9[U�t��M����oM��r�a]F^�����/�R3qn��m�:WT�aM8�Q�=&q[�`8�.���yO^����`)�;L��7=X���ҫ'�&��M"��x� ƕ�R�}#e�n��|<0�5XM}γ���2f���E~\rU�G���5&˹��_b�<#\[-�EL�##?m�7�>*�FTc;�BU�Q�2n\Gb������r��Bs�y0�nX�@<o�������g�T���1)�{(1�q-!y������XmI�~1&j��� ��M�.
rB*�u�����G�NR�KM8H���h)�7��jq�P��d{�[�gV��̿wN^��N�O��\���j!��G���@e+����%w�r��%��$� zL�:����&�[/qq��.��B�覓��\T��U�b���Y?�*�B���%�,m�0��x����偘��p���y���Đ9�����4������%	S 9*Y;ʞ|Sk�dI0�KK�k��~��a"��1 �����pe��W֓s��|�����[bE2yG��<N�:l/��k��c�E�j�(��#�Q6b��+����u����ɒ���Tj�'�Q��/R{�<�0��,��z&�����Ͼ��L9:���љ��Pm�`�2�ҋ'0��,�#k}#��-[�G{T�[c�l/O� #��\�٢�/4��J��v&5��\�O�՟����V��������'"�8�#0e�D�iٿ� X���\(Zn,���Ꝥ��,J����e(��ó���!���;/�5��`-G�j����!e����4�^���BZ�TL�&���ڡ�
��`~8�&S��:"�6����s�6EUV��S�3����Q��a�ϕ��������Rx'_�@��~CtΥ��"��jچ
��R9��*�qa��B~��3��zu�W"i� �PN�xz�3�v�����V�F��8?Q��p��6��p��s��|���"����s���ƕ`�f� �:��7p� r���3>L~.�,K�7���m ���j�*��t�yo��	5>�i�}h�B���r��5k��:�M���w��C%�Ô����_����u8����.s;`�'hF"��e3ׁ�X�+�щ� c��m�Ε��>�rF�<&�G\f��ƂSW��D6\a��DX|aCTob�Pj ��z� <� <�jJ`�S�����Y��z��$�E�u�"�h�uJ��ݹ��-����rI�ƽ��AT��"�%��D>5ϟ[��Y�5��W��S4�7���Q��a�F�[Ao%��C}���~��<GɄ ���pp�7ʁ�x�J:�N7���~�jT�B_
�)K��S!O��T�:_� �8=�O :�?���wi. |P�n�V�S���7��j�3 �D�-��� >��Y"�D�ER��?�h��&�{[ำ��|�	͈^E�0��EX���1����'��s��3��[-u�tw2{���n)�!���8�<V��.[.������Τ�?O�G#�Y����S9�,#�$���������|j��}�9����qy�-1XE�r94o�}
��϶'r�<[PK�����֨�D��*"�n��9+c��כ�����*p���b�hI�C����;���P2IX���_�� R�Ί�U;A~U���"�/hp��ڋX��#��V��%��[(;=2���i�7��>n-�Z�k3�'L;S豘��8���B�"P�vl%�<-�8����D����!k03��8PS�a|�y�� ��%�pӎͼO�Vͨ
��	�&hOԇ���%Gub]�庡k]I*&C�q����|,x3�p�}�	����#@���M@q�ڗ��K��C����%6�i���������Qy����`㾕�¨�O(��b��Mq����I~���u��[�����,͉��?/Vz�.b�#}��b��A�f$���4V%�>|N믧�F�X�סj��ϲ��mB���-�T"�d�b����C=;;%Ϲ�.	���My�K�7���z��N/`�� �����1/Ee$	�S�����N�#_��0�0�*&��|�e.bUO��_CZ�E���ه.��Bd���[g���L V�o�O��b+�K�`[3m.�����_�D��|^��$��������(�����Z�X�]�9�Y���#���My1h���Ø���ɀu� ���7s
�~�2#�D���=+��l(�	���W���v.�W��Tb?� ��:�R�����r�.$���	k��F{�טi�ʹ6/��k!�RG�<���7�PE&�ǵ�B��!�
Sǧ��,��d(K�o���Z�T�<�?�,�}{���	M]��zlzro�/�!*U��@��M�ۼ�5݄]�+��&���DYE}���(^�*��<H\FĈ�O���|_�%_{*U���)�^��s��8�Ё�~|*�㫱��2Pc����h��X\l�"��lT�@	�d�FG�?�g9��ۃCi�L1ø�e�g�������xUcVJ�x�;:�d!W7����������]A�� ��XW.K�B�ɕ2R\����g�8]���8p�K�I��x[ X�JT�� ;�_���
%��ݟf�4IFj�p�%�iɘ�����$-�S�t�'�Dd��C��}����8�}SA����M�٬m�'�����ED�g�5�LD�B��A*��!�\��]�_]�?X%��l5��]��8�G���+x������uWq����_��[�#�f�w�U����n��BM7$Y��WI�P����+�5���~�����&#�G�j ��A�<��������	7�RF�xX��JE��h���/�m=�~ʬ�6g��px� ��כu�3zˬ��gG/b��؍����<�|=(Nì��J���+,���-KA�6������>��"�8W�!O0ȭf �B;@O���������]�6�F9�ĩd�n�ʏ���Cr:�p"A����+�o8Q��s=s��6S���Hi�-���'��~7Ĥg����-٭�{��P�3z��u�1"~��܇+���!N����5�w5b8�rnhp4ȵ�?d�oKt�R$�w�D�W1�Dͥ�D�Q*��8k$գ��^�0t*�Hb~-���-~�Yd���@���vJ�"�-sF�'�i")x�Z�<���o����#��0�������%߉��{ɧ�í �a��|P����Lg� �1���F�����?Č`��E~��g0;�\�UE ��=�lZ$�\i��ZƔ������PL�x�l����b@����� dkd5�I�qR�ÁDObi����!�c�w��X/�b_����`�;�G��_-O�� ���v�y9��,���^ɤ����mH�Xg�G���Q�H�;u
���5��˟��O ʸ��56x�gBޘ1 �@� L�a��xC|���^�o�����8�v�(��Ī(5�|<{��������#	���0ɝd�j[�+6�c���)2�E�U3���;�>��d��!hkî�Z)�˷*55��x�A�H�0�JES3�4���Q�-VQ�PJ�=��U�}�1hQ�f@���+�P�%�ވ�]p�m$��s��0�G�����R�{p%P����匁M���/��^V�2�qkGȈ�Pދ��~g��=�v�Y��\=\.��W7��:��E�.��/�M�aJ��R�e%B��]9!Q��^�B�������h�rB�8����n�3�Y��k��t��4{�(~����)���e�$�����hu�<�1�n��������]X, j½����ƈKQ�:��rt)]�����Q�D���K0C�L��]�&��7�yX�֣�J�H��PƇ��k���˦rg������E}a�#`�����%F=IMɃ׬l?'�մF)$;"��9��2���9�PM]P���c�M���ɶ���w�Uh�*{�A�ۆ�23��M�x��uVI@S+���FJjy��4�f�Lj��;��N��s�A�f{Ȃ"���Z���-�]5��W�h:�\�A7���&����<>���4���'��z/�GK���bhn�����:kBs�E[�B�CQ���Z�r=��P�+6����6<���H����O��=~>�Յ�V��l+�z#'��.=?�x@��o4?H�z����C�=��i���z�T�E�d�w4�3�k�X�v"�z�42?(N#�V���0o�h|�O�ӏ���G���
5v��aN�9Iezx��MW!�w� ��4	4�����3>�:I"ϕ��i�)��l"�bQ<�n)0x]ٝ]D�"�����5f 4�#���4|J�V����N2c�\��ߑɾ3�];2Mn�'bR�������Il�'g9S,5Dմ~H)hCa���s���|��'����r_JQ�x��K�_!��Q���d��;��3��5�|�p�1��F�Kd9oU�\AAS��X鄂:`E�~}�k@YK�N�b���b�I�"vm�]�S���������xƣk�;�찁�쬌H�-��g���j��V5��AJ-�/����`o�,�G���'�.��7��h���^L@G�KW�h�@��"G\=v.&�u���2ALŬ�/�g`�]QZp��|�n�=S5�
}F��?K�a����`�grݦ��ҩ*�+�̡���.gl)����v�>ޒ�ý�1v@�#3�jޘB¯ۻ�����$�Y���©Z�����mV���1�����UJ�df��R�.�q�����ee������Ձ�*`�l�6"��w��0�l�h���)O#��eiƽ��Lp{Ԧ[�N��͹�x�qfZn,���G���T��(�[�Y����s�s��Κq�j�ޒ"���Ɂm��[���fs�;�b�QӤ���I.9u*.T����s�59��"X��y���
l�)��o}}�*�0�
~�6�b��$��$�]rD��X���6M��E�zl�	��[\I{V��G�\5�kڋp�d�Z�w|)�΢�����-D	R�����e������Au�s����<����Id�e�I�3����Rܷ�.S��J1ԣO��,��к�!��7��^e�����n_}h�臔ȇ0Ugk�-�������EA�,��=9�#s�|��o����Z�9����:$�!@�F�s9gZ��cޗ[�M����rƒ˞n/��)ˍ�t���}��&Ɉ��ē�TG˰�gw���U?�W�٫��)�����u�S����`��)�M�O��)?9#��e�����~�͖�yY��%���D�a���>���z����'ލ�o�- ,�lEPMEIM�t�Xv�J��ks�H�8d?b�߆e�N2��b� ����p�l�h�|���H�-Σ*�O 4��ж�|�%A���'�9�k�߳��fs�<Fj�����T�-ϩ�p�FpW,����f9y��n/���4Ws�&��1� p�M�8�
qK{�B#�.���oTX��"�3o(�Kc�I�z����T��>B���"�>Ƨ���Vwm���g4ވZ�w�:ޗ��H�.��z���N��%2�����>�e1ũ��cdYG[5��ʲyQ�/x�:��y��蔩z�z�I^�����s	{���l�L�)�h@k�9�?�I,^Tx{k�yi�R�i`b]���
4.��=&��y���R�5NČ�	����;^��F{-�kU��e�Ӭ9�� �9�x��������%S]�H`o�Q3��	� ��TÒ��H��]�e%#�����@��\yb֑��+~�0��W�� F!kUG`��e��=B�6��9��1g�^�w�d�2U�缓l�Z�̬B������`����/��i��t �D�����)�R�$	ת��V���ڒ�%L;�������MR�q�V.F��7��`'B�Bܰj��P�h�[��U��5#�q復7��mIÂ��Wo���V��g=�3|�RK�4ԩ�2�+��| ��;yPC�3���m�#��H�9e{��f�3~�d<�/�x�r��S���U�w��t�-ļ�����.v'u7V(�v��!s\S51�t���.Ĳ3�-���?��e��Z�Hhr����,����(����,'���Ů�;�{ JƼ�D�z��I$��q�z�E��l���A�-rv(I ̎��i�=v{"}�m��0��raC[�	���oY8U�v���p�%��!��äY��S3�-	x_mJ�9]���Q�<����e�����دy�����#�L�*Ί��e�o 3�x1!}�|I"XH³9vk;��&Ĕ�:<�GP%؜����F�Y��(s�;co%����̲���*e����)3%�m�b�Zf@���7(��e�����_�ݓ�ՔE��K���إ�2:'��|���yR��w�u`��xZ���̩�!hV���]�*)3�ο[�_2��'�fϚ�bQg4�"YUT�s�9�غ�6��f�q�U�N��=/���i�ƳT*�v����7 ��4���v\	����?Z�2���'�cC$�yB�6=�E��i����|��XMdSIּ�$��7����r���g����1S����R����g$�DV	�t�E�v��cM����4|�<TN1�NB���½:@���� ��q�
�����s��:�t7�@�1~n�տ�l^���jx��E~�ēX5�,m��n��G�mnG��a�E��92S��s �va(��<P�٫��
�<���j	�GJT�RD�}�Nm�˚��W���ڒ��ޑP}to�Ւ�ط�ǣp0_�P?��>G��մpSt�ab�8���'A�K�jWUP�Oy*0���IFn}�+�N��[�W!8� �fir�������n�,l���3��q86&5G�0뎸����i�-�ca�����%�f1F#">���c����=,�����p�.��.�������Ď�aU��H0��;j�(s�6�4��[�y��6~�_Pc��࿅�L�jjܪ�N��f$-����(	��]b��!�L�9����' �:_��Jk^uT*~�gґK!��r�[��['���2���Vx}�h��D�l:4I�A��X���?� ����8�!�q�*��M���ᓏa7exz��@�a�4:8Ho-�UcZ���"���l���g���G	�����aEY�/MLU\׮��j�-��1M9*���������."�qOO�Ԥ�9�u��HFKK�k�Z�\X�(�G���"�n�I��WMGn��K�{U���T?��o�w�l��C	^K�U PU�X8�Zb9�N����W��Mmg�h����8�Kޛ
�0�
7�w3��*+W'�3��<��a�eڼ����+w ��{�]�T�� ��~�k�l�2�bfgW����D����}�?h�$���Y���.P�A�@�{���$�6%�0x���ۉ�&�J�����G�F�y�Q^���K>a/q�Ux��>h��l����kN�yp#�7�H�FLtO�8ń�'�7��1��[x��Z�8
/��!��l�DDjV9��|7A"g`Y�ã0JHa>����	�\�ҩ
�����m�n�'���Md�к�?�W^�4��셰���O/:�|_���
�{��8Wρ'�v�^e�踤@�p񽽇���w/|҃S�X�TF��>����uN��~tʫ|�S;�2�����
=��x@�n��6_۰A0��xc���h��Rڑ%���-�X�(0�Q���D/���Nts�q���z��c���q2��1"����(����ܦ��p^��D�+��lR�Ǆ(Y�g��6��
Ѳ�^�P� ��48o��VƃM�t�w��!��x��0V20>���BU��IԬ_�'����do ��!�8%S��%]~�B��v����w2lO����&b0կz�r�����sj�a�Ӷ�x�Kv� ��}���u}8��Oh$$�؀����9'����l� 2��8+��Z���QxJyq@�Y���)���m��	�`�G�3B��Fj~�\|���(���#F�4�g���yAQ?���)u��U~������������"�ey��ʎ�m������׈o%�Gز�#���*#�TX��<\u��F����i�&e�� 
�����*�i��~"��t跾6x���M���ߙ����pV�I'�\n|���\�+l=�0hv��y�`s�Y��3�*�˓#�	=���+J1��6 �iA�ʐ2���z&�0B�u���xͧ	�Q���㎯"(����D~�`j�2B���d%�M�I�hz�\�Զ����P�DC��г�M�O!�~+i�h59e�4�mPG)�̌p�lA�o�"M�-=���#?T�+�R�"�r��Q(���-˄>w|"���Z��a�d͂�UMG���w��>�!�u�lѲ͹����G=���S'��Sr��;�(�=^����p`sDH�mT������K�-H�*1AjjI=��pK�̍'H䶹2���fv����Q�x��V�υ�2뉬M����X~�4C�0�-���"�H T�?CGVr�+��/%\����A��í^{�|�r��<%���e�#��-�1Z�	E�׻Hgm���FQ����8��Z�v�9e��S�ͦ�M�h6uR��hia�`A��+d���������B���Ab�S��5!ѓ9C��e}"��-޻�6���r�>��T��Dh�V��޴\��S)+�,��lN�Z9+�:�oW��5w�#!"�T��JU���rj�?� ��H�;c§	P�����Z�1�R��+f� ������j6lݹ��ܺ]�Q�_�i�U5kJ(3�v|�71ȭoS�����4�0�r����~��\���;�2���9_��k�,�3��:Pp�&D�C��=�F��=&�qй7�y���f���Ur��ׁ�*ٮ�2��s�pl����M449���!����3,i4q���t+�n�u�|x��e���g�����~��dӼ]*���ZyX�F�:��ze"3iޮ|M��߁��W߉Z�xE��й��o�ӛ��e�
�;I��GN�N���Z�ۘ+��#�U������v���Q=�M5J�N��{˪}��'s��o��GV��@n u=,�]��XBy女�x{�\��q��7	IPR9Odz�C^E[:�Q�9.�Y�tӯq�@<���l��Ҽ��mpwŤ�ՀTW7Ph,��L�R�Ɨt�"�S焠v|Ύ�0|�w�)�Y
T
y��}�Kγ��h����,4��[�,b1�+F�Ǟ�!�A�Ȗ�[֗P}G�b��!�Y ��mhiz���aP�K��#� ���&~��@���P	q�<�f�ު�Gc��T"Zs�}8�>Ic����a|ԩ�Qw"E�[��`�a3�6�Xy3%o_BjXVk���[	q&1��㗖4�r�.`3m�� ��˲z�_0�Ӊ�]�
�ؓTY}D�z*H��~�4���x��|�딩�t�Id����ҳ��&\w�8V!t%�^z����s�9yT���n���!��-N �+�}��1J�G��k�B��
���Gs�츽$ܨ����������Fj`3��R��%�	'~���a#dUx�ޮ%R)^�Gd��v��t�u)�4�V��9��cJN�=��x_)�9�^�N��@��y�#�*&!'���B�3���H���G�:�%6���2r��d���޺. �9��Z�=�R��/ Cq��H�I��s��-�a�E��g�~h˟��Կ�R��;�V�"	��2�[^�,�v�Vƕ9'NK��"��c�N���s%v2�bK5�A�LJ��Z_Ng$���s��q���#�4�J��=h���d�([�t�~�jģl�&�V}�u􈸉f1�/��@m��aH{q���i�;2^��j�ܘ����8�݀C0��ؤ�e�?�&��R��y���*��kJ�t��o7���9�#j%���!IV�d�T)��L����  �|G��1~��ޯY���	�/�ެdx��<��r �{́�/a���W.p���n���8Yl_������v�dGy�i�=.��;I�p���B��q`�b]J	��4�@����M=�m*jԵhjX��
x�V{�>k��q�W�p|�,�=צu(���KO0Ԕ���t�������E����(�5$ha�:�M�����=��ex1�c7������f�]ɢ�kg1���)���.�J�Q����H?6E�t��!�|+f"�Rgk�r���m�(�ü���ρ/�;) �#��I��f�	���*��&Jl�L<�1�JB:�5��p��*�6S��� ���gU�hP۽�ґ\Jճ_�ǆ���Id6�Ww&�e!�v����t���g�7�"W;�i.�淅��HU�yqBv*+#<r�@Ⱑ��@�I ���`ٜ�����I��E� �]�Xz�n���Z|�Y>��U0̐݁R�n�V��o��1%^	���	pD	\�ZH��GR�[��k\�۔ʆ���!b�|*f �wBl O�~;�{'Zb���@.`��~C<��m1.��?S���rìۀ��m��N+�ĜcsO���C�&��ȍ[�]�=v������<�(�{�6���a,�2ͪy�!Y�V�p����xKL�0rۓt*UxldB�|Q��#�B�N����5Lj+'��0��C�1���K4s��t�*+3�e�lj)���xw�����A����L��5���~7�8�m�Ē���B[P-$#�m�"�.OŶX�Qo���o�|��{J�ۡf@V�荌�[��֔T�e�2p�C�$����c�-�]i���Q��I�ޚ_s�O;�(/�j�tG| |r�����E��R�D��K��Yw3��ųIv9���e�߂M��5��5�ŒIL�U�-ҫ!�D��e �Lop��mvt+�D�a9����o����JO�{�z�+P��I��Ƨ"�C)%4D��27��I�'3���v��������S���;���iq����}��-I�y�pKn��u��0s1��g�g�eW��R�m�f�7 _���fI�Q��˧?���N�V'�����[�ތ��o;��FFu�@���+�|�/��B�����NfB��*�wб��\�xc�y?��l�ׁt(7�m~�|�7y��#���W��͏�F����]
��1��{�k�p6KA�'Jq�K�y�;\;Ǧ�#T��Y�Ϸ��t�`b8�8��1�v�ؚ�ۓ��о�ߴe�`nH��u�M2��/����ɴ��Mr��5��6�P�R�����Ko���͈��s��E�J�.&�T��(��ڜy!�Ţ�W�������)���^ӎ�H�I���iЗ"m�m�ݮ��&�F�1i93�����Dc)V�Ӣ�J�P�8eB�#ȭ�V'*KN����Պؖb�B�����i�$��\uVtƼy���Ƃ_Ғ��7����$��O�C�O2v�vM�D�{�8��e�&F��I��d�M�	���.�
�ٸ�Ԗ���;�ob���c�נ�AA��t��� ���ńј)c�yص��g�+1����=�����)�}�Z���޳����j%�ͮ�03��r>�q=\�ȇ[��B�,��{
	S�R��
�w��1�]�B缧@;�#t�$���h~��!��<�F_
�>qe��%��2K�+�dB�rئ��*�:��v���%l���j'�~D��LI:螠�O<g[�1IuO��^ۚ԰+�S����=���ԭ�E1�h�e[��J��VrbQctչ?�$i5q��ŗ�=�7����FF�
��e�A��e��#1E�qҽ���$V⃻d~3�(���4�Ƶ�,�r�D�����ǩc٨� <�*�D��:BA����7�f�jqƐ���l01�k��@�̜3*y(�VJ�����Z{��Ȕt�P]6`m&�5$N�����~��vZ�J��4�����燰��,y~��C��ͥ;j�����J2d�%�L�	`1I��Y.�V�ێi;.=1�>f��x��.0YH9�U�i?3��J7^�:���k@^<�(!�Qck��M�5,¤���/�B��><��"�0L$���i������6 rb#8���ӽ�B3��
:�g|��9[�C�T�	�Z�;�}��EY[���o�b�o�]��#� ����h&��d��z��/��>pM�h�t�� @��׽S���U���C�}Ȇ��	 �����?�9}3sQ��5j�� ���������f$�e�eB���/m�+�S����b?�ɋ������9��دp�4��������F`y�hU���_�Q_6U�٭�a@��ә���I����px�c�|-�v�&<pUы�è�L7|T��� ��{&½7]\� ����>�:�زO�)Z�FC,a�5vo�0��	ݔ�yͮ�¾��KL1D�,����;|�������o-��k�c�'�d3���w�ͦ�B@�ц*�F�d^X����ZA�uA�t�����q�
/��%�h'F�h���7C��s�]?�����/��cC�qC��_8�.]�m����n��C*�
{.���Pp�t�xFG�N#���c�Jqt؞��peU���w�!���3�� ��u7n���cjF�':�i��`�z�׾k�q<�
��5��.ݥ��DK�u�^T_��&�,v>�t�4P����ޭ��=��t�������Xc$�>��N�"F!e[���:I�A�k,Ԅ$L?"��˭���5K�@A����rSR(��̍����+��r��Яa�(�J�U�>;4���zؒ��� �G�)2-���d�p��^���4A͌�2����^����Mb&'9�f�q�ߪ7OPލ� �^T��2���Pz�bũ=��C��L~��xd��J2 �� mks;��RŲ����?�h#�W���@
��t��׵i:�(y`�VFb�8�}i5�S�܈��I͡�r6~-.}�?�)f�g��@��R���0���}�}2D���:kƑ~6QW���X+�" �n��"��\Kl8��V�=��r���j3�Cz�ע��sfM��g�{��2�]1FrG'�|��e�`�+P�~i��>"����6U���ㄢN���3����S�� 4l��Mvdl��x}܁[�U��B�͝(<�{��I���ZȒܲT��|��Ѝ��4�$}0[�-_Đ�b�<�F4%���R4�,R\�,��>��_�5^x�2_�rJ�o�U������:��wy�2H+{�:3ч��#J6�]�y���#U�-�١�� +��mJO
e'�c+g�z����{J,�>|�'U����2�꺂%�[��ڔe��)��#EJd����}x����h���H�Zͩђ�Iʊ>H�il���<����D�t}��� �k���J��pɘw��i[n�������
C���.m��E;�I.�*#ֿ(BB���,<�'H�*=�������f��Y,��>��d��qᣖ��%9#���E��B7��т����Sȭ�� i|�X�`���N`'��[n7�rEn�������ə 8T���-��3B����͸�4��w��r]�T����L�Z���Vy۾4�������9��e�2{yzԒF��iI�e ��w �&�����K���1��V�.ñ��x�|��]P��ϳ�&8M�b��d�{�`Tx��&X�������S���&��"/��jg]J�;
+o��׈�`D����H�-'v��_=�c��'�-�˿?�a�ͳ��*��e�#;�I/z�Ga$*����t�"�n�R�BЊ$Ҍ���j��u��s��s��&���2�:�J 洊!,����%�"V�~M��}�!������]��O����\�l�jMi�1�><dA���X\�]KZ�z���ɀD+T	�t�Ϯ��#h�`��IG���+���|�Q9�~��nF�PϪ��gG�b��(��m`��Zv�#���m�~��p�t�i�p�)"p�?���X�㵧T�dQ�O6둤���a�e������Gw��5�2
��$�{�(��7aSk����"_U@�,O� ����T�7"�XI����jل���g���f�r�hPj2a�]�B��60�ܖ�5yz�+�k�޾�@�X3�Ǿ�pI���o�#�؉�-Y�{ +��&���^0�:J|�<M*���o�>�V�?��Tw���mC��xs�lt�x�0��z�6��*냸��Q�C�~׺�=�T�c�<~+�=6!D���a���FNc,^s�<s�8��ƅw#,�����\I�!�"M�@����6��$�P$�Q؃��b������S:�Bk����b)������$�%�l�,�9bv�(.��j��m�-@�w�.@37&�(�ёtȲE6���f�؅��診=>�ȒS8�qv'�lX!g�<�~ݏ�s'D:�L�c�h�(|�W�� P��%羸����+�
9)�T'�=?� -��E�t���T��	<f��n�Φq�T�	Gތ�"E��1p��� ����W�\;kb�"Ɗ
�@���~fZ$}E�/L�Tp�{���:���he}��|l���դ_��*��t1ǧ?[dL+�����L����`���-���H~�:�G��QwYǥ��&�$��&qw�D�/�F�0����x���y4�`R�S�G	.C~�����#o2���f��qh�3x��+�Nʧ5����ݶ��:'Vґ80�b���m���"�<��԰ǒt��߻��(����<�������V]��M��
�Il��\ͩƳC?�),pv�A:.=!�'Bܹ!�Q��ii�kV�5\!�Q�eof��h�C;��T�:F�}M�q艖eh�����G1������H�H+5l%/�8��^�=���-pT�QI	M�Cd����wFW-� 毟/��������<��QR=��մ������������f~3��ʔEK��)_؈�9��ʡÌ�b!O����������s��"���*��s2�����TvwqE-�d?��0���l�Rv���'�����dT|C�
�F߹�7����FN��F�rE7R$��#0�`�b"���X�)�ńӘ�`�U�DC�tQ����d��ZJ��N)�C�������.����Ep��B����p��������u�ڶ������w�����`�+/���ͤvd�qU�T�G�Vme���u��G��m�f�K��^1�O�s$d�����Vk�����C�6� ���<EV�9;�B(����E�Cume�}.��\���l/)H��\sV��1-�`�p5�C�����*4 ����OJș�0�s(��ğ�(~��L F��GA:��σ.�2s01�M�Zy0~��{nb뢪�k� A�Vu�?]!��-�^~�˅��n�<���V���ck$�^.ak̯��Pմzg}�f+|���]]&�t�˵�N��r`{{����_P*���~�X��a3Z�)s�嶑���9���Z��%[�W3�P����?�W�>�l�g�|�03��|�d1�y�A{x�*�d�7�a��B�!)�Uy����n��u�����6F�+j��d�;7�Z��X��h籌���E�^��̯V�S���Q��N�_�D�\>r���hLG�6'��>�ƙl��i��l
� �L����ǎ��\F���Y5��!�1"E�+�������,�(J46��ɰ�_�޵�Ȥڏ�5��پ���f<L�����3�)�d���&�Vy�>PۛH��J��O�c��
(�*�P�z�#�Z��� 6�迤p��݁ze��(n�H� <��P�=M;{�jg%��Bbf�Ūֶ[���V�ߋ�;V���x����<�=��1�*Q��"5ÁL,I�S]�hi�ܘq*|B��e�]�ně�'[���ݼZV����h�iZ�����͋�=��\��x�9ι�s[�.%�b.9�J�w;�.�UUf������Jj��#l31��w�R=тzPAd���W\��e�>.C�5ώ����#����?��y�{�Gr]���b�x\Hi�ׁz�"!8h�Ɯ[�b(Uujr`h �Vd���g��j��s ]!�Yf�?�����JcƋ���0Y���Vy���;u��:�p!)j
yѻI
�6ھ�d�7�k\GWjs:�:f=�]Tkm<ė��� �W/^�.V��ƨ|������H�`|nN`�z��Wn��D�
NHj�2�Đ`Ӭ3� �$I��Z�y�a<g�ј�"�bx��eR6prp�!�H��>-kfƁ�ҸV?�Y?T~;���2wj���)s��6KW\XF��H�J)R1S��t�ڱ�pf��9���XUi��j�|H������3��Z��.��,v�V�s��a1FkD����]�Z{���1�~�;(+'ٶ�G�Z��˂�Z�Lڹ0�T�2$RD�,e��5vq�[�Z�smSN=˿F�c������ُ�����W@�����>�K�k����V��� 2أ��)b'"P}����.:=�m�B_��O'�Y<0�p�Q];���2��NkEڑ��X!�������.��E�2��l$zG7�)�σN]j�ٷ�������[+�[;Q����#�$�xM��;�c�Ӷ��I��,=>M�!Ne�f�,՚�n�Mʝ�a8k.�����t��.���;�)���I��r��q)���ڥ!qzS��[�y�J�<�I^2���B���-"0�);�%HDѸ8]��Gwْ�{�+���&�,qv�+ȍ֫_��cd���~�(\`�2�/>��y�@�ٯ���7�+�x, rX�[P��D?]�Җ{���+NÕٚ(��$����������7�xa; �'�Z�TL{��=M��)� ��ۤB ��4�?y[^�|2PY����37W?fX�a1�����z�G�ɦ�vK}�}��d�����(�9:;�ɡUy+ǯCC���(�t<���$��ҏ���)����/U`';u���O���L��Myt��p�Rm���L[\Z`o�e�o\Ӄ=���]�͹I�c������?�4M�ͭM��Q�Wƿ,e:L��J�\w7�C�t�"`'/o�-����<Wb�']uN8��sޮ�twY��e���Qz���dD\G*������s D*>4�&���el-5����>kÍ�R����'��#�Y�>"��6Q1M ށ�Zz�nh*�A�o u�
Ҵ0�my����L�7����ۈ�6}��D�+9@�����^�/��[(�"���(4;N\��%������DmNg!R)����[��Z����|�%���h�O+�F���d~��D�FX_=3 ��5`"Dm�����"�,c�ŦM(��3Ɂ$���8�'ڠA4�>Z������w�@	�%����?�J�Klb�<�E��\�ڝi��s��,��֖A���BmX�����)^6����B�A�lMח+QQ77����ة]��b�H-����w)����!|l�q�k�ӛ��dOc��X��n�~xU��3|7u������%��Ӷ}�A>���Z����6:�A�>���2d���<�� �Qm�<ئ�ё=>�;�zJT�S^G�����(�K;�k�38$���O7�Ղ�4�'-Q�������}f9�������G7�i^��~)�x�*�6��I͍���2C>��<��&lqP���kk�+�0��]#�
�#���܆o�u���Xm����ĕs�}/5]+e����pٱ?]�!򀳄7�{Ql�'�'�߻2�yb\���`�o�-�EI�M|��G[3(�4z�[���������͍�F�3:.j�;|� (ւ5�4M!��������7��d\A&�����kϐ�Y:Y�7i������7��7"�d����A"��*�°D�"��.<�g�5z� ѧ���<�����C[|���}�i��R1ùm�'���ˌ9՝�ۆnQe�4�_������t/��y�I����s#ެ.;KMP�I���i�DSGC�Zm��!Ҿ�g�a�!o��W=�ab��Dw��v�R(�{HF?+5��u�Z}ԁ֚����1�#0̄��rt�Imm�؆��:�{zx�8>����,B.Q��/��ٽ����D"� ��P�y�����v��p�<�U@#�=lu��۟��\i�>�R�TpBՆ��\P�1������$��>�T� 7�Պ�,2��:ZE���q>����vy�PSKhU.�]�=�?�S�U����$:��FjރgԿ��6�Լ���C��	rNY�I'>�Tb\�Z��[�񉨮ʅ2��Hyd~���I��,�^J7�Wb��rLȬ�D2T׵~���C������udL�x�kx	F����s�G��I&�l7��K�x�$�t��_��.�IItL����N!��J�Qz��	w@P�3�BJ���q�����"�1�atNE�����]�q>�į��qD!�k5�����&�P�\��B��1��kʯ�]J|��g+�����%{�}y�{�Ji��y\D�o���V�����?@0��2���*4�(T�Z$�j�G%<z�$/�%����	� T�I~��vB�p�����	@�mU�L��s�HI2�ƫ5y]?Z�VJ��<����K���ͩ�x���)�����rO�s0��J�5�����g-�_1��B��~�rB�) <��Y�Q�� ���M׵�2��~rƪ�i�Ę�^aO��]�+��ȏ)�XɃk�$̝	ó^Zy�)����1�����������r�;�s_'��u;`a/y��<�(�+�\L��LG��4l��0,Q���˰q�2���ƽ�ޕ3(c(���ؤ���=�_(��h'�r�rZP"��ovJ^0O��z���,޲w�lr��_	qj��*<C��]M++����oG���@0���l{d#������p*B'+|�0N��lR���B*B�,��F��έU����bH�JF"I�F�yӺg���}�`A�-�Q&%7�&yv<7i%��E��4� K��<�
����!=^>��e��9��J���C���` P	|x�V�}loت���+�[$!�z������o���+��?��'��ݗ���Pe��1B�	;K�����b�D|���� Ϭ� W��.ۦ�3�/[eݖ����R�/���;�=�/�3"^J��T�3*�P#�	�tK}�}��9��j�I�賿����o���I/a��8���+9�$F�a!�ۯ7�:G�u�qE�F������r��]ؿ�N�H��E��㵊��hm���c�/JY��%bQr[xã�b��>��
G��m^�:��X�#�sG������#�������if8�SF|B����Mk��q��pMz��<�3�Iq����(�~�P��������7�ȱ�F���ϓF�?�F���D���VFT��.���T3����l����&+{9_�`\㣶���`;.�hU�[ �w��0_/��T��&Z'��������@,�5�������p�L��q�M2Z�V>���5U��G��?���]P�^�q��D3����h����V��m�9��gXe�t9킧��ˏ����;�X�1��u#����2<q���mQ�������Et�l��"�*�+v���{/���A���I�%}yPfDG���%�y35$3��/�I�3J�);m�AĔ���-X�6z#���LV'�tGq#^[R���[U�{ż?��[zP*�T��,3F�H��K9�j�)Kɰ��R���n<����]���U4>:�STU^�	y9o��s2��$&���ܴjm^ڶ���1�����D`����o��(��͡����JC׮��#x��/G��Q���u���yV�x	=�����G�ޣ[�����&ft��E��KCj'F)��R�F�NNۢ2��`Fs)�'t	m��<E��������A��C�"��sj�vM��az�2�;_��}�]r�Up�|
de��1�F�X��d�����%Y���$�~% `���<� 	�l���̙���y	{�b�����J� � 6��������)��t��"l���C��	h�'	�ga�2�x�@)Ć}G���_b):���W���=O�X�#���cN8�X�7��ڈXV2d1:483�m��cED�K&8�2-T�@�����B"�@�A{(���n
��'�ʸ���K�ޫ�?HTߓZ�Pulsa����N��<%2��؊�������%ݖoTyJUf�bLP��t����F�)|�� z�O��K�������s�ք��p3��|�{{v|୷�	[��G�W��(���bh|��#ߠ8��0�� wHwr�H�a�tբ�r�`����s� � 6����@��)��t��.���I,OA����7�iU��NMy�^-�����]1��s`�ž��_���r��QJr���*It4-~��[����U��-�9H����yiQ���7?7����zB�4ǘ��[8v�����,�Hܳd�[Cn~��9� \��3�r0�Xo(P��g QI��5
&��k��g�ENL%
���|J"��l�'�!IM囟�8�[/�Cz�%6�Bpt/̘q���G�G�ilT����k������e���q�/�U f������
[j�%c�J]�9T�~��%8Tn��b�	�o�B�O^5�}iR@�T�"�����q���B��C�vt�CXQbWpq����������}�����W|9�NR(	`�4�P�eyGq8RS�8X�V�/8�)���B��s� �uG�l�sH��	n���(S�:�j���8�@T7��r>� ��b�݊��*T��m�HM�By"������·��HɽW;�c_X�k��g��m�x����C&�f�����2��:d��m̀(X��0�/ �s�J,���y��ihz�\�iT�F�yҍ&�r��i%�"�Ici7\��o	�m)U蔍o�`��G���j�1�k i��	�C+��W�����G_�98Fꄍc՘#o�:�iJ�F�%Kĺ�Jp>�\��Xω��gJ[�ﷲ@>��H��@�Ǟ�M	ҡ��WK i��IkȢ�����ݯ^�A���P�����&�a���㔅�?L S��xwA��@DA�ނ�YJ�1���l ka������K��ٗ#��Y#���:}�g�kDv.���y0��Gh2i�#q����7~��.�t��KqTу��ac���n�nR�(�_�nˋfF$�v��g�j�5'��[��\u�gM=��3ܑl�#S�U�@NѨ�f��Q�ɴ_�zj�9�Y��Mw�#��h��T>�Z��~7�x\M�:�[���taٽ��d^��G:1�)i[�B�d0�d���/HkN���l~������7b�0���g�q���?Ҥ����oM�r]��H-(V�Zz�l'W'��QPm��q�h���u-nG��B�+�RB�3X�����ت;.U�8�)��ً���^��Zl-辐	TF�џE6�f��{���0D��M��ٹ�蒜�Vb|�l;�1��O��`��M�/��� �ד��g��"����H�T�.�]3lA&�z9�3���q&��|ۦÄ��O�LCb�� �^J�8�W�uWE���c��Lq"���u��\L����ӝ��<�[9A|�>�Y�O|sf��͢㊂j3�I��SGi@稨�;��]�՟��Ѣ�S\���Â~�|䞃šTw�R���7 ��d,ʫ�\�+`=C���F��F��s(�vܫ����*�S�t�mh��9�dz�;�f�-�S�d؅J^��(����oq���|p�d(�2%E�|6�j�f�Zߔ�S�q�X���]�&z�U�jJ���Q�W�{ ;�ax8o���P������t���)eNh�E��f�b��Y�m��q<����H������Ⱥ�I�d��/t��=���oj$�ۏ��Xt�� ����@������E\�(~����Ӝ
=Zյ���wf*������q7>9�5�n!g���w=�LM���C��UYԌS�h������l�z�����L]xzh}�3p����v���j��2��@��`�ZCf?�+�A��QL�^pY�p,��N>"�}�
/�I\F�N,�+3��e��x݆�ܡ������dfh�{�nэ�'`Pu���k���]g=߾mO�a�17��>�Kz�Z�zp�M���w鑌��>�2�3Ͳ��v�9�?j_Ś����Њ]�^z<�/�S����R���~1PD�ɐ1�d��������4�I!L�#n���&֘��
����D��dQI��h��88A��Y� ��)�s��/r�r�Z��7o�8�:Zn%تhG�`��_�Z�E����������>j��>B����t�R)�z/�Cb���<)Sg��z��veQ��7��A)����Z#Ug���D.2���G��:7��X~��1�k���;6�|���gg�M�T�+�1ݘمC���W�2�o<	�i-@90q��ݛP>�����r ��-괢LR*B:Ǝ���|�yZY.�|^e	 �B��������*,��^z�8���@���?���vX%O�!� N�����){�^Z>o��:+%W�0��U��h�%4�S�/G�l���.yG��X�R�E%H�mO���,���J�p��2WH��d|gfϯ8�fy�C�Q��k@cp���W��eOa�TT�6�-�������������/���m|�LQ8K<5���x�ϫf�m|��t �PM˿z����'қ�bϪ��~茗Q�x��>�)�����,�ی[M����E4P	���kV4ax�*�=�d+�; ��Å�$;�=m�b�H2�R��:��'�#�O��|k�4�*4�� ���=xn r_g��w�sAZNH����޴�}��?�J?��Q?����B.�sy�ux�OtU�?�x��*�1��~���8���J1�v��=��R���ƏhАB[}o3�ܑ��A5TzhnZm��k��&�T"9�|n�-D3>7(\#V����/��HQQ��T�O�D[?���1p����øe�8m3|�K鰥�ԅrOU�	�m��m�=`��k�֐�+�᫼Yw�W{1CE����i-��>���S�Z�n�� �[��(��2���s��^�'MVެ���B{��T뾳�n4͠�CI���7�9��^�✎{�=`�!�SY�qjn¤m���S�[�����]�]څ(�$c��\ыL��H��Ь�d{�k��� ��Zb�8��&�N�V�|s�h
ԼۯG,�{I1!���<��Уb1�)��4T}��
�fm�C��
��}�����N�+n��/�,zlϣ��������!WW_Ց3Y��[X9�8>1���H����zIg�i�L�^����\��9s�ZmݩX�+����c�ux;�UT�͡J��EN~�P����Nzl�g�	�a�s���F�^�M�Y�4t�W��&dČ�]vn���C5��s����#��<�>&_���t0�:��+�6�=�zB�A��=*�u��\���9엻�L�͵��|���e�,M�������y�{��am0µ��˙0]��I&���5xfk����>	��-�1�	Hl��T�����cř��YfjÁ����E���l�oKz v�(�����d�[>�8ô~� 3�;w��+,�d��m_�?��	�>�ά)D�.�a��Dj��R?UO��9R%�A��+�G[r��1��X\�k:�ʹ���K4��	�v
�e%eZ?w�a7��O�~���'�p��N���HhR�7��L(ѓ�[t!��u�B7�QAo,��A�'��'��t��ȐA���p�3��/�L��%�cn*(��f�����^�`��|f�A�x�=����!�կ���4�	�ZHA�?Y��o^ˌ�'T�Ha�k(!�<�t
��-�w
�i7��j�`_�D|-łd�c���!�Ga�<!�Գ�\�����7T�Ήr�2����K"�P�C�6If-�i�yX�e�~~��Ż����ʼn��&�+հ!ެ��J��7�L����=����[����>)Ն���Ϫ���/��a}�?� ݵ�(��,�ެ;?D�P'�R|Y��Xb�F��3N�a� 0��&�m�u����!�#dI�~��N���Yc��6TZT�����i�z_$��J�L�QL�.^9"vNɧ�XU!;�/��ƴ�D��S�_�_�)D#Eq�P"���_�_�ڂ��"gR{�ξ݌k����yZ6�-U�9�6���M�`-�:���ex���?YhWom���ǸCw���f��GS�����9��Na*u|I��,Ili��U1H�U��,j�>�Ar����6�$4C�|_����G��,�)�<������n
��5o{$>;�e�{��{����I5��+-U��2�	2�����P.m�7D.{1L#�w1wq E[�]\��p�G�7���o�������G�Or���Q_�V]�T��O��.}��r�,���2a�� Xce�C�"܊�}U��c��1�K��f^���O7s,ȿ����$(����n��"���6���:�(M��݇��������Q�/U�=���F�tB):O3̚xR�ͅ��c�:3`kk$�ãj,���P�Q1��_ہ�7t�T�`��"�_󷯶�X�l0G�>�m���E��Zw�
�cu�!���::�����{�vC���A�3�+�/��V�����@�3�f�c�a;�陸���;�����25u$~��}.dT:�+5�5u��[���������-}\��PC%�]�O�S�|bl�ˍ�����Лt��ѽ9?ɎH��.PyPn#j����*Κa!��9x���}��1�%�#v��6��̍�q+�`pC:ʐT�&pi��9?%��S+]�W̓A�2����}MqwƆ7���wb�`lf���X{�'%9`�C�.�f���ҍ�ɩ������4UB��14���j���C@���mkd��1�����ܖ��.��ʎ�TL��!��aw�[L<v��t��M��E�����Lπ�H9R�~v"N��6 �7f_K��\ i91�Lx��v~�9��ؒizB��6<i���އ)��Ru� �
�E��C�EjKg����( ��AԔ&�||	/)Q��� ��k�e��9��Wkÿܕ��yYג
�4:��?3���k�[T+�mI6EO�ѱu:�kK_��;��|�Ť��i��1��n��1(��.G�����(�ʜ��A��W�9�7�K�iۢ*���>��0�Ԏ1��������X�@(�'Mj���:�Ϣ����߇F`����}ks���D1L�X�c'�� C¨�'�t��A);��E�HR�����GČ��? wsvu~��;9�;8[��mS�	����B�ye�������Bu�=���b�'#�YޮyiV�#�h [�P�"\�L\�8Լ�E �1� 	��/�SR�uh
���޼��)͜�����q;L����V2�~��|M���T��'C:x�5�j����)я�V��5}k�T<Y�����G�f$w�[1�J��5<�Z��A�>hR�<3����N6�ȨiԬ~�f�D�w�:/B�Vd����ͺ{�Z�W�~�oB��D���$&��UF�����`$',?*0�`֡�Vn�����g,��}����k�7+���DV�Y��1i	!,�3 �"�iyA��,�!�Q#��Ƚ�3t��<�����[V���W,�f�*������[ĀR3��1\d��Y�)-�oN�M`�P�Kw�/�|��)�w�*Xp�e��.��i>��v+G�	��S���P���t4-���l����`(9��0��YǎR��t�c�V�Z�ffl�7�#L1��s�@�Y�?�����U��4'�Y������O�%�ar��X�����U��)��n���uc�IM?S�g5�H��
�aUI�S Csg�LT^e[��E���Ѷ��yO�G�g�WU�&��[���n�$na:�ϥ��c��j�	��R�� �#yr���jg�*�<�?|��,˻��H͘�bkt	� �BJ	�<P���/�fX�/��-=�2�&����-u���GD�!�BȦ|�BL�+�Qы��\T�E���(��6�oªK��y�}��^a��U4K㴈V��f)t%
���2-�Ǭ��~Ǉ		��LX8@t�qER��h���"�������oH�m�����,<��{�u,nU��M_��4p�+tߕ�n�j���i6Jo�i����ŭZ>-�@؞���u�6o��rK뺍NJ��cs���}LsB���>��T ����uc
8ʈ=���E����U����fd�c[/g�D�h���/:β]��+7G�0��$�$�2;��f�9E����e�P����gx'|\X���� B�#y��솋uŽ���Q�KK�O�,)�k�n��2��Us�~��	=/�xɍR�-�g�0����t^��t����Ѳ�����	ќ��<ntIOx��
�1�xg�A�[9j<)�4ש��wƿr�_�e�c8�w���N��Q�[=��5��"���|��`?�jr��+g�HO�S�6�R#RC�i��W�9V����@�)�O	����QX
���=�]���qڞW���h3�'�ĭ�P:%Y�y>��5۴�Ăc��e��ί�4�I���K�@��ݷlI��n�E���lDC�ߝ�Y��"xZ�#tL3S]�`k�kL���cTC��\عOs��fU����a^�>�m0b�ef_��^i>b�b���{��Ľq��:���}�B$�h�(�ڈ��٥�N���]Ī��^ܢWO�B��Ma���� =FҤ-�������>O��	��{��9C�k����9/^�P�)��jaR�|m#]R#(�P~<;.��h�Z����&A!4�;ҷ0�Y�IW�z�*�aou�k)W#�|UzޟՉ�ز�H� ����~UP46'�0~�m���h�2���ۓ���n����?Y-=��z؄�VmOca/�C�6Hb�����r�1pQC��I���,�eDVp��ip䖧��@��O������rڨk;��i(uu*h]X�����;�񆒯���8 ��s2�,U>Z�&ߦ8���k%�Ù�o6Ω��9�qxȰ���KD�a��U�M������kG?U�/�*3m<l���+2�|�u3�A/NQ4�Nq4����q�P�*@����`}�q?ݦ��0����%X�]V����E��Al/֡'��P��̩��C�٣��O��Q��`B�c��.����`@���� Q	�
��/w�"��nt����&-�v����en���$�]��1��Ci`��v�r��r��^G=���_���/�hY�8��z���B��ٚ�S�yB��@�V�����$̓�G��Qj���s-g��tn����>�rx���L����Yۧ�S�n՚<���2� I��$���k�����]\b��EY��<A�9����T��?��O8� ����-�`C�@	j��E�2L���0f@�t���S�0�{�Ѻ;��YeC�f*.��I@��޻�}�
�J�����y�.��#��Hy�3e9�Eq������,��C{嚾�n�;�x�g�Ǿ����,�C����D"�!ojcH�����A
��� �n�����q���X%�P"��	��s�)ǐپS��7�]v�����,>.�$�脧��ĕ3޼DZ�9����L�ٮ�l֫���1���8���(�k�7�f=2�-�Pb)��܋CL�'�o���(C�9�8�G(ٌ@.�Ŝ���������0�������o,���q�
3W�i�ƨp`Z,�n|���x�a]�c�:L����x��έ[R�,�k3��#����`(�֏rEc2r6�PM6�W�)�g�%��f<�|vтc�'"t�b��0 �=v;�C�QӃԈZ�j T7Y uE�:t$�Ƌa[�B{[�p�$�֭v�$�U�Il���}�G=�$W	 ��	�>rDi:�,q@�!�eZᘧ����Խ��I]EZE	��W���������F���Z����2�z�)�qi�:ں\mPx*��$Ac��+����F_�ʬ�|��e�1$,'ى%U�	D� �)^�������o��Ҟ���1P'�g�u��	R�0�����㕪X1�8 ?�T�@�^3:C�O�3��x������� �q�W ��]�\,���d���������sA+ ��QB�|�����mN�̈i�?֪�˹;�󧥺#
�y[u����qt���H��f;+!r�F"?� �'�����gţ7[S�z%��~�1 �F�P+�s]�1ֳI�p��M5�N�`�^�r0�����{���0I�r�fӽfc��#�|AvQ���S{�c12� �0�K��F�
{N��-�C@mD�+/L����&��g7@_����A[<I���ʓ�B���:��p��C)�!#=�Ο���;����q�x+_��~��Fh���`��4�S�qOI��\��#OA�;ϝg|�}�P@���5r\e�pD{�T�6�߰0�6|�sjg���M��n��i_W��@2�wO�:P3Bb����� �ä8���0�����_-�o
eq`����qy�ZnG��`5ds���/��yor��$`\�^ 1���4R�����2�d�v�hӐ`i�}��\+�M�/Zda�o�ES3.�*��LR��A.%;�T8��o} lv�mz�:�I~����+o�A)٫���.��?�9=��>x��'�ŶXd��b�O��M.���]^�bv�"�t�>S{��,���D�9�h��m�1J>�0���Op�Ҝ����R�CyWl�6�-��M̞��1e�u[�N��!`��� �*4���ԉk�Iۭ�w�h�Y�1n��~0�{@��=������7 =A�{m��Ba�i��yc���[
;,U7:lDcqP6v�Q��f�a^#��,U�J5��}Xe'�i��cDez�O\�^-9i��N�9ѱ��p�Z�,�\��gepT!SU/!>b���Uh|}X�A���/x0��{���v�X� �S:�:�������cn��_��m�B�зs5K��H:����0@6Ks������Os����'���g�~���f�1s����غ�٦d�����g�-O?�8�#<����ƿ��Y�k9@_����U��Tm쫬r����$�Z�\ ��Nt�;�n��S�=�̤x_���w���ʺ�`y�RO�}xI"4��>x�c�!aUG�X�e��LB��a'�hp_�Z�I#���_�t��"��i��p�ΣC,��S�2Ȟ��}'ٿ���}#��@=PH�OC�����@ݗ�W��<�§[���1�*�Ĳ��%��a?�_u|YpX���l�f2ɜ�лa�U��' g�b<�� rAݠY҂N�8�^j���c<H�Ϋ��~#��9o�J��a�CW!���F�Q��p�k�5����Ԭ�^:��˕g9�a�D�̜�	q2m�i�)1v䳚�k@������;�w���^ΧkJ�����&��=�G�P�Y�ۯ����#2�{e�W�oθz|�y�Qb2��0��t`�ܪ��v,����w!��6�\]עL�1�i@ٳ»��
��?��|w[���q?�
�
k���\-�%J���f_��Mf�������j���le �h�&��������o�a��[Sg���a�6���S)a��Ǣb��,}�-P�m�/fǹ����!�����_�����1�����f�8���k����M{��5	>��:�r���B���(ҙj���J��5�3%��̜�Rc�Y�QE��Z$;��O�����8�=�+*b��i��lћݫ()2z��s�h�:�Q�oi�Dm�r~��G�� ,��g���UB@�B��yI�Lc6~�?��#��9kăǅ�����M��=�����KR3���#ї
�aL_2)��_4a�B#A�Yq�~�"�}*���"�����J͚G���r�O;�aVqJ��}n E�ˎ��
-��WTQH~>	ܑ���[����Xn�[BI���B�.��G��$x�����<C�Kw�J��}N�ʕ0C_����K_�N���� D����K�[t��fM����>�����ˬtm����n=oLD�r�`�� |����&ۭ�֛��pRX�VԖ[_��,����%j 9*���o��>�aq贐h�;]
o�n9=Y0׷Z��,]���Đ��B��$�m�s�N�)꡾@�@�nZÉ��%O�g���	�0m��4D�=�0�K��Ф}9�����2�������Z�pM ���,g�1uB�R��iR�y�"��(~¨̔�Z����S�L�R�{�w��!���P9��V�2�~�?N(��~F�>��RX�F��N�p2�"SW��9'�&�AN~F�k�3Qj�:���y�B�pn��������*���+�:]an��ѷ?� ��%�Y�x]����*9��8�X�qbt�#M_�o�E�}6D�Z4[@�������,Nٸ�d���@��F���C0Qb1��р"q������4�e��عV���eRY���5��	����^��1(zU�ܕe���[��V���Y��H�,Q|2���.�fUS��]z���Y�M�'T�����K#���ȱ�-���~�o��M�^?��y���*�м�
WD#R�vj4�)-A!�4��݌�pB);l�`�k�/>��< +��#�&�t�����A�ˮy��	���4b.�n�1��F���[U�%ͣ;` $��o��EbQ��(��t���;=ܖ�������L�Rp@J,��4T7�-ݙ�wQ�*���J%����D�Y���0=�0^����K���)�#�AA�Z �ʟk��M>e�P�4�_���m�;ͥPXp�!V�7���F�kiQ��V�Tޓ]�x�����:�K�
4Q��aZ���[�NayJ�xH�?׀=<Q��.��A���5ص�OR*M��[x1�����F,YH�#:N�����Fy�j$��Cw��_��Ci��&廓���lTZ\�b�l.�Ih�Vo�/�����l�$U�3ֶJ��o0z��|���@�}j���v��8|c�'|M�Pm�v�[Κjx8��Ӂ���ƾ��ng�W��\p�z\zܡ��N�%#L-��Gى�y����&h8mg�v���������zq�L�%�~��]�i&�����(A�u����![eWV�k⦆Z�GW���xu�W��G�#���L���:Kݞ�6 �a�i`_
�ұ��D�՛����҅�?�]��tja�
X�̿0X�1�^��F�^�����c(���u�;T��%9���ZӖȦyZ��U���L��.���)��UK"|}��\���T��{G[�%��D���F��rj��x��J��yvD��ll��#������h�Ԓ�G_+W�l8��~o�A�}���Y�G~��l�8�h.��B�RݧL)��z-�eB`��$�{��'3~�dUV0T���%��෿"PJ)hw�T�0��Uw_�o����<�3K��,%���ٖ�v�� 	����&�͏j�S��l�bȗH<����b� ��C����B<(&��>�;�@���s?����QYB�kB�~)��j�"�MB��t�����F��8E`ӓ���%sH�$T��6[���s���Oǥ����B����P��?�w7�܆������ߊxYa:���D�78=q���c�Ek~t��;c�t�r�M�=�E�~ ��W� H��"�JQ&��_��bop�Dl���K�{W��Q̴�<.='��D��`/_�)�Q	G܃B�}yзո+��a}��rۈƕ��]���T\�Z��2f�M6��8�o��1[�}��A��IeZbŌS�|��.T2x�S ��[8�Su0�ɪ���,�B~y��۹7��E#U$2�;SD�C�q���5�%oXG�{�=�J�P�_�EE�Ha9aG�̃�o��IQ��/��k���sK*Tj�F Hl�y�
����ޜc?SA9��S�[5y8чL�g�6�ؚW�(Mݴ4O�N�/��� �k5%*�Ͱ>͢���+���1�P=�U��M$�cH��%�~z�v���	�v�� �a��3�=㤫����VD�c����C���}D�N�j�	�3�y�6t�)3�¹��_|�&���/�����	�[ȶ|mQh�$�~�������o���k�N��J=�dpvY����0/:l�� �UW/���[:j�C g/mə=�`��X�c���k���s���ן�Tޅ�v"���
 zU.E�kq�0Y,�Rg��k�¿b��s�E�5X��L:��B�"���=�z��ϟ������,���_���H �9��t�KQ�O���i���]u�#l|�R��-���ʜi9�i�Y7��	����~V�k�/iG,�*�sB-���`�/�Y�A:�;E
(
[�?3���e�(��RҪ����	Uۀ�p3��w������~�p�=��h��Ç�����,�g���	a�QΏ�Y�M�W��;���Vi��G���sĿ$����%�D���3�Dnl�w9Ȫ�v�8�MH0V7o��������25�	��n��ml�:ܐr	�����x6.��'��k��=.YN������[�	������M���?��z�%����TKn����1��+��^�M�>�%(���]H�~|�C���d���b]�"c~0�n��5���R��_Uqc�b`s)O�陣�G��/m%0�Hja�a8���P��5����\Ub
�=�/�qs]A��������x�{دdP$�j�Àa�r����b*���:�i�����MH��嗚��W=�K�'E���ȉ�qz�f��wNv�~\G��S}a�o���d��gg�e�%# 6��)_���*�/��P���gAS�ֆD�/��� Mt�M۹�&��*Ɯ���X��+ְ0�P`>ׂ�O�����p�U�ށo�^�"ʹց?��P4hZ:$��Y���B�d��K-�奨CR��[�`dk��3$ƞх���a��]:����ټҠ�@��!��$�Ҧr�R͎XW�T��N���7	�B�D��^�h�A�L��vW�F�9�K�i�%{��ڭ�M����hoB轁�5ʲ�v�X�^�[X�S(K�)�K�b�h�<�QW���Дt�t�����t�tLE���l���]:�S�(s�{�)��0E�)��n��_H|д ���h[Ajyv�=���q�<ܟG�[
]vI�&�1A�e�:�"�p��a��*�~$�b�N���1��>(68C:�x�����i׺�m�'���zM����n%|����l0���v/R��?�l/��'o�%m���f�Yd�F;�z��sA��*�c�Ń|���#�m
���Ztp���%D�-gm��� {$��A��$P*�z��c �p�=�ΦeT��7o�a�����=�|�7�Ŷ�4P~|��}y݁����%b���ݴ�TD����6�,F����ڼ?m�h�1�R^�����a�}�#�ʣs�g��X/z�r����r#�j~[�����!_W�Ϲ�#({w*v9���CǢ�u��MqK�����z�`ӿ�<֒��Z!�Y7Ǭz�}����sU,g�FzcZ��1eB$�+p�C@��q�"9��cg��J6Gb�%�a�dʪ�v �k
m�8}��_Y�G�Ni��f+�J��s�����۔ %����_���	�e�v3$۸hM��nu����~9��砋d͓f��x�7�����j����}r2!x�9��&vӥur�h���xe�YkH�ʯ�r��X !��%�����4�8-�P����̛�Y�]խZ�6�	/1.�9y�^�p�֭ۄњ�,b�����̈́a���9�&�&��U�z5�j�]V
A��:S5np��Ck�/3f͉�����oߨ��$��W�)�A�)ﴽ�9�r�:�h�bļ��������M�%ɾ\��{�վ3I?@y�A?Fl�`ѝ<�V�U��G���h���>���\M������ukU�xN�v���ȱ��Q����e�]�	�i��2C>L!����d��^�$.|.ݖ��(ޒZ���r����c���|���l�1!�(�S߀��5�Ai�Ϻ�:P���n`/��U�+�f��+#�JJٶv�Ia�����&Up�W���W�������@���B$�ޱ�Taey�L)ٹ�\�iX��#��b��6T�҆/�Ʀ��p�'6YM��6:��:�`�/S�Ǿ�{��%��0��ku�%,(o?:ݰ�L�(Zxb��E���8�h.)ӳY��^��ѕx� u�~�nW��ɢ��������K
qPܥ��fG]^�r`뫺v}���W�C��>�H��7C?%�x�@A�֥���t,Dw���ψ�><��ή�D�:I�YN�B�ꦵ|L {�-�9��D
W'7�!#�A������!�8V���	� be��l�k��ZD)/w��	�m2c{|+��1X:t�s	j�8g��^��o���Ul�{Ɂƫך}��Hl�v�����b�eō���lrURM��b��~������]�%h(Xv�-�?Q��KC�$��i8��iy���J�1gx!��5c��N�]������W�CvŊx6�?���a��	Zس�r/����9��/��q��!���Q���E�N&2=�^��#��Ʃ1��)?t�a
	���S!�B4�ϹP�f��τ��e�����r��z�jЇ0)�]^��ItuRٿCh��[�E3^���������n��Ɓ���ԺDH-������r����i���� յ�'�;���Ƨ�D��������t���>�nu�K-d�$M��&�P�p��rY:4�%f~ۂ%��)�^ ��XNfp�C1n�45��lQ,w���A��5����b½Hw,9��q3^��7I��U�T���nnz���� �@��e�E���+���_���**�H(�g���K����UG>ҍ!At��+Z�1��5']�q�UYd?���I��^�X�Mecc`Y�HQ�|�V�O�
e��
/�,ǷA@E;��١�(�顿�t�bcI�wB�����Z�	���������A\CB�~������5�%�e���������Z3���϶E1&�5c����.8
�f��#�9��z���2�\�lQٚJ�S�ݨjw���
~u�\�6e����w/>�����tsNx�����FJ�Ͼ����V[ʏ���R�1�2��c��yS6���)��}ݥ�Įq��IX�/��������>w#�c��=Ӑf!�m6ِoc�|�
���AgPɵO��*��⿑���8�"�9ķ��[>6ʅ�ż�}�AV.���_Ph��9`���Ov�2ӫ��!�L�&_��R�X�$�/��)!��}�^)��f罒����Ĝ�(q�b`��Ƣ	 �IO_�U����!<y:��y+>3�e
 o����)� k~� ��0��z���S��kL9����
@��������I�lK����͠��������&W7l����=� h���Y��]���dqm����́���V>��^�C�P�Ù���hlLe��G��Chm|��1Γem���xh��)�P����_~�&���V*�!,E$3�jû��_�C�=s����ֽ;��=��
�����	�=��5����C��!�_¤N�ٚ������]��!6�ȯz�:�B��Ĺrh�f��m�=x>k�z՗0�2iX���f�6F�n�O�9�!��⛞p
�$G�,�hUb�͆��|٥�J��C�6R����1�X���@�f�n[�P��h�ѕ�qo]&ijWg��ŭi��-���P��<�kv�0M�n�L��C�V�0!ӳi6a���u�)��U�Өd ��NZ7o� "�^>rA#��V��,��傘E=���4�U%Y$����2&���MA�Ǝ��u��/w��v�U��?X�$���T�FC"+.����.�vR�����hg18��=��@D��G,m3��W賥�.!!zL�E}�A	Q,��*BUs��ǅ�q7�+�4�p��ّ��.0�������Vްf��_����A��,�,���'v��X��G0�f!腂G��������0���C�y�z�=#�)�Q��h�-t-L'��j)����!��U��a<x��)����/!D����XW���&�K�wε�փ�=�(���8��-�E>w���t��WK��Q�e�jѢk�6�E�R����
|�*S�NțO��@@�w]w���B�t�l2j���vr�04�I���<����*f���װ���cj/܂�\����[�N�=��=cV��"f�s �a��ϸI1�v}0H�|H�%�if@�]aq2Њ�q�.�����^n�"N6d>��qع kvF�����C��wu|���
�Ɓqž�AU�F83d�e7�H\��[��V�`"�K0��O@w��gp�� O�R����ń�+A�){�-f�t�;sžƴnТ���{�G�b��T����E���ƌ7=Ce
OG���+7��yk=��aO/���.Ua��&5����Q���5¡�	���X$�r��j��h�Q��_��p�7�����Gq�ӂ�b��i�k�λ�������P���O���t�E��UO׮�5)����$7"}fz�P?�취���VI��Z�c����9�!�.�Z*i%]�u�[��=�P�*D��?�^ٌYe%fue�"p�x��������_�*��\[Cb�����<�)��,i�2H�A��I<���k���Yܠ�\Q�4:�JX�J�{ɗ��YP���v�H�}����	�^sz	��R
�=��i8�#A|�o�[lxt?��+��>2m|�u��G̕}�D�j$8��Gl���	W=�J�'�G�bͿ������欄�Z�B�+*�|m����g�(���RY�Q��· `e�F�!��zc�à��7JS+���7ڵ�U�#[+lE��LĦ�=\8ԟ�7��YP̓�+Y ��@A�NÑ�N8=H�;-}~���O�֙` ���Mĵ�e�&b�
n�R�z����Bm	_�����1�#����͓�O���Qtn�05�a֜�� ���x�]���!ѱ�[$�y�̦դ����e�J�{��ᝋ��[T�f
�6�*�[��r&������v�x��=��_���|�����q}.�Yf�q�1s��>}#���#��V�Y���-��?�{�s����':Ei����$4���t&�������&�^�M���aqg�W6����-����r�A�_Fv��"��
F]:�X�xd���������Ԏ%5������)9�OՎ6�c�f���=��������}(�k�b�����o�����ѡ�_���ȏ�%�Y� Q���r�Jڷ)r���H>�ї�����GIV�~u�>
�L�"�E�U��F���
QY�ƾf�ARЈ��Ǵ9w&�L��)�.�6���{0���H�rqz ��CBv�l��9CLt��;&�b8mMw��ȯZ���r�8sGޤ_9$�[Ζm� m�̥S���C��ߌ�� 1�[ ��6W���5x���aFa��Ⴤ5����r줯ޯ�*Ρ�g�V���}X�]!
s_��@� ='II�<(:��ݢ1���FT�Cb#C�� }�R�y��^�ќw��� ����T��}��l1�Jm�,�D*��c;�:�u蟣ͷ����(����r5�x��d�|I,�Z����<
���t�Q��p�Qɫ ��1�xĐ�; ��~�RTZ�+@x��\�rd3칵X��s {l���M0�0��g��@[�E���|�?�tW����$!X���ݜw@O�>aԀ��p��eV��Y�󝙌Kb�h�����h��4-k���dv��>}^>����|.s4F����sc[ܜ�A�|Ad�ak���� �Aɵ��$��a������Ҋ�jc"q�G�TY�p�����l$*�����@�B@H�p��!�V7b�����-��W��"�s�2䂔��us�k��~�*$��&�nڀ�n�8e�"@\�⻖�چ�\�����D�ACDV�{�������k�u�Ʒ0V��	�N���GagP���#�ah�AJ���4��	�|�и�X��?1�z�nə���U ���ᖾ�x�a��u��2r���%(����5|tb۩##{��Pyz�����&}��� ��Q�p����S��zn�;~C��z�'{2|%�1��p��]���3/t���Jh�p�c�����1�/@���|��^#_��c>�|�ڀO�#a��[���-���&�#�*`��C�[���2�~����F��O�"�0B�Uq�v\��@�m��Ψ��G��Y�d�ӎm�#jd��G��󢪙娹a֞�r�C!$�H����O��·����=������PI������5uIC�7{#j@H����d.�
�9���MRqCx6�%�uu����;5�mr0���b��2`0�� u/Y�^/����B�ͫ�Vh����&�J��
&٧�o��g^?Y����kg����7S:U\p��������Q^����[j��x.�ܡ^ܓDp�h<m����S!��YS���VQ��V��y�&�^�֙�+U7�.���9dYa�/%�P���Y�����:������퀃-.��:i#�<bA'�y��LyD/I����l��@��}lK4]LVF���A%�)�a6��,���2~Z�A���u|�ku~�ԋ63�\������*m��Z�~r�F����E�̓zh��1�:���O���җ����ǅ#J�:qu��k}H�9s[צI	�RKE�[6�iW��X�[�����W%�����mqhA5fQ+��oK��cH�OwlA h30��9)r#�����ӟrQ�B	]	�>����1&�*Y`��q��7��a����g�3�@:~�FY'>H�}�f�������$��՞��J6��K��+����W_�ΦY.^?Ҁ�=��S�*�
�ڦa:a G:�&Vg�w*�x\H��ۜ����|���xS�1�H��yj�:�	�8��h\�U*$3*�����.A�g!�M�#"=�;�ox����Ծ���i���JwH��6="ӫY3R~V+d,
aY|xS8��k��_+!?u*���n�V�,F��%���jd��j��'�I��-Y�V,x�!ù�"IOtP������-�����S���453���O��jf/�n��˒�@l��6�l�"ĄhR���B\y7��%������f�����i̺+ ���^E�[幦�R��w�Tb2�7G�P�ɨ?��f��)����5�Se��f�r�6�fk�v3�It�B��N����?�y��Z>sƹu�_V!h{����BЏ�(fP2+��;���Aq��X��V����ԯ�����g��|<0D�u��m�;B�f�s�!28,��>��;-�%�䑷�釢�v:���i���?�%��"7'���y�8�˽s�����/�UJ�����C�A�y�Z������0@"z"|u�R��"<�~�9��+��z�-�S�e�	4*W>��^��&V���� .h�Mg#6�����}�u��**����)f�f���Q��� /�#P�����{���f0��*nj����Q��N(A%��
�['�\��#��ϕ�M�B�|v�/���HZ�zr�X��{K�K��)R�9�9���'���5��ٻv/�#��mesc�<�\SN^�"sP��9�l�;[U�;!�AD��j�c����XdJ�+c�?`����h��޼G,BY�2a���E_*�f�0���ee��#Wmk�_����$7��м]IN8��.{�d��DAd�yB�4×[7���ƞT�srȢ���{���6&���)�*�l���)���a����hͶ	�Tq�1ܱe8�\��6���s�0��V�BJ�<�o��<õ�{�c��4A��+$�U�͞r�,��XL���@1NZ7�:�*�5e�&�R$X/��5�U�q�()!0��o*���S;aӮm��q7��fvO�5�������ٹ�~������� �>_��h���D��:%y��N;���-:VX������Z�@F�_�S��p��[��߳S��8z�����.�ۮa��q7��AK���6��~�Icl��{R��[�ƾ�}�x��`jҳ��޼ۄ+��`~�0UY�9c	.F��>��Y-_쫞�\f�X���ÿQ� >7��S�J��[L�z[Z�Kh
أ
��~���cT���4�Y
[#�R?/��MQw�}j!�i�+��{�s�rJ�s>�ǔ盬X�I�! ߅49��Ѯ�I�����(f�����鴈W�4S5�ע|{w�O����{�Q���AK�J�ƴ"F��F���}}��R�{l����mD:]�005Z��6�_nq�G"-1����:[.�ݷ���T!�N�F�������ne�r�����,qũ^�3U�Ja8[�G��ie�z5�O���E�G��~�>k��^���ڊ�	U��(�N�&J:'_6Э����a]-��DW���d�I!��:���5b�J��<��7���r��&��o�#Vn�a�+��I�	��m$������AK߷���:�2���pHD3	op��k{�d$���8p���o`����0Hm���f�H�r>�YS�2��4C��|�����{9���qF���8�̾l
��#�م���|hp��Z��*!�=̹)�z.)�x�S�����Η�����G��B�`L]���t�$B�<�_�ǔ�Dq�N�Q?�K�m�T��;�P��!.�}��p]���85�e�U�J�+7�B�m�e��!����s����YS�Uw�֫f���[l�(�9L��W�`?��f����85D2|�aMEQ�*��d��	9ዠ�h��B�<��п��짼f��5za���>��Oa��y.������?Jԙ��?��$�q�nZfx�>����i�nfBKH�w��H�A�y�S\A���_�qLL����,ԑ���3����P��J�@)
�����4��R�=�e�(OM�+���/s�hLY���6��_�s7�J-<��=���
'�H���X��aE/Z�-N	߸�QL�P����11��� ﷇ�"=CyÐ���J֥n�[��˞���m$a�o����v���zĸL��i'ʣ��P��:^��)�4�T�e��긳�}]<�j��R���8�d~�����L]�D�gn#��P�-P�8��g�+��\�@�S�ZBMf�ڐ�1!0���1��8����\r`�h8������)��-tQQ�=�uz���WzM�f�#�}HL���(.�R��8�u�oխ�LW��0��Y��4��D�W���{j^�d�	ϒ�ڮP �\e�'�oIT��7X*�.��G'��,�4����N��p�,a@���{J�,W~����4�9%�O�]q�qQ�`J����%&�L�.4P�K� �TQ[ƿy�e�A�*��I??�o�Ê���N2z�K�-DN[���F��[\��bS�L�[��ϯ�1���U�65H4������&WGE�e^ɟ�f�����p��E������$�a�1�A�=��91������� ��Dohq����.�~�f�����q��>͋^���c�TA�u�i�|v��3�i�b�x�I���U%U��X�����c�R`�D-��ɖl}�;,��N0�kk|�M���y�X
P	`2Y�*jk�*������:���v��w٪Mnf'���E�!�jq�C����e����R�iFS�P������MǢ�:��W�p��V�X�:'���x�ٌ�P���جW�#8=��LZ�a��kU��ʍb^���	K#H6�ԓ35�$�%�I��^�RU ̧���ϝ!`ژr�5��H��1�ū�*&�H�؊�*�׷�0x!I��y1rPi�wAX��<����jW���]_�s��l�Z��X�s��Ё��M��!�,q�����dC	T��������0a<�F����
~ӏW$K��K,9��[OZ������^���~E�-���c���=���o�Z�� �K�s�f��1@� �,X��[k�}�A���Z�GMg�ID�_P�C ��U�"*�mQ����y΢]q��Ô���Uݤv�kd�,{��}�v\��DN��f�W���Ѽ5�P1a%uj϶�q�h��!_��)��PK�� ��`|r_��ފ���|U��]Yٕp>���ُp�ۗuݩ�3w�#G�j��5\���"�i�D-!��\7�������,�Mo}�F��tl�T�E�<ğ<��S��A�M���oР�fZ�Pv�-&�zaO�w�0�6����i�#&� �T�ї^?9��h��L&�5����1���4��m�b���!Ƨ
k�P��9�D��=��<9\��� 3��Ub�}?�xX�
��|�����H��0�g�ǵ?a16��7�.������<W}!�]�p����x���I��� م�A���n�B�,wA��p{���� &&KZ�1�Ξu�q U�A��m���P~��I��._rh��0
}�I�t��s����b=�������c�"�LhP������]�̬��::�;��Г�Q�+��'��c���p"/� ��@7d�F�_l�Zb��%K|O�b"coQg/S	>�AFQ�i��b;���s]R_(���0�(]�2�������	q7����h���z
β0�ܓ3�M�Ѥf ��պ�e��+s�+�%��ʐ:9t)�y�
���k�*�J.�������g��U����b4�{�4=�!�^�X�ՌI]��%r1j��/,<��UO�9�f+o��^����JA�Q�y|�)*��4��Di�)�U#���d�]��+_���Q�Ĵ�~P�|���.�C/�߭�?9���q���g�1Fm&��r:w��J#�"��6(��t�	�'=��1�D��X���J&�o���C���\�k���K���Y:W؟���66�ž��P��/wv$1����w\T&��iZ�6�.�%�yz��B��<*P w������I���= )�:����C�6S�5�����"��s_�:iB�F�Ȼ�𻹌Z�7�=c4�� �\��ym؊Le��k�C���Q�ظ@wDT����~���g��>2��lh蜟e�Ő�}g���k�D���W;72=��q�Q�Fh1t�0kTO�>�@�i\E�9��Qᑏ�ȹ^�B��yA��a(�Yb8����2�;���x��כ�V��p���Y���Ҧ�j�8�)���}"w�����FZopG`@��	p��d��Hi�|���8��y:AZ{Y�3��EA�H7�T�%�s����y��������'�G�}	��p0���>e��49�E���L�op9�o����a�M�'K��\%�[�J">T8O�b9�W���XM�n{�V[@G�����(b����ĒV����f��C��\���������r�u�%f��M�@	�D����j�h���7U==I�uCa��v��,�/�5c���Tf�_����k^*��Mj�\KH�{_xT��
�/�T�Z �2湉�M�s�>e�<m�u ����o�X�C��5Bz[�Ǯ�
��O~mV��R/��9��J/��Y��<^޻����i�r�@_���y3yT��0+>���9�TL�gI��"�۝4�U-�f��<~My�*+�zl�QZkuQB��s���-�ZD�&3��%Ah�����/�=Zx�A��mW�XG�qZ�kl��|�������k#�A�K��*;�Q>B���HЎ��5`IM�0�bӨ�e��5����V�Y�K�p'1�ҥt�Z��7/D��\���'0��$f��"��}�F��P��:��|�H����t�o4����?�lE ɒ;xO_�b�K�P^����	r�) �� R�F���x'�/R;�DA�A���P�E ,#1��E	^��3*]�uw�q6�H3(�����2K�t��ogG�F��'��/
RR�E����%<��Y�B��ݏ�
ʸ�6�X�>��?�j/^��pCְ"�,��_�h�#e�ڗK;Tr��Gjr���(s�>F���{I$�����_�#�tr�x��L��,������^�t�LhR�9����>������z�i]�bZ�����i¿�s0��o(�)��DL���ٸ��.���'f}G͹ӿ�p���>��Sr�1�\!C��8��Gi�:��W�$wM(�m�����Ҥ�_R��F _�kQ��ŃObeMq�{݆��^���Ǿ��oI�<���N2ӼO40��*��v��	�,h�|+?��=�f��Ts@�a�1�N��n�*�S���ּ�H���Jc���D\XK�.1,Qc3+�^��w��TB��F�[�vkev����N���[;��4bH��x|w�-�n^�i�cp�k4V�Fc.�n����J�B�4�J�k� �BBh�
��:�X0�\5L��g���IZd�@Er��]�N<<�a����ʱ��6����_ۄD�A	!jB��X����@��T����̸&$�y7R��R�\���o����Y���[�UV�M�XT\g#g���D�<E�'4���V����é���±:�8�EO��K��?}.��G`�L�1�T����¤=ǅ�y��[�9r3�n�%�
E���pހM�g�Β¬�
�*��� ������i�0�,M�f�+dj����4"�'3��U0#��A�k��V��AL@�$�N��%�J�I�3���bL<$WJ�j]Ď��-������[�:�u���_�*M��`��2,�����J�񗑩�Z�2=s;��/��VEu��7�!���V(��2S��Mc澭2�.����Bul��\�^	���\��P�jŉN���xIMI�����sF�������׷��yH|��9$
�C	X�@���.Y��O!��Z�_��ՕI�Q`�;)�2$z�K�Q�NR�����}��~�|�|�<��z�	�����J�(�u�����Ф2\��$�K�ǊA�ܱ+*'���4��pYx�m��F��j` h�������9�c�� �&Q����Ɠ�[�֖w{�*�� ��#����a)��|҆U��V�F⭢��Th�ݲ�3�2��b���'��YJ	<�G	ɏ�V�(�*�ƽh<�;Ӳ�����YU�_�FW�`��
���80�i�O�����Pw���jV̱�	�T^��K�E��4l��w:R�w�Fa�7$��K7ՒE�.��l) QJ7Tx�G�R
W��rqG�7�/>�{��ⓔ�K`��fw=M�#�:� $A�k]��=���_pqm�q�x*���N��A��х#DL��nإ @���U�ՋF򺀶��}:�4T4�����L�Q)�l#!RA����0[���0+�'}�
$�||�P�a��r杪] �v�C���;)n�`2��2�_��n�j'�JB���$��ϣC���.��JZп�W���*���,�|,~�w����Q�ꄦ��B�ї��>6<�������g��C-I�ɉ^�Pᱫ�[������`�{�!x��5�{���f=|sh�C���c�bȘ��^<Y��E�jk��[�~��������l�2�lQ��� �ў�j�;��op 2�W�kِ�Ì0z����$},�K�/(��a3�Ay��tN�1���
�jJ��1V��f�:��D��y�#��h�?��M��+���6pXw�ڽ�����F�ORN7J��e8d���ՔN���>G�3	M;j1�<x�K����"!�NY®��4·S�x͵�0����
�����o�ٛn��-�5����p�_����!V����Z��8�������}��[�Hp_l�Jm��A���x�@ N;/c�;wf,	U���No��#��je��ޞd�Cy�7�F�ys�δ;����G�poZL�8j�ƶ�TP��4��9ѵ�̉T�G�]J���������NaQS�L��� x��H�O8V&rI��В��d�<�-�(���Dq�3��1��ݷ�DA�Π;L0�J%���(�<w{s *�ލ�F�j�e~�0m�� E��VbI�c
����;�ε�6�*S�NX��}hPC����x�r"*I�]s �VG|	dӍ���I�K2�=��i}�U�_����$�6s�\@Os
8�4��=	q��?9��h��HU��B�!r�&��������݇��ް�2�`�G���H	�8�G'��&�$Tj3Z��")���!ٵųYFWRǽP�q����:�Fq)~���>������+"J: #1T��G#J�^Q��$��b߃�:�}�mk���Yʳ]�'���]M?P��<$;/#�T��o"�WB��7��}��`�ψR�Z�#BN,��������3�v�(L�c��?}ڡ3�x��*!�Ej�	@��3,�5�p
��`L4.6��e�}����O��9��s��@s�7Y�
h�]� �ݬ����P�$��nKO��oX^`�|
��lYU����%�� �S5�?K:������_��?8&3!I���n*�d��;�b��m=o��!6}PL��0ݩ� �8�_7叡kڳ�_�р�G���ܯh͎�xM'�IсV���p�<'��g�y��{��U=�a���mJ�e�6��(���%��U���0�O��hv�%y�ܳo>�k����t�] ��*���Y���_9&a��|o��z�I�OZ�H�ǿu���Q�HR8A)��UV�l�MGӶJ ē٦|�m�ð�������Y^�@m�RYZ]n'LA�<��Q�S��an.���Z�{C<%E�P/V�d'Ŭ��O�P�ϡ�[)�"n��ty�|Ӎ�g[�ԄXv�5tpK?Q'��㞪;����˨�S�dY�[�������޵XU�� ������O�8���8Ig�GϦd�gE9�F�&�^��*a[���yBrP��R�s�|�w�����#4���������r��&��ﻡա��3%�s&s��OM+��|�A��&^k�Q{�Oa�a�g�+�/<�2"�=pjk3^�[��yF9NM�p�L�&�ׅ���S��;�H[(���ő���NX�Y�B%(һr �SH�9e��[Ē. E B���^��Ȋ��1��m䱰��+^�TjY�L�g'O����	������DĞ�?h?`�z��%���qCO���<;�Dh�~
+)�pC}pN�#�L��_�/B?MSYG��Mx�H4g��ʯ�&����dw��q�B�"��oL~���n�H!��٭���	�R�o��<Ȝm�^}.�f���� rJ�p����Eq�E��:` ��eu�&��k{�g��T����V h�]�p�����{��R�[�B��y�3�F~�ZV_��c8��Ȭ�݉{ɾ�Yu[h�xFG�?|b�����q�Ou��V�Q/yYف���&����ܮ^-�V.���+���Ok�`�IM�݈'Yڄlvi���J{p�0+pڳ)��뛥��}9��pLݾ̈́�9}׊��v�&�YY�n��֮��/����P�R?�p�u��#������6���n�i˽J�L��@���`��!n�e����.\{��7�3I}l��n�0����^-�:j�~�P���O@̥��NgM$mG�ൟ䫰�2��k������8��a=}锴��cJx|m�/�$8�E�|��+H�	�b�)��;�T�`$<z\IB��)�u�
�g�Q�q�2&���X��=���ZӺ B�S����dW��P����{��E�����_���@��"0<H@e`��:m*FJX6toH��lDmS,^�1I���	���:�p\͜�o#��TP������_Px����	�W�D#�DO�k��G16�x��&���E�C�� �%���k!a_#Z-#̋���:�=ܜ?�nVH�/>E��r`X����Es+T�-�sm?�z���_
��u/�[�c+f������T�U�s���#f3 �{��.��S�\}xV�f�����,�)���K]�>5V���۰F��Zc+�`���`�J�l���5'���(�/���H>�` �ۄˆ�E�c�ZB�)��o��
����k���6�гذ΅�pܻ��Gc��ot܁[Y.JfiR�Y�����g�|�TIк���7X����"�PP��o%"2T%C�ʪlAa�l[HEvZt�:��}kWY|�zLA0���8�ѷ_��_s�y^7,H��4n\�/@�ڧG�Ϯg���K�q9�����{�p>���"
��<��9�S"�W?Q� ���[yKbN��[���D�x6ye��*$��41��ܺ��Qbv�_�\�xFW/�)��uТ��Ə��٠�7�b9 u[^ų�O��S\xg�DK/�|Z�,|�J���٤^�[�H��ػ�$'h٥���Z������fD��M�3�vT���e�ֳS��q�1�z��l�V��v��n��A�����[���m���ӫ�+��� �R@��ƪI~Rl�ه���C�Z����z��m�/ �;����4*�PI6�e,2|�2	�ІǴ���
�����2pʝ{�G�$x��G�Є�f�����D\Z���V�o�ڋ�X�d��Q�M�Z�T��^�g����Y2��Jc
�}]�b�ɮ�礸>x콞b	����(�PT�(Ү��6��V5�'�-��<CZ+s\�|@8���JN;�S�s�S�[� ������ՙ�B���W�Rܛ��^Cp������� �`�ASf_�,���J8���8��_��� ��۠��^���'�)�o3{�2	�h������%�+��>�Yrٙ�)���i��i�;�R~G�Tь�����^��Ob��u��iY��������W�����ै]mӯ`�HIf�o��4X���
�ý�S�g28~r>�9����=�����@0��)�5�p4�4�OV����2�[n�����	�c���	j����ف���W}9�]	.�Ʊ�Թ��:κ���0�P$�(��&�\�̘���~�@Kʸ�_6�>23Ls/C,�4��-�-+Z�,�q�x�/[����,t׃��7M�N��W�t�C.����!�TeUa�+�m5�*ͬdBݓD坶�nۉ֊9;����oK��H1	�i ��]�5�xqÈut��o�8�e�X��Q:�f
Cu�ݦR�ٗ�0��?��Ku�ܑ^���������=	ZY]u9�Lcˍ�������<jH����՚1��?`���
�o%MXH�*/�^Ȉ�ם1�F�S6J4R�p�{S�q�Uވ_&� ����6�X��X>�i`1��מa'ݲ��#�B��_H��?Qk�۪ +�>��Noo�G���#D�]?@��N��<��X-٠��wH�Cn��<�t�aV������B��1){m���u���o�/��F�(���-L�Ydw���I���-,C����a H�[�|��Ý�9V%��$h]׿��]2����?2D�Nz�l�P��N�.f�PS���@�x'�﹓΢��Ҏ;~4��kߝi�:���p�B�-��ktBxY9��t������\�a2����m�X��U&����d�X�i]�κk$a0��U{R�|V�	3b}ʹ�W]ys��z r���娐ؘ��-^����*��<�VF$��c"��F(�q�����"��Έ��Va�z]&��MhX�ŒI����W9�+���Z/�"�A��
$ �-�xc�7���}���F0��+P����EP�	U�y���K���������;�Z:�[���	(!�>E����8ОH8�@�7��i2�d.9�
���l��>��9��zyo���@��PM���R�>F��Vx9\��p��˸�O�-V�UO+"�Ma�q�ADsė�?��?�3E�]�TV#�}"�]�"M�QA]�6��Yq�9�D]b`[����
���$g�r��1���ᚎ�0�&x�i�JN��ǵYK���`�����/C�h�@��9������^&�,�Y��W�C������K��/�I��~]v_V�t/)F;�@���.�3ÚT��8��d
x?�A�_�T����-��\?F驥OSs�$����ٸ�x���A]����([,�I��k����i�)�_�P�<����
 �����+��Q���U�e'���Ɓ�/ <���3�z��c�6M�594Cej4�3�<�8v��M��N�w�4s�»E�}�5�v�rX���i-��5���@`U��홳���R(z�������)l�l=�	�+�}l�
����}(�9]o�-�n�Ts� ������!�������\'�q�����Rq��Q�����I���Hݔp��%���D�ƍH�V�
#�/;��AG�1hF�-�7��zx���w��Y_ �j�����!z9��l�R���2�G�P�<�O�'4��2����
��e���,����?����, 3ɕ��V��7 �w�e��bο0�{�W���zm�)TS_����jX��_S/�La�Ɯ�y��f {w��bj��/1]!-�zC,C�jOh���	r�*�����-4$Ořx��g�/�;A����I..����ZT�i�VwFEʬ?+��HcLX�cW(��"vC>�38b�1۵�4��A��g���OW*�w?1���fR�'Bڌe[T��u�u�u_���2�d}�_T),�Y�\�^V�$�\�ѷ/��JJ���G�<��Aa@)U�����iE�e���
��[)
��"�{�6"���;x��@�T��%�o)�����xU߹�����r9!����}y�t����A�N�c�s�"@G���|��o�a�����f�.G�7G�rp�O.�X�܄S_�X���nΖ��x�٧�~��-IX9�z�^�,nм⨉j�*�eȻB�����h�LÙ�^��R����L�k���`˷U�[{�^�B�T����%
ie�� ;�V���P�Y�d��%��*9�L~��x_�z��hA�!U�r1�,Nw۶(���( q*2��|� h�w'��(��h��a�_FF�fYt��1���e��