��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� ���L����ѳJ���ף�6I	��7�"�D�}ے-��KpV��s�h�n]��[��;,��*��_�H1mTu�<'�M� ����Z�H�H�#����*ծ���p����*�R@�>���Vx�Cl/_G�b)�z)���e5��=")D9d��R�d0�� x��Ġ	\�{���> �Ueڼ{�g�_ˡ����T�x�\mB��޿8x][������v�	1)�X}� E�� �_ð[#�b�$Xt��C�
w��bGe���ʹ����UG٣�ɹ�~V��e"ѦΙo�ɱ���0�-�y�v��CPܼ�Fڀ�2@�E\1l�GN��Ϣ l�iRP'�ϙ����Y������ T�*�g���DO��� f1v�\�w������Z�2���8.�QV,���W��K��� *�,�J�6��jH�;�B�n]��CKxv���R�i-IJK�vC�?K$�Q�Ai�L�����I��L1�Cɂ��[�������x�9ئF��ty/Y��Tdto�	�^�S���/C'iy��^�,��)�:��K,϶>�e4��D��#��#�a��ÉB��� m2���pv �Ah���q�ݩ#��?-����A�1	�)W"�"Q�T�y��]�,�V��~���zZtˑE�qv��C������+	�i�����Kc����|���F���o�|B5Q�L�ν�!������q�"��?����z���AL8����B��<�x4|��<I�*��m�}��E�r{���K�B
�8� ��p�P�ĥ��X���@;;%lcKrʓE���Xȉ+A�|�7q���vI+@���dK�K���.B!xW�����4��P\�T"�8O��y��_�e�d S֡R!�vqA_��n�D�fn�O����_��8y�W�y� iё\'����5���ġ���a��'�^��?an$�U�p >6��?>VT��O?���}נd��l�jnl@l�h2:پT$�NϺ'l_#(��x�$RL���n���r�?<=:)�N��:�g��i���]�L�hc���}� x�}�祰����Х:��^)��c�v���/>�,λW4��'�>�P@�)!�k��&x{]B�J�J�Y�xe���Qb��*�m<VyYWr�:��+��a�*�,F�+�\	΂��	�1���L7�&�|�prY�Oq�@ű�⌴G]6\&b�6��T_
�1�E��-TQm��z?�̣�Ȥ�Zɉ�\�_�Q[F�o]��ÉE�����l��u�	PA9�~��$�˓�Fp?d+W����8�`�S�ڂ�I��~BT)�� �)�gd]�+�!#�Dq�49��ͻ<1��&NC@8�����wH�' |���%��K��'����b�)���=3�,�NKHsOȫ��� �B�p;*Զ�G�EW_ذ�s��D�`L�ri�e�K�,y��R�"���D@����P.���~�o�l�o$��|�7o��	�������3�R�^��X=q�`"�˒��#L#,���H�����Ց��ʐ`���^�(�h�i3�K ��*�UG��tO_Ņ$�,���D�1����ej,
ߨ
�NbP���
f��mm�ѷ�T�Ɂ����Y��|lV���8(�+<����}�D�5Ow	���I{�+���������@�(�E��{�Ftt1�0�YS�����c+�L���^L~��%]�&Q��u�ty��o�z����*z;�b�<Z�y6����Bi*bq�WmcC�{{��E���7��N]�E�YWL�~=��x2�L��AJ��u��ȹb��N�I<�R$ۑP���^���O���ZJ�J.1��ߘQ7$�_��H������;+at��7!��0��ҙ��I1�0��s� �2�	�y��@ӕJ��tʓ�#4q�.�n^`��<�E�����E�����p%g����δK4�b�_*Ȼ���咴�Ql��e6�8/5�3�s�^OL!.�ǐ\z�A�W��osq(4�F���c	��t!4;q�W?�j�,�Ey����ס���9V�;E/����(S,T����b1�1�����{�����I8ْ��z	��+�)��m8Coϳ
���R+O��}��q�J�?Ot��O� _���14�7�\K����w���/V�I�ʈ2mp�}�CRY���=�ѽ�i09��]�xYe�����J�����߻tU��q�8w���p����Ƭ�'S���6�2��������w�}!ÿ}����`�k�a�%������4h	]^�;��z�eAR`x�Z�������V ���O� ;Qn�2�JᗌV������(t�x��l��M��8�,z$��w�0� +?���FR�h�-*�����X�n PD��}�ݞ�ɶ0V��6ʐz5Fg�;Ɂ������Q/#�t�D��y4�y��6�{V!n�_��c3�h�[���f9�l�~C�u�ih�G8�pe�֮1N�H,�h/�����5i�H���PZQ�c\��g�rV��`����iM�'��ˏvs̽��(�o��J|�hR�ۀ��WM��ԸKթy��]ū�\�Z_���!��~��+��V��z8��u}"���1��D|�\�q���8P�����4�1���;�5��x� �;b2��dT�t�)�� �S]o8���������nL�Qא.��/xε&HMWZr�)���YA��(�4lC��oo�1N�hh��{�2�����y����_�Ɵ�w� )�I����Rh�|¡�8�dQ9����Gj����;T���A�je�;�p�&���z��19�B�à���m�M��_�yc���!�����3�zQ�#b�ۅ�`� BP
�I�2���`�ș'pR3�k��k��|i% /F�Bΐ��qbY�cH��&u|�h��1Z�%�Y�v��Vd�d[�0�5�5(��� \.1��[(�0j��p�?-ՅK�F���|X	^�)JR�娽�㨺gP�0���������yD�r�M	ͅ����f�e{�{.y[$��0Ӊ�F&|�[}�YB�V2�M�m[�ґ��B�h�(;�

v����Z�!�oW�K�\C�n|�6��ؗ�1/����.�D�v!�#��
���h!��&�ƴw��u��1���=~;:%�������B�,+�E��T{����;Mc�а���J�� �)�nr
L_q|K���v�,��J�&p8��>
D�?N&}ޙ�b�c��ȓ7��6r���w�78g���O?���.���I�+�V(�� �M6dBC �P�������r�3�e�"�-5C�L�v�R��H�ʛ�t�1�.F)�s~x�4h Y@DJz��g��l��C�x[|��jc
*0'�4�Xy��<�V�~��瞲��d���u�#�}�!�k0��@Xb>9;���Ɯu�³k؍Gi�a�}����{#�V��6�¤	σP>pid�YkfM�@J�;rս�,�S���;3�)�[XZ"Ź�}�}�X%_���_\E��:�>��rD�l��9������S��? �H)������3Ȉ.������+K"�7��T�7�=Ա���f�7U�|@ٺ�=�ȥ���މå G��m,p�Y��0%z�+N**Ek�:{�+�s��?���p��ꮆ)�j�@���N�c�j�����V��!�]�yB��߾�q�:� T� �L��q�f�Q%�J����d����W��y�Z��,�"m���<y�ޱPd�:�T[��9n,���j�����j�I}���}���*8�-����U�KҌ����� ��$P���]��O����px�������b�8O��(of-?NU��Z����^�����h�k�}	�V���4Y��/O
b{�LYC�;����Q�
aك^�`V]u���� �>r�E��bA��Ь��k:ԅ��`h%B�;:5��*�	]�īv�E�Xô�ͬ��Z�OG���Rp8�!�Ĺ���q�$|�3~k�W?�
�ڶd�-�� l�c����{m�A˛�M1a�^����~G�|*��R*c��]�)���]��>� �����
���S�{8�o�{7�g��k��x����N��s�F\��J�$���|��bq�>����E��Lv��C䠠c�hH[Wz7�������0=����F�dV\\���ۖ�Z�3 �M>_f,�L�񤝓Y,������Z����^@��l���O��kq7*�&�͙
�6��#��ˊDjC�rb=�\�ig��j pz!��D�3���P��u9ū*����;��Rh"qo�#�`+��^�Q��.��B]���2��S�Rb��z�/`�l��!���� ��^�#�g'�7��J��S;
rNһE$���*�W� �l8��^ܦ|@���ŕo�|�1����ق�:Z�=ǯ�U��v�=#��Ca����P 6�|R��aj��59�љ�6|�yLϮ�����؞=S�Y����kf�E9.��m|���`E4m��R�h�g� �r�-�ܸ��mQIH������^�x�����hF�Mo=ɪNz�v`��@�D�AE��!��Uc�e	l��\�)��"�g�te���2n:"4�Ʃ�u�R��PHsJ�A�+`�`
�P�w*�u=��ǿ��7/��U�3:�ZP�b�����Ā
c��o����xܞ(Vջe'd{��h�^nޑ�νT�����g~�"t�ǜ~��n&�\��xS���m���=>�X�q�^���{õ�6۳() SM�h�O{��ͧDv�H��kv��~Y�Jt��;`��V���t�����Ce`���hp��D*�W��dn���_���ϐݕ���.�1
=����3�0�ʹ�\�(]�O�(xn�^���g*�^,Uu	�
��J�E���?6@zd"҆I��;��5o��}������T�l62jJЭ���&DRȴ�x8���Ҝ����E��\����fְǻZ�n9Z�-�F�%��z,�u���!���x�/9� y�
\WM���}�'�1����2�Q�tQ��o�O�L����A$��g���V�i�DYT��h�1F9�!��Ɂ���H���v��4�r�?�(�qE��U�(դ����z��p���;_)`̮�[2	�`��� ��_C!Y�ܵ��f�e�	�rSS�	�;`U �j���Wdbj
)Ĭ\�jP�gQg��h��B����<u\v�����(^6��pr�Y��1�B�IĶ�op�+�Y���_95@�OCf�6�~�N��.���@��Z`���>��E�өQ��)y��T��A���Ɣ�7N�k_�-��f�-ן
���`��u�U�f�oo�m�-N�5������I3��˕ޯ�^�0��w4OS�*�$�w�	`*+�����$&�/�mA���^'���a���޸X���K��{�:�>F9�q�ڞt�?�#���2k<��!����}'�g?0��9T�H�[�^TŴ��Ⱦ<9�e�XLD���هƔ�o�#�*n@"l�M6U.}tN��G4�����&�D��O��Ϛ���a��'X�Ĳ2o��")��FK�͐��T�R,��a��-��x)�˘��]9_#f����'��[��*�{�.h��G��l=D!=�wu����(����&$t9L}�D^�M��0�OT	��#g��ٙ�W�^�`���L��X.��6���G6�ȿ��� 9/�O��Ԃ!hK���V/l��o�W{�Z?��ݬC�� ��7����g!ݢ�����~Ԃ��ձ�T� ��`N�h����a�����V@vk�Kڇ��x?�Em��G7c�k�.�aHn+�1�cz\=���q#�@An�V�P_q3mn9�cxX_���̼�2	g|IŦ@���"&��y�Y{�y���}�o���Ey�6Y���F�C!P�NϷ�S�<�Z�^�'ƈ��D(Y��G	��t)�\hP[,e���r�呃��A�j����b�?�s����>��Rӛ�~��͞(���6��'Ew=�������uu�Eg�r�	)k}�	7K����T���~-��G;,�+�Y��^b��1�/�A���+�"w��sS�֡�	����J��TY/�����0�*4D_�҇����6�R�s+�85�33��)�Ţ?��t,V��� V5�>ܴ�e|!$��6TV�#Rj���2��s#�w�W�B6�ߣ>�srtM�1ZNh�V���ZEb�~����O���5���b�����h zJ�oD:$���T	g�r3���$t��41Q���:O$��wC#C�$N���#nv�U���D �����_m"��]P��d�+�8o<t&|��iSak�u�M�r%����X]��4�8���,ݨ:���� �3��D
�ʁD>Yl��C�M9���	��`H\���㐖�=�J�Q ~�N��!��1i+B�.z�?b�D���n�a�@�p<��r��\�`d�\n�\񋙁����%L2�3Q��r_Q:�� 8���3�f�͇�N׌C��)�Dx�i��9:Γ63�fa5��/~U��F&4���~��������7Ӯㆻ�8Lm��k?�h��]ߩLW\�9��JT�A�k�m������,,+j�iki�O,���=�UE}������� �ײ ���:^�ļe�~��)�j
�i��/�j�⇜��u��0(���TR$4�F�9a9J�C^`; =��I���mm��&����U��<%��
�"O��' N��J"3
_p�!�j(}K��2^b�{E�����8�tָ��5�Q�������Cס���0я�Zp�7[��Y�o<��%j���f�e$�P��*�
Wἦ�S��4��BLwO��˝XNq.U/x��,��H��k}Bu��� ��6�a�w��泓Y�����յ)D곱��R�u	�R/v���(��!���J-�V�UG�*��qɷ��n#�6E��.��X��-lG���7�$�MD�b�{�������ӊ�1�y@,{�%`=�vES1-�� +g�s�_-9��3�~����O1k�)&��j������� �%|�l�ƿ������7e���r,�x��+�U���(�e_%�� �'��̼�J\,e�1��p����'�E��ʞ{G&������lβ���0w2�z�5R�e ��	 q1l٤�f���r�}��c��,jSV*/�D<��w?R�RXB��ZJ�5�ce�W��"S\3v��զ�!Tβnmq�_��LMݓ�L��R���P�[^E�W���� �q0Q\َ됂�f+;��Z�V�OG��:b�fQ��z����x��iϭ��*넲��R�`�6��}�A@ã���Q8j���#-P62t�u�xX���A�;��7N�6�Tͣ�@�R��1�a ��h�N`�,��Qsj������é�ǖ#<�玀П��f5@��\Hv����1�5o�}�E�k�:â���ݎ���ٍm
�;����U���ʂ���,�%<���1�PZb�P����.��Ȼ��w!t\������-�/^������{{RR �n2 :*Ǻ��@���m��n?;�Z6g��=@+�i���C����B���2a��]@�i(�}�H�C��g-6Zh@rb��}���]��r���ƙ���w�Q���x���]�[ t"v���:Wg"@���A0&@�c�R>����H�/�i�m�Z�ڜL������>U7{ёW��3��k3$��'<&w1.��xe������ ��!Xҍ���0Ck3��2�-�.���o�+�)���F�T͑��65��T�-W�5�8G��Z2��B)��
��V��}&��|���w:�G�(��ؑph[zڧ%0�)vC���[8BVbҤ�{A�$�If��M,�������M3��_{����+`�i��ág��k���(�98��OZE~-����\R�}��+	�=E���5_"�shX�,MB��(�s�鍕�X_h�,����R3p�!Y�
��g���񎜻OxV.v�n�.��8Ļ��Ү�"�e�+XtD���W��e�����g����(�o�ȥ����Z�[}h�?���-#�x�a�Î��[Ax����9���n�}Z}�C]B��@��ADHͪ'0qv�����4�L�B�(�J&�^���f����`?���̳��qd���j�{W�r�����P/-���ޛ���Oi�����0�Qմۘ?0��4o�OR�'!���0YO.�b�6�y����Q��z�e��<�a���͒�K������?w���w~jsTO���q�*م[���1Q[���|�����F��0;M�?��S^��IuG�dRx�����M36v�*n��{���>�R�ʴp"=���݄2��!�#��X=D��Ya�����׾6\n;��9�0q����U���:r�|�R7w������� V؞��T7r��c�8�"��,78x�q�]kz=h���Js��*z�kM�e�y��V��<�}���Bu��/\��s��Z����Y�Nq]V��{��w~%'m���F�6O5�{��g�wRS�mDXX��q6v�Jv��N�[0�r�#�7��s��5��wzGfd��M�͓���*8�;dʲU��IL"���ּK��1���G�볨��Ils�Z��ڗ۳�n���[�k���H�!G�p�0���d!w�'Ue�-�	�����S�CEӐ�f��u���a�k�?�X�ʊfo"<�{���m�
��L�9�$-�F���\�^�[:�/��͆���b�ٲ�d=��bU���B�(�H! 6�����,쟹|j��/�=��ζn?��r$��N�j3���UT wnGTu�@��KT��/Ѱ�D���V#e�ݔ:T��wK���,V	kiMv��/�i7x�XC������i�a<!%��Su��?L%��6����V���^�'�����X�lxsj���S�jmA!Ա�D}ݗ����Q��.��.6���F����x]��ܭct��^�̭�t�r��k�O�,ah�DԊ:��K���|vw���ͣ3���l��8%�D��5U<lE����Hs���*��5I�5�1�Ep�<��_V t�B��:�8��_���@��"��kfzY����[����[oPm>�d�Xx/Ϥ�f��qVuV�I�L�L�,�6:�;t�|�O�h�2"��d��J�j�b�����W6�jι�e�-�t��[W���h�%���!|(4+�X��(��3�������
-n4�����@�/�5��/a�,�[s:�ہ�����?�wG����W�{�=�WAs�NM3 ��n���`iy� [WVB*5�P����:�edd`����)�裑�?3N2����+�z$��Y��NC|���T�xYZ-� �s�Cl�2M������p9I��H)	�|c�Tbن���밟Z"��]�C��s��6�";�p��,	]/8��M�L�Z�k�"�m���ݾț.�ѐ�F	�:q�)�m�L����j�v���^
7m����ݽ�TR����k�ve���8��p��Q��B��qf�+|r X�=�&�)�X�.EQ���vۆ�o�AG|���e�(W�K)%k�Z���+�$�Nc�k	ح�u&xSG��`<n]���\�%�Z�IO3b`��2�|�cV.��v"f�lr�]�x4��i��v�0[��h��D����l�"��Vw��V��TN� *�(KD WS�S�!���g���6y,�Z/��W��(�gR�����-|��j'G*}��X3G���A\�u��C������l6�P28��\��筿SV7:�����h�a��|�Ⱦ�q� ��E������f�NA�#`v~q�H�tqn`�� f�0h3��h���Gl�����
]��|��_cX�/Neb�a��!:�0˸0��7$el����F}3N;I��p��9JM�<1��7���;R(��>l���a����j��]9�� �U����U��0����g��./�1�!����rSJ��{,# �9���Te��ٿDn}R�\����w��E����U�;z��Ձ<�ϭ���`���t�P�;b	�2<w��Tԫ[�3R�߇*�]�i�?ı9~�ߘR-A'bs,ٚ[�5u#��H��:f���V�{t��"�A6��۲r�zz�B;���Ʋ�r����aq%ɍ�����m2��av9���O�����ό�F�I�W��G��4���n�`M�ol<]b�#��:0(�&֐J�qf�1Y�y�(J���6oJEh���Z��c��}{?�1=j��1O�t�Z��I��fG����F��@B�����ڊӎ(����������ˍ��}D~[?���G��ٱ�k���dU$w{����}{~���Aѹ��뾯.[B}zrRpL�����QGgt�c���������m2�Y�פƿrT-���ݱ�xgζ������1c�f�nS�z���fҩ&z����6Е�J��XWcd2��ޚ5�􏬛JA��lb��
G�r��ʞʹ[NKS�H vq /���y  ^���	���G<�sGwi��_ϩ;|��9-�ӱ�J�h�\�ZZμ�%[G��-Iy�/�)�HG"%����╯vj�G�$�Ԩ���'��/��bVH9  ����a��5L��un$N����)�HO>��-gb&>i�"�e�=,{x��x����wu�; MnpH���G�i�[�l}���NM�����m���2מ���D�u�n%!�`g�w	8�}� ��T+�����ݸ�x��n�٠O���.Y�@d��]r +r�yw�#;x���|\:3��Q��s���$�Ǵ+�%���+,>$
Sj�nG
�d,̳3ȭ~sMkԡ���p&Mn���@}������Rk���^�j�R���-�	x>*q�b6 e����4�k��	�R���*��(sV�ӵ�qYM4Zm	�c&�
x ��,��<��!�*%�ё�0,~2��)[(���zth�; �	\�*C��P35�k��4�����o�����Y��4L@೧�r[��^m��w���Ӳ���Qst..���a��Φ�`5�W��S�1sM�������F+e��:�i/���x��8h����T5�W��5 hNԺ���P���%���l}B���_.�?�����؎J�eM��a��
��[0m�I��Y�*�h[����s���g�A�m���#G�2"�rgR�Ǽ1F�����y�в�Ui$��"���gI13���f
�w������PD؃�(�^�=���/v\�����E@�
Ӑ�st7��?��Mlv��e�ٿmma�&�D�ط�q(�H�����Y��'u��ʺ�9*.3q�5"m��pw�N�g��k��Gf4���)J�&�xJ������*�%���B|����(}�r�=�i"��,.!U|~g;]vp��z�Oz��/X��a��F��%�La��5&�	�}�:/��n��1�x�vJ��;��u�F.��c#�wo`��R��¼�|{��Þx��h�lΦ�������i�����Q ��\S��NY��z�sPvA�/f�is�s��k36�9�\A���ΗE�E�Eg^Y�@k�*���WBP&��(��)鶠|�Ea%s_ ʠ�(u�v�"�ݔ��t�|�<�\�7f����>Y����0��z�w�eEx��(���
��Gl~�T��+L�!^��-L�+����޶�y�U�(dlS�me���c�v0��zS�jv�Mդ�̮����c�l�=�*�Bux[TQ ���F�����(��~Fs֊f�p�bL]²�
9��@���)G��;^�M�lU�r���q�^/NM�8A���� �u�8_�����Wy�a�.��rĎze2(8ɰ�e���|�{f�
��k�}5A�t�'n�mCZ$\���!j�b�~pIa�P�����W��~����<}pk�{�7�V!��-��,C$No�Č�����XJ%24�zFY3	+����97�x�N�C���J�3��	�s˶��	mό�GȈX�����aU��ڣ;��� /�J��d����E�e|vȻ�_�`�f_��3��no�*���ϊ�՝.������9�1���ֺ�ؕ��f(�f��;����d8��5��g�g]ӛ�=������#��XM�|#�z�z��ь�Em�T���٪�lYP �awF�ClC�<Xf����C�p�ꚦ�\!5!V#��N��ߕSy�����+�fg�r�C2,/e�	m@�����u6֒�\���;�'D��&�t��k�N��YjŒB?�0��ȌIipgs������PgBs�-_�"b��/�d��2=O0�N�8��<���|}�t�zb� �o�{5����P�+&���9L%#8�8�.����"��w5�c��
��~[�ַ"oR4ȷB�����[�bڷX1EuT����J�����F(\��;8uI�Ŝ�E�5�g�V�����`��HM���m�&Q)��$��K�E
�1ϱ���I�'����"�i�VUS�w�U\,f�tq�yg���#}�9x�>���g	���<�^&������~K|я���z
���$�hH�c��2�=�w;j�Ŝ^WGw�����K�U��_O"5#�	p1	|6`9��P-vD6<D; � �I��O�)�R�s��e���6�!1te�ʐЦH�5s,v��Gir#v��u!���$7N�}��V���z3�'����#
� $�ࢍ �ZɾL��'sL��qRY�dn#�s9����|�afZ�g�`��݇��Aآw�-��K��}y�g��/4CYj�4�l|���ї��gzgW3�@�lF��HŶ�kĹ�9�+�NP��=�7�&^lq�כ;�yB*�) �❇�����۶�����/��r�B�Joki���#K(�1ѩ�26I�c>A�����)F�>2�;��k<Q��&)j�_�w��h��\���TT}9kVV��$��C��E�>�>M�#����O��%x�Еx�GE!q��Ӻk�Q� >sߌ�u�~.�靴d5��@G�C���T��h��,�<�c���f���m��d1w���I��Ƕ�~u�=1j����Y�q�A�Mw�YTZ;�o��%�?2GhHQ���U;�C�M�x_�I�������#� �U,e���o ����(�@1��<���B��'��z��a,$kGi��e(4-Շm�!��ւ` jvѼ:���l���g�Tw�Uٜ��b�FY������G���/�~�{Lu��#xF*�B��
�qwq�{'�/T��-s|�Whw�y�-�Jq�ts�_5S��M23=���zmF[��ڒ�G	?w����+Ԗ��ϫd�K���C�v˒%A�Pd?�*.�W��)�ͥ�!
���oC�_5�O{!�9uk�?�3 !T�+�۝�0��B��B*��5^=,~t�3�B��'|�.�r�������q+�ƚ$�8�H8��G�K�h�~��8�'	JH��f�������ڜA��dip��CW��dG>��4�,�{�z9��߅�U�CsA����d��9�3�4�2�[��e�cp9��S�.g�R�~&��3���6��� 6gmp�`�7���Yb� :m'�t����a�uߟm�ڞxCVᤡ�>��5�·È��?�5��r�_)>nV�$4jK�{zN�崾��a&�(��As��f���`m��$y/[m�P=)-V�>&"
�HnѾ�!�� 6k�5��Jץ���S{���̟a'څG�Is�l�I���w���q��TVvB�9G��߁)�nu���� ��-����2Kf�GC�
�ϵAϪn�K��6Wy !J�0�pM�Á�re�Q�%ҀJ� �y�Z��4ڍe�Rة^�)g	�ɂO�k�W�X��*\�',E#�\�C�d!P�T	*�;*-���=c���䠊K×��U�(})"jR?�n�M,$�+��_�[�9�J.l��y$}?�	�H";aԙ�9��^m�x���
�ྭ0
�'��+��ŧ��X�!,���?��H��c�,
�y�x�(R[������8�}#߄�l^�d������f��U�ꑡG]_E�A)��^'ԍ������۪?��p<�K[���Z��p,�y�]��^O���%��>g'nO�A�t}L�%裣�c*��
�����Q4$�8����,�����TW鐾}Ʒ���9P��������K��rZ�:�Ti a�	��u�ԧ����>�\ �z��-��fD��m�И⼉ē�몿K0'��a�q:��fD�i`st��B�@*Sս�N9�?#��$qm���*;���\5aVXvz�iz�2���<�6���=����,��	@����ET�!dK{K-~M����wNeIm���͌3�=�&#�Ac�2�����o��S5�ӣ��эY�3r(o��e1J�b�Q)xR:nx���^����_?2��(/�#�G��W��b+}�0�c�(=S�ݢ��Q�y>,�f9r��ǃ�O�(-���?ڳ�j6�z�]R����؜@� ���Z������ k_9�œ����V��������%o��mlA�c'�G,zI2���(o>�q�����R>�H���o�#9 �/���������#Y��P��ٷ/����#-C�`!.���S���(ۧT+�Y7e^؏9_ ����`T�G��Z�g��ĥ "S���M�������1@�-R� �5w4�^�F$��{�B~�A�PC����Mq
V��&�@s^���[',+�t��5�"�X��(�/	 ���an��f������T�]�<�s>���þj�����焧*�����;Q�ץ�����6ii��`-�j��I,H�K哻۽EdB�?2�S��7E��c!_�����
�ڡ��	K*�QX����B�X�&FQ�����
���N���u]%}��&�*H���g�tׅ5ëҴ��N��Pcs'Ā����:\�d ���0�D�Ή�M%���U�?�+��;������dƏe��$�$�:r�(S�e�D�C~OQN���{���jy��.Y�5ƻϭ1-�ǖ����Z�7��]P������%�>��Xrh/��AM�C�{#R8�Pc�\�²�����ٯ��
��熸0��߮)���}�_ ��r��\d��`#M�v��Z:��u2�7�n/'�r\�(��e��1<�f ��(�v�&��|h�Pn�ǡ�aM�D�rx�~_�|��r��`�H��Rh)X7�d���#���p�^��ѽ� Ѵ#1B�62ĮО!7u8��Ϝ�����(�t�y/2��}Ք������A�e�
��REv�	c��En���IA��C"�� �	��U��V�R�+���v!��d��r1������f��Q��93��{.���~��5�x�&.�?�a��dc1�7v��
�]Is(mm�z��"�f�	(�6������Z���x�U�e�秒XI��������5A�N���;�E֕-+�M�`9�}���o��*�E`�]+������o)�u1J$�,�i�80)u�M�l0rӔ���2!l��[y�NB}�Y�/�������v��e��@M�=W�W����ϫ����3�"�ݭ���ǯǊZ`���4��lrX֞��Gf,mjdx:c����a]0�~z�B�<���m1>ՔK�ԈK�L)^O~J�Ux! ��g�}�E�[e�k	f|��tq �,\&طս���6��ƒЫ�Ls�t�^w��U�O�_��P[����M,y��5s
�����3���xDcGw_�����#>Ά����в� �,o��Q �'[��4�yY4�T�c�û����b�ˇ��NC{q�� T�,ז��ɫ�����Jt������uF�B���a�~��ƃ�Ӳ��M�w,�k,h^�R��GaÉ��vٕ��~�0VJ���j����$ܵq�7`V[q����j,��M�҃V�����3:�	O����<��2�^L���-�dXi�+�SZ�o:�`[ֺi�%C����p�*a{��)w>|m]��2��\���w�\W���3D%����0���ʛ:h�92��d�F42�����}L��0C|l��Ñڭkʣj��8p���@|UB���tP�i�V^l"M�e	������j�4��)4��d]n�������]�~(h���>��j\ *��.�%k1�D@~5fe�^d��E۠[����4d�R�1��}+l|4$-?|����M�KLrC?NB��P�1���Z���������C�1�K_���ダN5���6��V���@����L�=��/)�;BN^��V��ץTKg��r��O�z����C��y��3kvld�����B�QT='l�ߓ-Q^P;�]�1�+����ޔ�d߾�2�%J�u�ȷ<�w?�{}@vXu��r���K*4��w�u2�zd�M�A�!5�Pk���M��cZ�7���6dѼ�s�@)	5kb���o�X�*��ž�;{��A�U�����,�ϪD��wT�p���w���Vj�����W(��5������[I(_����
�Nlg6cSp9�1�t8���gQ)���D�� �&�u��õ�W���M��=s_�~$��&s�VO9�YG�Rƥ�A2ךۘ�/v����)�ѭ7ě�y�:D�w�@u���؊��E�j��Ȳ?^*�d|�mTы��|��[�?A�bn�=lIL\5��IA���{C���b#�[�'����~x����k��ίm�(��}	-��B.U24<��)�e�����ZV�m(
���ѺU�2�60kX]�䨍�Z��E��Iݤ�L���ᐢ��z��(߻�'�߾m��#ē��'�J9\��x��3� ��s�ߩ�OW�Ei��<s=y�8ހX��4���+;q��-|�����M=���:��(|�)�t4z�ˮ4#a�o$7~\�8���d��T�W����P�p��T����^ܔ�b��v@'���ط���-FH�y2��0hf}yӽ=�un+m���|�t&��xw�΁��=H:1�aZ$�{����T��2�Ϙ�C��l��~��B��^L�����-��	���d���{�@�# �9)�x��H��Q8	*8EV@>�h�x���`,��a놛~"A��H'�
~�;?w�v�ܡ*�}	����������.����^�%�nB�}���N�Q�Pw��^���8�5hB�"����~=ڥ��- ԣ��=٧z�UܝV�-K�i�p��y��I��t>��ʸ�T��a)!$P(=$�^���(A�����I�]��N��u�TKU�� O2x^Q0�M�Q̎;$���.9��`���"���E% ��L����ʊ�Q3�.�%��//:�c��nu���mǙ�i;qğ�	X�=��(���	!�乚��{�%����@��\��
����pQ�n�ת��r�s��lm�H�xs]���#��\�*	��k\�Yp �c�T�%x	
�_oP��_4�{t�Ś�m��/��Ɲ��رh�%N�5Y�S� �z�v�XqeQ����)��{��)p%��rksx���[�^��X�3(O*���}t�H+� �WI���{63��{��y��C4�Y�ʃu�@}��Į��Y4�&�c]gz�]���_�õ?`�)JPKP֕�=�J�E���̿O����el�-��ǒQ���Pw�V47_؂0 �|�g�Ɋ{H(a��j["�A���`�+�0#�2L���M�?ךW����$�laF�Z�a�ʎ�A��O�)z�W���J2a.�*�"�4H��7d�6�̐^~-۬��D.�v�*:���/�q����g�J� �؏PU}��X���ElW� ��R�V2�A O��߸��6�0�X��X�5��f��d���\�m��R��/�Q��ڸd0���+�mû��mF�L�`:Q#����U:����_��j���yS��EdrE뫩5ql�$�8v#��;ǂ/�ȹ�Dt�$�YWY�F��M9�J�W�(�0v��IY<x��N���r�ۑ�P�gY֑�����'��k�t�l���Ftɱ��F�Ӝ'x�n�l����j�.B���� �K2�Kޟ���K�D �m���W,�*�&�t�?
�3k5(���Ly��ΜB��[���1�!F߼5-N�Z�R�e�����)PO?֤�g%����[��
O��=�
GE �3`�ˋ�^��W^v�A	!��{J�µ�3%u+��Zm���@��1�o}u�������jj��Fxmu�h�>�x�ll	�W%����	�G؈E�5�6����h*b��A
E�^@{ѿ/��߮R�h�L0�=���
L��D(���4He������Oo�%�V��|��!����Zj�
2r��6K������" ƃ3N�!�&\(�c��Da�#lk�����2�����V��	�6%o$��$���9���
R��l�F��[��i��x���S*��s�RС-{W~ލ:V�0���?F��~Q�𗷶�-LC����^�B� ��Yk��]=o��K�t�ֶ��*�0u�G���س&@���g����@���D� E�����$l�ƨ&�35��tٟѾt ��U+u��y�,�����<M,i�k�]�H|�@�]�8���H޴_1��F흵o嘂
81Ps'��+ޜ1�{ȕ*�*;�x��d3LO�o�@��ĜWs��.�A�3x"���N�����%� ��9u�5j����N�h˫��}�Q�Y���W!᫜~�MdJ9|�R�� 1U���.���*�[��F�>P(;N�j��Z�VA{ӈc�|O�uI���D�����5B����&)���3Mz�y�p?��r�T��"�JCX��Gc��k�X�)���+���<8�Z>�M�@wC>�=9tV"��a�����d��=r�>.����r�k���NwnK�"b�Hd�C:�
	@�v9f*5�.��9P��\�@��$�%���tlB��6�8F|�8/��Rђ��%ɸ��J�v=v��JkHL���o�m��PK6e�d�.�q)��T�>�]����>r�[:\��o�6�?~�&�BR�̘�.VA��iG����3�DZ]ȓ��5��/5��"����S��``�G� ��x-0�#}T�dJ漿3>��t������z�x�F�A�>e���C�5H�hcU?��vtX5,zXwk� ��+�ȇ��l	���IM�Pf��l],��&<�m�(��Љ��LD�wc������MEi�"+��F�Þ���$��Řlkz`���6M�x;�w����(p��0T�u�vJis�Ċ�2��5�����憺�z��㬾T�N{��O�{��a`]��+o�$���A� ����������ٙ2�fL�h3��/�4�0�4��_S/]������׺�5�Q�w�c'IOs�oٛ��j��
�*�����9��Mmǯ5�o�喳M8o"��k,:E�O3麲�Ȁ�>�B�#�PH��`��3{��f<	{O��- |at����~p��۞q\��)���,����j�*�>���Ȇ��7
����P�z��C��?���z�N`6��(�R������3�.u��>)*P�Q����f��˞rFh�Nz�m��@�\�i2�ԛ?�8Uq*�-.���>� ��+g ��W�-���E'���m4���iD���|�f=��S��In� �{�;�
:w��S�ΖL���|��W̛�.��t����9�ڃ�V"05$"��R�-��1��O�`��;xw���/' x���L�j�
�}�닄�C����Q�KY�I�i�!\�*s��nٸ�����X�n�ԆM�u(���x���m
����QfXyF0�1�'�yU\0t/=]�d�0'���2��1D�qvq��C�,2�Ek��g�Pކ"����(j��yF

3O����ޭ�|/��8�F���C��]e[���0��}����4ϙ����,t̻�h/�ڦ�M���RS\���3��_���Gf��DAK���G�3��,G���HwAS��\N�3,ۭ\GRF�!���$=c�dS��A盤���m2������L:���a�Ua�����KQ�e���e�tlR��fLy��c���";P�4���,���[�+�i��mCC���::T�1��22�]�lQu1,�[�2�o�-4�'UMx0�^�X���oU�S�RL)	kݣ�o�mg�,=��}��~�.�X.�Ug������J?�q��Ǩ�ǎ��qܜ�s��}u)�et��0��B���GaL��&:I,����[�3t�����3�6"!+�v#v�(�0AC�G�j�z+0�!���%ψY	����T98�2q��[bs�q<�M�&E��5�]1O���+VKq(M��l�he���#��~?�7�i�m�����C�ic���=����%ͽuR�����ł/&/$޼��*v� �_B�gW�A�WhN���/?գ��ݮ�y����7�g�������20��<4��r��a�ʌ����hY��������7��Q7�8d���7���lwUT�5���̖y�"QR'�?��R���2�L��"�R�'��@��K���A�w��)�呁���Z�b�l���γr\��s��i��&lh�o`eRƦ�U�S`#Ė�ك�8�\� Ơ+>�a5�)�v�8d�B�^`}%ֹ�O��V������~�Q����ux Y���׌�UTK�!�� E�O��59אT��0X;�':�X,�a��P�Q]9��?s�����4��|�8��\�j]�[]'q��ƵR�3�u�w�@K��l++�07��-�!�:Ȁ�\�g:�۪B����V���`�P�o��8|��{�>�+㌆JY�vmY��Ԝ����#\a��Ҁi;65k�o8��"^d�����d&g�g%9�&��ۿðx�S*KK�]L�[Ի^]�Ѷ�� ��5��V}�oh>�C*�7���l�`u8�'�^��`�!�"�RS����TTd0TF�A�恐b�R�w7�X��oMHo�^��վ��K�HR2ݰ�7�͘B4ʲk>��O��J�����:���~�����@���H�"2��3�,w���
�`� �qi�0�h�+�0�~��	;���U��|߄/��R�z�{�sk�u�F�����+\җ:�Z�)���Hɕ����"hdNŜXZ��5v�k����J�@:�u ȵd!��u�X�D���y��҇���d�y�I��'�������p����qL
�k
Z�C�^����gE����r֕ߥ0�Y�6� )YiF�<?#��m\�
��$������5ԇ���vK�%2�+������l�sQ��<�x�����gO��5v����]x���ҧB�� "�9�������+�y9M9�l����� ���������2�Z�\�J��.'��%�WZ@�gE-�s���4�9�	%u,5YS�Ͼ�e�pK�z�8���4"�s��W �1
�g����jJ��<��#Y@�[P_u+���rsw����%lq5�+�2eڱ��ӑ��i!�
��1��©�O��!l�}��:�	'B��O��@kzwPL�#<+��3_UĦ�r���v8��,�6�$�$؜�F��#��	�u��������c�u3�5�"jƛ��bG��^��M)�������!��`�
��Fѫ�F�ڰ��,���WUc���˺�+J�SϢ���
w��L�.�-Gg�UBYo�8�:ۈWq�Cfih�Bӫ۬�	[ɔ����)��5�"�������1�E"��;A�ܒ6h�:���%��Ƞ �9�O�̲{L�f�6� ���yt:�V��<��b�]rp5��H{��f9�0�Ċ�k������?�Q�̇�-57gr�#w��#K��靸���Q�'Z]�ő ����{hp�X����9ra��-��}�I ���Z)�.-x�}�	���6�G��z;��؝r�4�
�,AV�g��צR�}�%'َ`���(H?�*��b���A`�&	�[����W������|�!m4����Љ��J^�kf �I~A��7;�}�T1P�Le:��3t���+�$�g�/�E�VJ*�Y�e`�� 	��[~x������r�|}��^+�TR��3$8���+���.o��az��7s��Վ[�0Ma��/�,}l�G�?��s���Bs��4<��! #�0�u�9�H��k��� �g�'<��ג��l[���и�b��/w:��:NQ9���ߺ�g@���L�����k�Yr�x�>����z do�w�R\�u" 7�HOQr��nLTs���jL�?��@�B>(p0�(~�^�½2<(��4U"T�f��L�?�}�v���#�zQ�>Z;�3q������9F���=<P��r�99_m���i�5`�0��Y��?�[�����ꄻ�os�ѵe����NW}b~Kzk7��?M�WtcE�b�<�ǆ��GfW�0>�m��̨�hg��'���nl9�*㧭�{���l�gHo��k��Wj�Z���J��x�gk�^�>��6jd8��������8<�2
���$�yG,�� ��3����LN�j����! �B(�Q�U`/L����!eA��n�%F�׸U�ԍ��~ua�@��$T���UT2]޺��L���$�_���P��k�����C�O�6�g|�&3��q�h�+�Q���]�]��Y����'�b�̰��b�yl�1�D[@�jZ^����~�����z�����2p�8���sĬ}�����'���ʃ�u�{�ǥ�>|X<{:ڨ������AW�Bc��>���*W��w�ƍyK� c�m�o�!��+�[���Y]d�]	�����þ�b��\�G�����Z�2BxA+��x��E������.(0�#fm�Q�@<�{J�qB"i�P0C5=ֲ���E����=(|^�F�hT�̀>$LG���R|�!��gh_�G}U�0A09�O��$"Ѣ�=n�L��\LQ�z��gcm���-:/� �,��v���P�RS�����heA��	�>��_�����9�:ɂ�?�aX
�~�~[$�{�,�^��U��G�o������W�Em��
�3�ۋN�`����+��Utr��3`���pG$�6{ �36���X�ނ ����K�x�ս4�|6��m�l�|��3 ߽>�4 
|I]#�����<	
�c9��<	z[�1��?Wmݱ��a��E���0d�-_���d�]�۫4��+���aR-����m;mn�[�ź��mj���H��m�^�LJUP~Ń�JB��9k&���kA9x����B~���Q!��ˉ������r�S!ܙ߹>�x��Ew�d7NGԡ���n~�*٤}����+I�؋�A*Y������ĝ(��ӞT��)q("�T ��18����$�r�h�}�s9�4���&{m7 �����lw�u�M��5V�J���;���);���[A���҈]��\\�@nKj/G��FY�dAS�R�`�l���"���c�X�ȇ�t��n&��}M?�h3x`�g�;�N��e�u��仞a���xqQ�AT��;֬�%��e�����s�;�*g����x�usy�ǔw�y�W���	8�N[݄fo��&���� ����j�я��o��-+�x�sl�7���ewn�����>���{��p�q
�mq��Đ�7r�� B;[@:7��Yf}������)�V��@'#��IJR���;zg
Y	�|R�B�n�Ò��\״�,����>!����J�KI�T�ލNk�4�������;j@��[+�yz2Qw�/\#�֥�G���elk��(]-J����8���2�$��@߄F�.�vp;O�T�}%$l����ԑ�W�i�(@��ê��'� J�<��U�0C`$6./}�M�q��	�G�G�6]HF�-<,/����I�L9a�zzKVB/�B9Z�>x����53�!��.���'vIKQq�p�(�;ګ���w0��s/����R��0XĚ��8��������� 
v7k�.��?N�W����*>��$. �C�6��#ܼڀOM묮�Z[��� ��r�M�{!�L81��|��dLC�
*�����C(�4%�M��ˎ&U�����?٧f�F!M�Y�阄`�В�ãڗ}X�`�0aXn.�3�� o�>[{9g�A�a��(�0��%jR�T�䡭��;���.R=������]�����ys�aU����ꋴ6l�i���yǛ���`�OPSkK;���`�dc�kYƐU�ٝ�Yʭ�r�_b6�l-�Z��U����L�D. ��P��$1�$�/����3��E�\��>��I)��5	7=n�%ã�������T��f˪.vB!dD�۹&����m���Y*�g���7L�܇2H?�b|�<B��[��Wd�z�yD)C$�y�SJ$�x�!Ox*~�Q���@�38�Ӽo���|#��sq�c#b�؀��tP|Q����g��h�����j�`H@��0�($�cP�0o�ubި�)��g�0�m<n���R��ʻ��e[�DTՇ���%	�ux(��N�dB"�ce�3s�Ya͊}�f���f�^:����#|M�'�\�}d�k��&�%0���m�|M|�����w�W,�~�]ŉ�o���2~��#�c��Aq�(����g���J�� �mP^�GS9���2��;�M(/��0��=MX�$}�zS�b*5��u�0����i.��4O�y�7?�-s�!Zz$��	5�2-'�h�����|�^�ҕ�X��[iO��^/:N	QrZ��)W}�ɘ�{n��NVA7��i61����5��sj��ndzC���Z�Od�C�r����R4U�&v���sc Q@�q~d������6��M@�j+�Y9��q�����&ܻ����wwH��"���&T_D�������F��d��b��$k���٣kɒ��o?�"���{C�!�;�� ���`n �����Qθ�	�Li΂���9�(�[�=�����o��U���-7i�WQ���W���^D�-��cØ��1
B�p,��~�8e��8��"�2�Z�Ǩba���5�Ck��E͔��ˀ�%U��E,x"S��'���X%���V���������C�<ߓ��@e�w\��v�6�|.�P�2�<��U��BF���ws��:�$�o۱{��]��_U2�F�C��g
v���� ,w)�ԓ��"�s.h�Jj�y2Ѿp�D��VQ��ڊ������ ����s�wN\ӣQ�<����|��)���Z�����+�q<��B�����_�e�&�g��7_�3���Wp��N3 �=�"��4�2{XuX��׏�v���.�T�cS�㱼��o�,9dyd%� �z�P@�c:��w�>��f�-H��(mv�!���iuNVy�E
�����]�K"P.�?�a5A**:~JS₳���t�&��R����� t��SO�2����� �W4�h#�љ;wr5F�Z�`� Gړ�-���H]0nڽ"��2]bPU��:Z ���B�M�#�<�>�@ؚOH ��Ț�Na$�\�(C�-o��>|k��z$Y'��֪��&L����?̓�����t��A�b�pz��YvŘ�^9t�mXN:��~��-��k�L{�HXI�w�d2�[���l{��~o����_�r���7H��Ɨ��^l+����ޕ�d�	G��T���#&|zh�̓�ȫ\��U��~����VX��,0��T��,+���g�,�΄���R���4*�](��G�^q��Q\B���d|�
ɻ���d�0ݲ&��G.^;���C�T���Fh��?;��N�y���W6{H�*7�RmT�@8 �nֆ5��N�cD��vdGXe����Ś��Z�A�3���;��Ȍ��=�~����z�*�ۢOB�y�k�[�+��ܐ>޼�'_�"vH��po��7�[�F'm�y�f��yi��%�]4,ZӲU*+��]�c�a�2���7	��t#J��Lx�v2��5�a����,Rz��D��5p-�<�x��$CH��Y�vо^R�O�Ί��M�y��X{z6�H�^���z�Ăh%^�$�NT�5�!Hl:�ŋ���*#^�6 Y��@��m��ȞmV���Ą����yiW�W�4���/�sc��jm���6�S��>b�w�S"m:�l��u*A��dL^���G#g�#R�L�U��v�G���<ʎ$�p	
�Ą(��;e����+�pO�zS�t[�>J;���~�7���#Ѱ��+*��b��,N{�)9�~�T�ȂG�i�B�6�����w.�T��j-|�Ȟ�K�.���2��B]���M�
��p�"u�l�$��/L�{�p�Q�#qٴ��bu\���c,3�>I�k�G�W8��9�jO����E�	��������K}\��Sz?I�
�P��7\}����T�,"�1�J,]��N�iS�x�-��Z�X�*H��*i��`��;�b�:�Q��C��7q��V�I*��xu��s�O��v��*��s��"\j����U��R=E6�~{7s�^#�'j��H�c窉��8�����ؽF�uۯ�$N�$�.���T��@��_/��XVL{��N��c�V��,�=W%������q<�)y	��cǅ������� B����c�|�߅�)�k~Ӏ���I�۞���T�G;�LaT-�f�=�j%�dͻts������ZD��&g��mQ��i�MaE8���^��*ĜV���%x��'���.��6�����ٶ!���3T��a��u����ʀ��t|���ݱ`y����E<i�����I�f�%N{r�Z��z@�<�~���T*�oWyc��e+���f�iv
ף<,ծ�&�Ļ��{������{T��Xm��Oٷ��%��a��q��"���xm�Ӳr�l��J��B(��]3����:���p�X�����H�)��0�>%t�+���ɒ�U�X���&?�-H1�'m:C���ff����Χ*n�":��O���z[l��)���B#�d.m8J�BҚ�s�u _]�|\��"Q��Q7��g���7�[b�6�uZ޻z��+�,�f���hrܜ*���'�v��{JG�����2K����|��OfH������� U�X�W*&n9PJG�'
�� �]�A%�KM�1^�.�97ζ��дo��Y`�b��?'����Qr��z|�7��҉�gt֡��/���2H`t�hڤ���eY{5�FkG5|..TGP�dG�wd�l�;f��h�:>'��H���B�s�������:��W�6��̤��;)��ڷ��Z�ֺ�R��E;�g�^8k�r��[H��l�D�$me u, &����j���jw���]��->X���0�\���.b�7�L'YϦFw�u+n��o^��Y�Ja��C�Q�~��߁�ܭߣ��g J<�Cx}O�4�94�v�;����.f����JT0�������>����0m��6ތ�pf����(F�q��/���ih�����[�1󾮌�1Zq��h���©��l���|Y�C<*²f8>�:\�����4U�:!f^�������k����ݨ�)�c^�=�ڀw�A���J81�=������1�Cսc�lB�]��f�M����2{A�э��T�n�I7�CQ�o�(rK���9�$��V�6%90���z�Z�(~دꚷ{�wtt_l	`��0m�(���aI0��z��Eq���_=2�P�A)� ڇ,V?�u:���#�.J"򖩨AJ�Ŕ�0I���Ā�š�E	5�.?����K��Ԓ9o3�㉕�>��x����B�]:~x��G�*��t�P�������*c?���ƾT�,�[x��in��λkB?�4uC��w\�����rD��*n�|�f����Ұٱ�n)��:�vC�Y*���Ԃ�H�Q\��o���[���%G'Ńɬw@���b��1OQ4���:ҘP�;r���/�������6nPr?y��n>��黢i��@g��-V~~+Ohe�}���Pgp����j_�HS`��S�y[u��O �8m��ƿf����� �})H{�ﻝ�� <F��a�H=Fi1�p�(W��CNk91��ধ\�j�6�_z7��A쾥dSR�Z�r<{�xs��Ѷ�-+��b�n ���/i��1�ِN+�ɸ�L�$�)�p���<���:Vl�փ XH,�m����%��=�66e������#VG��a��b�W)<���ߝK�O�"����^sNZ-$qo����_���Nr���ʠ����M�|t�S_O����^��{$,b��8�q�#H�j�\S���X��V}�{:��p[1��ރ��{'�6͠KA_�F��L�CԙEtf�ǒpȧ2?p��;�����rI϶CAh�_�߹�����rGdlԠ@V�)���I�{��&���r7M��}���ͫ�{���^��!YRo�@Ԕ��oq�C��˶:��7rQ{1U-�2�~���Qn�ݟ��N�]_]H	[�[�1|�zkǃrLa�;�,�.-�"ɀ�B8�N|�ґ%�m���?R�6N��9��R@�0S���H�������/��Y����sͯ�٥rk����O65�^)������g�]��c�U�>=!o��j�abg�z�O?��W��h
��aT�BRM��'��8�['�W[C���7Jۄ�=D���m��P�}�1�-w��+�R>:niN-��R��Ѭ�R9X������$^hX]���0�m$D'=��z�.\�:ѲgF���u�מ��㲘��]ysJL�36<bKE\� $��y{#�G�z��c�^���9_����d
�(�mKnTO�E!��d�j�>sp�K�C�y����,sT�:�W2���v����g�CJt8�TX�q�䗅���n�aD�� �//ۡ���(~�]��#�-D\Bwh��I;"�^�L:���Z��T����T�'n�Qi.7=�ϣ�J��pY����v9P�Q��� �6@�*��|#���p�3��0�dq,v���ز�/#��i��c�":F,KT%z���e� �=q���_e�b0+��4����{6?1�:n,������bE�.-�0�|T�q1�9Ę�
q�ʫ��6ٯ�bDJ7F�P��&�AH�s���m���-Y�����y �؎�x�@��Ky���ym1�P	�(~X�X{/���@��N;��*��w �݀�z��(�z:�����{�?�x4^1+������L<M�!]���� ��9}N�|��G���Q1xnQ�+QM��D/Y��cڨp�r��Ϸ��%tE�D��N+͘�s?����E�(lA�٩�as�׏`ao�jޏ�/l����N�����q#u��U���غ%OP����
����������p��mam�+�E��5�X�o�%A�<	�#{L�f�.�2LG�'�b�0(�{�*,.��q���>y��?��Kt�-Ti�9��P]�R�)����4��fd��*ML#���-č���qve#����_���D���99�8�SΚ+�ۀ �<Z
N�������=��s\�>P��.�ޚ�#g���Ok�U�:�]�]� ��b��*sQu<$�z}'7�[����c�#4E�DV��1�r
ϒ��t(Dtա�"w�ٳr�I��Hn��WK�g�����D|�.�ۦ2�^8�@�j�r���\���_��������K�����CL/���Nē�#[�N�݊X���*c��1?둞E��!1����db�r���Co%��|w��^(3ѵK�MI�'�mͳ�ml�6�d�;p����z$���,��/%�c�?@���F����9��T���	0�������'=�SJ+��\G�� k %nS�c�-��֚l��zI�Z�������_r����#S5X%�Y	�lG��mR^//����T�E��1D��G6�=��x2b�q�l���CO$�@NY�f�9����p5�ٗ��l�a�E_��(���L�GT�>��K�΄�����|������$l*GR�y�]�ޢ����[��^$-�����ri�M�6F�(n�q�����]�'U�n�M�%����lZ@�����{C��4���+�@���R��	f�b�A ��tP�'��N�Ր����YUM�1���I8��n�r�t��|u��␻� ��S��R�������X~uV��tE7Za�l�u��ŶEBw�Qr��h���E��2`$hT-O���m�v/�V,��9���~�i2Ru��H���*0_���d�+��=�?�� �g'�%)��g��|ޡUW�6�g��APi���:��;do��)i ��X�w�~�0�����4��gA�Z��T����ݡOc�eؼ�������%�p+{4�[������hL�+�r����h{��-D���ު�K(F+b�
�u�5�����&tmR�@�gU85
�ȑ
�idȄ3�z/	¾#�ib'�S]����[r�bǪ��`����!+N�����įڟ�`%����[�b)0,}ѷ�h�$�"BuhN�%�﮸�W�l&5�(9�W�h������:W����Lf˽�04��u�����Z�Ψ�MKV�r��Q.�������JC~&��T�)��%V�T'�`��/�H��%�Fe�N� :<�w�.m�E�H.U9�9�z{}v�IAi�SU������ME�&!��͌��тц�1��A�!���[�g�O��,��#��{�\n��6�*%&�7�SS�)Ժ6'¤�LY̓{�&-�6i@!������y�-�-�1;�'���_�{@8��"Ѭ�O�;�p|�R�$�Q�0�����$���f* ��Vw�۔IO5�@���=��B	r�{��>��i��X�x�S6y��P/�-&Fr�Ц�K�C�����
�1����o�������a�j\�R��Q��7$,�N�������2A��B\i-��m�X S���B	^��~�<.g#RDl\�,�9\�U��F���7��gqb1�q1|r)��q��m����@�SýՁ+���:)[�� u2ȞQR��L`2yR�� ;T�{���4��d䫶+ɁB�����d)����[�۩��ϯ:O�pֈC�4�d�[e��mZ�_���f����z���Q�$x�뜏!s�%�[ѥ�g�F_�U�Z3�f���ū�o��#�����c߀�ظr��n6����^(RǹÃne�>�Nb㽐��-�V5��tM�C�!���X��Ά�[�uD.֪�?�&������8$�Y���p/� "����\Ǧ��
�6���K��J�����<>�M��p۬�u%+�J���1�* �M)�P�C�0�������^D�G��2��@Dk�Od�L����&�s� �Nhi��̙�t���'����[wrU�j����>Z�]}�-
ۍ����帄�l�5)u)'K�"?\MT�E�*�cW=z@"6NS���L�T��i5ʔ&���ı'�� wG�M���qS�����䘜y��� ����]������d�P#��ӣ������A �I��=kծ�8ҟ�¡;67v+7$� �q=��Z�:+���y��ќP�P�˫���nGr��Ek��K,A0u���k��t��[�z��R9r�� ��R�{=J�@v�j"���o:�97E��`SXD�шK:�u�Α�6&��9߰�|�ʠ*d�T�M��G����*�\�;���y���ݭB��ZO��ʖ��1zv��tjďk�\+67e�E������I���=��i��pϥB��bw(��A����=��|=�tn�꧱�hq�/X���C��S����&���tc�R��F<ީ��o`4�%uEz����`ec�-3; ��Y4��R�\�Q�3�qn) w�y0oC����\�م�Dmd��j��Y[}����`�X��"�:�*3�Ve�;�3��,�ɒ�X8{S�\"���?KJaPa�Q��Pъ|kԫb�rA��܍'t�����V�#�;��f yz$*�i����a�2�2�E�d�M�&�g���AK'L}�i��.�B�]N�c;_-�C<:<ؚ�[�����	�����T}Iw�[E�! A����9��{��*�{��C�_��$���!���	���]��F��o��K!\d�#��;����v�K+�9�']PZ�ж7���i"m���k�z����HO ���vţ������H��)O:v[�6�غ���)���?,'��(��\RX�'$('r�{Ok��t��Ko5U$�Ӯ{�O��'rw��g-�My���\5(፸x�'q�F\L �SB-��(����C�@������1gBD�ՙ���ܑW�q� ^4>�O6��̜!)P���ȋ�����]�1XՇL
�&�_���2O������Kb�P������j����ޟ A���[� ��@)BWF�c4u����&ߜ�X�>ˉ,QE,~��]�1Ժ����̄<*�"��
NS�X-��dxs �὎�a���B�0�U�[�E�5.Y�J
�V�o�Fʶ�����RZ��)MY�����6����~��p2r�"Ú�(��x���˰�8��6Hg,8�Z�T<�`���z��:����Ds�dwlK�#��M.�����DF4��Py:v�Ǻ���Ҥ�#��o�-��	�#��8��4�-���n2���f)��r0zE���������@%�� �G���r.��=�(Yf��˽��6Y�Eg�+�C�A��d�Pm.��ټb��
ٴ��]��4���aʩ��o�7�.�а�$FB��Z���A�� +��`�$��b�؋@�!+�G	�,����F��A��v�æ��l���g;<�р�|� :Sw�s��>�����&`�w�������Sh_��vK�a��Q\{!4E���I������L+�w�-;Y��/�-������'�Yq{[��X{�v�Fp��� m�n�oMCuE',Y�)��$�A�o�3�;�쒦Ao��s|e�f���nz*�[�$E�r|���yQ�kCl�"J�0F��Ca�v��:��qbXz�-�������#�\P��>����<Jq�/M=)�ȱ��[5}iJn��j����7zIݾo��B�
�ډ��J0������ ���Dx�5!�G����O�c�D�bLK��!m#0-20���+j6��6�G��c�79�8�k�C�`�M��.P8!��M�5��ݻNlR21B��|F�΀�K�p]t�'E�%���t#��
9;�a!.�(�嗚��H/�9�LVb2���q��4��X�@�^�N�d������C>f'� ��1X��ul*0�Ha��,�K,���q)���o`�P��s央=�y�|�]��b��E�Uco51��AjC�[�W�	HO��U8�Q��A�X8��� �[yV�@5�U����6��������t��8���\*X�����q��U(�8�\�_�z���C��JJc�<���B��#�A(͟��-&J�P���V�S�-{3�9&��oHx�U��
���/�9�y��֘��.�8@'�˶����>e��g	�8�zQ��o��
�_�:�@/
��M$+́	VN"n�u&�DٷRf��Q���'-k������J�6%��%-�`Boy����w���:�4	 N4&/=�[�$mշ���zKcv�H�wk�^g��}�@,{4��T\$����ۥ˱���fm�FM��~z��B�_F�V.�/��E\݋�A����y@���
"j�*`��VsI׿����ʹL^��b������U����w�܂eq^<�|&,� }�v�4�?����I��Г^X�O�Bυ�}/i���!W3��qo{�s��!�s%�蘶����o#� �ж�V�c�p�=�hc���6��̙s|ZP�I��Ԃ\�i��s��1�U@�U�vR_�;���Hp�jI^O��Z��=p�<hPJ݂�!�\���ih�޻�VKo�`�b
���K�4V���3k3#���5|6���[5�c�[�#c�~L��
��m�F���͉Ū}�Q�[CV!E���ҷ�8)�k�|R=�3"9M7x�z"�MĹ0��a�e�rv��]]��NO��/���lWǌ�k�4K��fw]c�<8��{�4�򼬄H�X�#�g�Q�5��mG��
�%8,� ߹����;�_�����4�TfjS%a�C�|g��E<�������5 �����)n�@(�_���\��8�s�^����G%uļ~��)����N,�Y��e�҇$l/YBS������%E��Z����r���0���V6i�8x�G����@��M�;��-ćh��Q���-�aFm_\N�����}k�f���W%_�3�	�]8��/�b��!��:��̦M�,ǿ�����3Fo�f7��݀��+j5A�e��BC���x����Xr�Ҩ"�X��~2��{�A@��h��2�~.�&W ʧ2���b�K��PT�)ڣ�j��U?q�V� [{�N��@��Iҷ�qUv�KYQ'�Z<VB��M�X5�盛Ct/ȍ��)�n���Ӑ�>0�xv��6�ރ(ރq`��!�\h��w��_;$dL��ό�)��w*[�*=���Q�G :��[�yܟS5���xOѤ��"�����b{Η堾�u�T�f���gM�\�6�[/��Z/���`\��l�)C6ꪩG4�sӥ�܎Jz�%�F$�Wp�?�����5j��vV��эS���Z�ƭ��̘�����M�7����f� �^�JT���a�Tie��K�T�L��"^�������H��3L���"�'��yp����`WӔm��/��,�e�����1BWc�jP�qM��Y������	'߽�!�R�����٨�-�/\7E�γ�MB���+H{��	��`c�j2�D�V����C�����~����Pw�Fi6�W���%�wq|'�r�	�#\�F�Wï�sWp��(�,t33�I'��$��c�C ��'�C P�+�b {8�fGz)���W?���L�E߳�ձ%$��tx��O4�rS�_���M�?�%����W���� b~�`�ro�%��e�:���JZ�i�x�>Ú�B������	`
a��Ն���2Ћ䫑z����޽b�m�A�RuKT�V�h�6��߸F��t�=������WJ&�sz�V��`��e�Y���QM� ?����l$Y�{>QL��Q�{n��(����#o���U���Ȼ�2���C�v#U�����>�� �4��!�����}�N��6��Ϭ����D$��O���KS�Ƀ1)Ch-7�_��Y(:o .�t�*rĕ����.���ggC�)x.0"Ѯ������}x� r�at���9Ĭ��&.�����فt�xl��	�:ɚvmP����E*a���w�](�U�'���1���<X���]۠��� ����d���R����Vp�zu�z��\�1�&�M��{l����-�Fθ8�T)�S�p�z��e]���"gK��jU:��ӦX(�e�A83u8r^���	e����+IPC�y�
-'������=%�-q���D�A�]aF'�~
T�H<���X�gq�>�D �ÑOkJ^S`����\��W�dplg8�|���F�2v���I�f8Dmo����C�c�0d�����s��X�����/Nܲ��r��eĻ�$�z��_�#' �6D���2��c��4��3Z ��P��֢��rE3�����s
��W�h~���ﮙ������,v�Qb埛�PGf��|u�{,�,���H�M�����&cHe&�L,�`.!_5x���tVk�+p��H�ǕI*0,�`rЄh��=�����lWzb��Lo�,�W�t���uT{i�xx�/oS�����n9!����O��zbG�N[XȷUNc~s|7I�����+d&<ҿ=n�������]#9�g��`�ַ'ߑ�i�İ`y��ڑ���w@�ǅ8�����B?�9��ݫ	 U�7���v"	��^7���t�r(��ݏ�Jݍq#o#����|�L��簟:x�XC���� L �CT���(ח/Vr�ArF4ﱒ4Z]�d���i�խ?J�h��=��e�iZ�=�ѐ��N��}�U;�<N�w�Ǔ�S���a���W{�>���2��Ob��Zh$ #�#.�~ #ԉ(Z�+�q�&@�tFѪ�����@M`���P�B��{������B�3���ӛ$��u%�gk��m"=�%(�Mr��B��T�M<��v%uh;�	i��N�ڶ�Fj5�6�'�|��!l0�v���~*YW������K�
�d�"�O��N����Tr�5v��Pa�f��*M��%	�t��G�)�<ȁP�n��^B3(���6�$)���P%�=�v 9�yGҋY~�[��Ƈ3��X�#��(e%OϷ���0���;tQ���K�+�y�/8�T�����/�aN0�'k� ���ِ*RNc��z+b�K+GW�`��F��I/Zߝ�SK؜��DO'u�!���b��n^$P�M����<�����݇B��[��:�y��z�X��o<�������h�',s��N~#L5s��nuJV�-fDS�{b��;�ژe�26t��#��d�o���ǭ �/jPo������{��:�#'<�)�3���{����SR����C1��I*��LY��i@bS)�66��F*�����]���]��ȂtD=����j�XUNg@(9�U�̏Uy
=;��S�YxА��,��ǔ)��%��Lv��&$�m�{�3*{�f���d��� ��`���k[�֘�h���~�{��D�]]M��h�m|\bN�^���������R�H�`�=�Q=��As���<���a	e8$\�w���V�%$�u<`�b��g�R)�1����$O�
���C�-�,A�V�ㅸ��lY�;V�����V1)V"B(�kc6O��K�<d!��&�9�1vĽ �Zn�cNRr(����{U��m��/g�PӸS�f��XG!`6%щ.����Ce�������B}>� �`��u�\����v��A,m�6�f
���H������K���%���$�d�hi ����V&˭w�����y�e��QYծ;&�n"��
�{���I`%�5�#���ǾC1kU�*HT���fItk}��s(�����B�4��<i�m9dNE�"�x����`�zSM�Q��@:IW��Js!�s]�3���I�V���5uY(��C(�ӱM��D?�㐊����������2�+�QPD?�|gɖ)�׽�馈�l8_8s�JloהT
����ֆ�3jP���m]�(s��+FU�`sM�Ea�⫂����ӜM-���f��'ys���I��Ї҉e*~(��
��_�9��`TD Y�p@�6 �8�.�@��A�S�T�͏0kyK���c�s�Q[\�<H͐F�?�"�zw��E��8�(���f�u����1��<ۺ����*�ZK.�iهɮi߆�q��hF��� o��������8�L9�B�L-'>	����L��%$3w�3�g԰a���9`�ʔJ��o�(�:m�C��ƀ�8|7�����F��T�42�v}��9�)R�4��T\"�)�P\W 6�*j��8d�[�a�.���2��DQH�ڲjF^3���(w;�'+��n�+`\@a�&���s����/�z4�'�+�(��Kˋ�RN�.�ısz91K�´;�v�?�`FG�nt��?�,_V��FZ��^���I�mC���#��~��c��?vU�9|^:u�f��M�p�vR�c�~�dBod2�&�>r�%+�����T�U�Ir��ws�'K+��3g~��n�sDL���X���ߧS�5��7��^M���c��U�i�'߇�nGF<��}i�{�AW`	�.�(|`��5^Z���:��w�'�{���hy�k��9K������^�Mr�u����h��4{�8��mʢJ�l`���hs��{D��G��,��ɤ���r{��G�
OLl����F<g��@���[��.0�Hg�޷w�IFh�Τ�-��V��NˢLuN|�6��W���A�3 ss/��kB�?�,��^>���֖������0�i�-�X��&��GU�қ�l��_(aJՅ�*:����{t�����|����L*�}=(C}u��PH�D������!V��D����L߳�	���-݌��6�r�ֵC�������-
Ƅ�� `/@W�x���e�����'4dp�w��8�}O�C���-;kn=�yP�k��S\.þZ���y�wZKЬ�k����u�}�aŞ}�,0~ΜE�yxy����m�S���ι�Ǯ���:y����2Y.����X���%� �*\H�5��	�s�m�3�R�:��ML��OPRJHFk[A��4{/�Y��<�ƿ�N������o��bz�ɕQg
,�K�����KG�||�Rn���q_*��OX��;�
f�Sb(T Cg��ߙ2�S��N Q���.���J*
���[m�+htI��Ŝ`?>�<$(�)$*gw����n��[�%`@�fԿ�����@�� �g�?!�
�U��G����5��}��z�m���w�q�;�>�9�����f�,M&��'@,�9Tr$%[H5�[��Oh��?n-�l�l��!���9د�0R���ڇ�#.�#�.�y������,ų�v��}:22�r���<v��L�]{(C��0��y'9@c�8,,6��+�t|*\�S�����a4�r}�<1Ӄ�hF�jl��6��xg�X������80o�p\Myj-P�~���#9�,����$*�15t.�%�DP�z4��f��:���D�Z =в�_L�����^����ӧ�C�A<bV~��+�!ͧ't����Yq"�{G7CfOfÓ�h�ܹ�+��x��,Ns���;'3mČt/���
�D�n�_ e)5��'���\�G�Y}�S�9G�-���p~�2L���t� ��ESb�)�zK
oNR�Ї�Ca�0*J�f�Cl��j�@��_p�o�x�7��w�XF�eq�+��㖓t�N
���zx ˼Ge�L�.�v�=g��PV�zo�D�?�Z��c-��f1�߄p��~BSp��!h?���}��'w��r��h��'ܠ�y���"I=$�.�0Ha�� `��9"�D.�Lk6.��;�h6*���(?�n�h	{�<鯩.8�^n�p�Ȓ(�ן�����9�S�c���iu2��$�x{��͓$z	9�@S�]/��r>�������\;E��.P<�K��2"V����yܿ�a2�-%����YJ�,M3����z�d;���Rpf��r�~��i׼'�w��Q�`�%���[�"�VX�;�\�[W��S"�Dd9�ȅ���)���"?�h
��
0� \#eʾ~�B�������+m	*�JN����"���5����2����z� )a�{���Wh]�$kS�s�D��ɽkͱiov[6M��]���\i��sk�a�sV��ز�`��>XSy8��<Nw�k*�k*��)��.�=$a��ީ�7�+W�I��<-.��hB�8�����I�{4�7.	C��K��ޜRc��q��	+��P���ե}�^�#�����ǋcB�RVݘ��SI����tϽ����/k�O�I�bN�0}�*r�r?'=N�}��ڟJθ��S�:�zZ·�9�m%s 9���Ab�nC:Dc^VBy�_{$���,hM�yų��O�'�j�2����M��ӿ���E�1�Rqx��J1L:����X��H7���� �:����堛A��ũ!H�:M���/�>!	�YMm���&iO��X���h�4�����y��ѿ%"PM�s-7���m�p6����U�}9�_�Lm1�<Rm�d�g����(�7]ٿ�䂟>��i�v]��%�d����$�N6�w�I$kl��%�/�NLl����]��RD�સm��$6�G
�A?���^�q�0���p�rY����׍���(5
�Z��cB)���D�1�\}:}���mM-���1���$Ec��kfX�f�m�+���ג�(2T�nB0{����f8��re����ƽ�3��������h��E�4�]Z�o�������-�}�~!�z����8w1��X~�цVۣG z�z�M�kc?�)�[���}��{[�w�e�'�,�:�r�r����8��kh%/�t�]h���s
�q���÷��嵁i�dC?��ҏ���������y���v�(Ͻp�cC�;k *qr������|u����Rd�|[)�N�L�|؏�*�29�e��H����卩�]�}����b���m;#	���V1ƻ�����`c�FҖ�F�״b�c������xM�T�94HSĤf�[�����E=��X<���v%t����1	q�K�[�e���ıy�H�9�Z#.K�b�m?�Q�$#G�ZHQm��Q7s[
 X�&vz �)G�ď]������[�'��)ӯX$��D����D�UjPC<m��蹥_�)��;��Z�5�_���� c
�EԠ�/uЖ���7-� B`w!��c�~Gj���<1���
[~ehܴ�Š3��QsgYu�3m{=�&�ɷ_D��������f�E��O���B�\R�Y ����N�חf$����h�;e�j���Ek�h��G��,T ��3�y
׊��;�i:� 	�¾�s��G�e��cPB��J�@����J{�Ru��P�5&��Ϳ�7�u������z���_�.���G��<1W�;y�������˟n�9/Y�3��<ͱ4l[^]��h��&�$��'���Y{����Es���7A��=������ ��$qB9n�%^��G��L���	�1�䱘��j�j8>Ӈ��ޭ��v�h���3#y%��a6��is�r��[cW�����ٍ˲�|+D3�iy���( �6&8!wՉm�t�����&@���&*�n�FW��&j�7+��9�4��8��gݥ*�v
��n�y����<^���-X�2����N��K&!�h�_�A.t朂ͮ��y5
J�.�@�/��g��W%ON!x�x�P��Q`�p���Mu&铐��|�96��W �=�<�+�ulP�L���΁P6���w��8^�̎���q�/[]複�8��B7iU��b��k��o��^��E[\���O�dP{�X��d��q���1.���D[�U)����������N3{��#C��T�R�8�\B�(�l4x1���pk�(�"3��Ό�>�@�z+�F~z	�V��, >$P��V�˦l� ��<�I�o�@QX�8�Z*��=�����J$Dv46*|�ԫ[�!���B^ms}RRR8�;�X�`p\��	��Ft�p��eN:i|�D7��-���F&%V�=�w:Q.®X�=Y���p^��MT��.�o�gۼ�Ԅ9���ŉpHv>W�7��oPrr�w$��R���9D�j ��&%y?��D�-��`��qeL�`Ch~��V��������v�\�7>@W1M*UW�y�*�eMۥ��t$@թ���d��"k[��e���� ���}�GO�ܷ��Z��?��'|]9�%l�&�p*�YO�#�� ���:�e���P�hd��H�*�m Uɮ��6��Up�l{�=n4����	�Ne�n?�)}����sO�NT{��7S��2��Ǖ�iZԘ��Y��u��+TJ�\T�KF6�ր{фDX$}&���&Z��D���y	ք���K�f�k!�&j����b۟��
ჟ�Ʌ�^��ϟ�}��gs`��xY\<M�Ddf��B��;�
�
�iu��V�x�hY��1_�q��Q����l���7D���5��%�(��(�j��]Q��o�V󧌃R�� ���1�X{��M�cF����Y�]?�|����kti9AZ���z���j�Aρb)DJ]��H�ͫ���C�������U��.�Ȯ�Z-� 1BRk+0Ŗ�U��H{3Y����"��_���h)��@�d\�%�ͨte��B0d���2B��|���ko>�c����\�ea{����kmh��unKa`�N�m��h^�Ea�[�$�z.Α"KJ�L�T@�ת�g��d�L��zX�ȭ�GG�`#�%�1�����W3�H�p�X���5�A�<EF�����ש\�[�dҨ��4��7����z�3 ��ܿ��=�0��Lm�%,�%v��I��h���1xt�n��AwI��,U��[`�ep�/�: �8�r^	��i a� �O����c�U�T^��>D����9���3����u��w�YS�����`� �=<�r���ߵ\��Q��o���?�}D�pP�:�=�5�7U|���%s�Ԟ�bD�=�Q���O�^�Y&���#5x$������l�?+�W{`�/r��4���:�u�(���Lbd�*H������ٝ��]ٹ��V�	��!���*��R�R?*}�h�{r@Fv!�.�`�3⒦<�z�e���)k��~�M!����1Ng�$'N�إ�`Qt,ӫ�/�N� .�O*�qS�F���e��I;�Uح9V=l.�vk��A���kL
p炇�h6)�/���ŊU?d�4��Xo��D�3�z*�����0�^O��T�-���@�sD����1���@VR�46��_н��|�R�󙛉6�� �)\v�β���J���j���[���:�#Jl��k��//���HX\BʵZ�)����@5A��-	�l+��
!�P˧���D颠VH�y"�Dȹ���x����e�P�0��i�p�`�S�s�{@��fD���j��]�2����K��k8FS�����N��D��`ӐD�2��^�pbns8_N(�d��� :~_G������ljKt<f� ����-�iչ�z5f���ݺ�k=��v(�t���t�BS<�i�q���0Pl5x���zm�]�"�uQq1��{����%��)��	Y�;�d�x3��k!���΢��zpч�P�����[eu �qC�1�����9�~�����1��aĸh��l�L`ێC� ��
�_�fg`�ȋ��?�[�����aŒ�~�+�]��q��
�IP'�a2k�&�X�_��e�`F�u�E!6`�N=;�B�g����� ����X���i">�󈒅9u�̮zՃ�u�<t��9�?z���}t)aY��9�PqbD�<��8X��L��X�`%�5�^N����̜�ҕ� ;?b	�6��%%�)I���R�(�yr�uB�*�-w��8 O�J��[45c��9�%��G����8d���>ݯ�F&�EvݰX0�VZ�;�1,��"�P�,����U�z�<M�<3v| ��G/���$��]��O�h�����(�>�t��~��������4���\ozj6�90�?�H��R��Kn����2?J��L��ч�F3f�s��*�ka���A��հ�V|��h����=��K����\�H1�1��|�v>֋� �[w6ɢ&�/���\?��O���ح\����S�5S������hp�9�I�f��$sB0�� ����3K`��H�V�,v�_H�F�[���d���Z���E(�FPoL�<��aX"��Q��hy� K~��k���;�m�]4�w�m��zLL�s7ǵPF3����'œ�m���[z��{;%;xYlâ��I��V�~nub�i�Q�sd�����}���̮~o��|�9R��Y��m]��5����:vF�u�������l�m�R�EeeF������ Z�̮�)��u�fz�T��U���������9cZ�8�p�1<�4��(W��J ��N�lI?}�-LWdT�@r7't��s�U}�%5:�F�vedm{�f�{{6�!�$�47���h�]mbV�]X�]i���KS�)��a޷���$	�%���S:��ίZi	��iӒ�FBK�_����e>��!SNT��>i�� ∡0e^� ��?!C����6@A�/�j/�*�K2��lV"&1ZB���3�O�g��u��*��>����'a̹��4��Y+�:��n�I379�Lq�ʌ\|�+s軫�A�]�8�D	T�V#�3 L�9"�`��zƌG�]���ot�!��E[v%��2i�}��\�F�`�.����`��d�U�QqM�%6�k���
�]�a�mҽ{�ؼ����Ķ��$�*q)�e��*̔�r�Hk��6;���Lq)Q�
�'XX����nts=�6��*�4��I��EN�M�j��U���?:���A��=df��m!H�������d�;���ǂ�*���+�Qs�/>1�Q�U[D�E��!�����VyR��nmb�WC��ݳ���)�L ���	M��>��1�eMg^�����G��R�AV�D�i��h:��Y�,٭��m��ϱd�5��*�7)� �9�󿓲E�3H���`�VF�	�½fL��<�ܼA��3*#~�S{C�2v��^����G+�F��`��z�DHph̎T�L���3����]Ў��5\��v��Ω��|Ĕ�Ae���l��,�)��`l
�I�\1��*x)�[�_��`[h�u�Y��.�?':��a< ȍMN�T�&£�*E��p�JD�z���.:�T��㇧�"l��pw��j�&u����5�!��[�Y�&��e��8��AEo�h��*�mT0q�Y�5Z�х�$w%����U�EC�l��PK�O9ҝ��}����S��i;����X��l�ȢBq690�dĎ�'�����T<����@�qAk��6�h"A2���E\<�c��k40W��0m�u�BgK�h��=�0�Z93��t�~�"��_<�б�}���{��qn�jY�{?GVk�r׌u ��Ϣ�Dbu
�{v7i���i���;�n�Ѳ@6��Pɓ�tk3x21Mqxd&"H�J�1"�{sd���0�)���ξTT{��>~<Υlդ��o)ȔF/��X����Q�X��t�(ꇱC���V�@���k������PL� �5m���<B\�q�å�fy��3v(cV��1]��8J<?�lw�OЍ���WE�"�����'� ���V��ǰgc7#���ʗ׉c:fE�ow���~�P�YB5u�����5yԝuN/�_�yN����p�(>�F"����A4j�h��a�ìXd�\�w�XЅ�)��~���غ�C
�[��x6��h�����(0MG�_�}P	��7IRb�`����='x �Yu}в�g��,��gf~3^�|:s�H�nT�AR�i-͛�6	���<��JC�7JN��T_��R��Sp��o�ݣ �ފV�2��q>��\�
Fn�o�H<}6|�u�����?���P��j?5?�����_�P�u�o}���m�}?_��a�}n���XE�d�����
~��TP�Jjb#�A�?�3PRc��A����^5���4�OK������0d�<��X�CڂX5`�#���ZU�4�x�#E���q�In���Ų�7�E:O�����wa6�L7 x"�'��O7�s-Y$o��:צ���vH;�4��yd+/��cQ�",��}��b��z��pl�����kA�����5���eK�l��O J!�\�q�l�!���c�O��mv4+@�>�N��\w.\�x̨��kw8ܵ�tl�Aޛ��*;�*d�Ra�6��.��'��a:ޠ¬���!q00���WW�n�4>�e>�ؠW�"{�����
����X*�=���є����Q>㏵q��	���{��]����X�1�F���G������aY��]�y8������������m��a���7�z���+g*�.��A	=���s���Ȓ��G�׆2�|����*��V��������ӧ`�fH|��X���#r�έ�������j_y|@���H�gRط{AI��N��#�4����)��_iQ;U>6=
>��
�W_��D�Sf��y������P\/�t�n�h���8^8B�<O�K�~G�� ��84�&�'�4 �W��ksKc�*�BzE_m�V�N�!\��/�GY�{�v��j<��7?2�D� ����Z:ֱ�ZzX����Jo�0z��w{B�����rI2�����Ӟ��>�=������B���sP!+�TԐ�}��8>;�} �-P��P� ���;cR86PE���S�|�kՓ��}o2�P���f,^5���T��X҉W�EsSWD�Bj�\˵��"$����$�܋���(�8S%a�AO,M��gO+|�A����;�K1���#����bG��G	��>�A	ͨ���UjD����O0�_ѝd�ۜ��%�P��45 �hY�kc�5��j,C��60u�a�G	u��j��
�Du=t�F����r=}�S��YQ�)�A�Z��gt=\_�i��3��n49�^�����*��e��zܧ[����_9(�jf��I~��W�����)�k��#�l�{������|p~,�8��0�����p��Ә�=�[��0m�6�F=����/�w�_ޣ�Q�qp�9��_uy�k�g"��NM�:AW�@�L�ld��_0w�N��)Z�u�ӑ�k��F��#3,�j%/ꐨy*����[�Ŗ��@��8S'J�*������F�$X�����й�Vn��O���\cM�o��t��$�B���c	ۦ*�L4P��T�C�#L*�?#�j/�����������+�Jj7������Jh�����j~�Ѝw����t�}U��)���G���Չۿ�u��y.�{� )���
����-P�����.ǖ�=�z<��2�1$��i�)z�QJ�D�%N��,����`p����5l�ρ^�>}h��[r�Z��4[�W�O�+�Y��J�W���'/&�����f-���̆U޶~���)�!�$HJ���rK��M��W���E����m�d��?�EP���{�^&q��&SWt��Η��@�;^4��ܝHe���zٞ��b<�2�Y�-c��Xh���ۺ�~���6k�(u�z6�q����WQ�8<�aT�Xr��`0;��=�$|%�þ5)� ���S�`�9r�S�e�_�b���[���)A������=/k�ߜ6�}��D���2r�Zꄻ��d�W��<CP����x+)<����@�BN:�4u�ڏ�k�5��⁙��Z�>���"�q�h8N���e&��$ml��y����@���v�v��%!q��Ѩ������r����+�k�|6V06�d�:�$���h�����.��uW����JG�hD�Y��h{�\����v��*�ˁO#>:�S�N%/��' 3�D�D��ˬ��{�=\89��:T �2�p]=�j����4�9�vw�Uч�2�����q�Пc�D���g9|~;��Ok1@O{:��m�I�_C,��|��<�'�����8p�SGq�)��Ŋ]�0/>�:񾚔�qT�{���E���4��#%�Bƭܳd����X�E�*�M���Ќ����9P��M��-֥<\���G�9G�"�W2��z��Tdc'�LC�#{Pe�C�6u���������@�擺�ɨ���fS��G���\	���''�}���ɩ�f\��h��v��Z�)�Bۨ��O���30���1�u��7�F8��،���������B�ّ�N������U�A�˹�p�Y/m�JME��@
5�ctB4�4{���Wkhc�)�_���h�9�5(��������z!���JӖ*�68���td?�k���\]9�?�z�eP8j��
�[G��w
�6��HQհZ?���_G(B� g�!��L���'M�ٗ车զ�s^���+P����-.�� _���,xq;=��eD=��$��y%nUU����@:�k���vh���G��EO���d
�|�w(�D�^��Z��P�.�bf�+�������vU�vئ���?%lth!�fK��9S��j����:�a��L���&�Gxy�e�u�<�v!���~�æ�Ο��r���|�e���&�����Jm�CV������a�jk=�=ё ��<GVܠj:������c��W؜,������^ �sg�S	\�p��&15�?�t����\Y���Q7��͆�L�%�!ٽ@L�X�~x��q��6�O���9E 7hK.hi:�<�̣=���(�����L��Ȳ��^Q&�䲝+�dx>rAFL�菮׻JE[��̈�;!�"��v�\���']z�_�oGm��{U9k�<��9D��7B�._H�&}u�a6��J^#2�~͏O6>uT��E6"�y�ώ�2��ֶ�\|��C�~ťm���O�����n�mW-�M3������ȝ
zTۣޕo�������Z�����JJ�+I~%S�mib4�����F�����u�ة��(v��};��'�0_��Ko����e�7�9��MV��	�E	�|ո��}m���6�t9�6�J���1u!)4���Y���ޔ� }�&�V��D����T�O��3;2r������%�-�����_�B����_��j��e~}qȕ�Y�Rg*w)e���.�2^��]���֎`�eg���J>7~$��Υ�$����$�N�Q���sxG�y<]�Ơ�:�7LŭZˮm$?����i����Bl8�(o���
a~�����I�5Q%��)�E�^�>?�����T�U�k;���Đ��A�w�(X����DK�U��A����h��0oFYu���� B~?Z߿ɢA2K>��p��k��.m�i�����!�`�Ԙ��X�;����Í^%B�������3կD=��7\���\�~���m��R%��{r#,�P�^�D�R�RC���y�e���n�Ί��̇b�M�L�^0���U�hρ]uu������f��qT���|/E��ѐ���O����h�K��]
���I�pL��:�,IE�k�p��`�"h|�����"�_V&�_�eb;�9���v"�ͦ��q۽�鎪y�qG/m��a��+�Qg�e١������QĹ��\lh��Eò-�X6�#1*�����װ( ���M�-#0Tt�r��d���J�6�4���r��/+��1�i�M����� C��e�3��0�j�����Q��糁�k
����#�F�����\�ߥ�+���^^��*#Z������Ey�y:H�D�� #Un��3t��*u��'w�BL:����'X ��`~�=��ؿ%<��J��8_.2�Z�j/$l�]h�P3뢷*��)(�,�4���o�K�h��X]<|T:t%�?��k�d����8j���"�]����ݑ�y����W�H.�Zt;�Ȃ�S���4ˢ|�2 ��m@F�G="��0���eSV&��9�4����3�Ѻs�l�j%%-�4��v��� -v��>�TՀ��=��}���
ڥ��'M��	ŗK<7Q#�8g
�ʱ=�y�N�o �gm�����r�#F����za6l������`��M����g�1��B
q&=��	+�q�<6,-l/0��0W�+|�.T����h&��ZY=�CF��#�b�2��#]6�)e���I����xB���x��-})^�����߄����'Q*��8R�D�N�%�.��?(��)�|��sW� _˝b.�o�(3�Z�L����<�������`�L����:$K�� �&�� O�ʞ��x���N0���<#����U���r�M�Bu��aY�4_�Rj\@�Sx�G-Gb M�<�`��5��u��0�d]R~JQ0f3m1[�2�-��1M(�!2��$��`��r-�զO�ha�{�$X8W½_�5���"͖�u��n��:��W�վ�4�N#��DǗ@�*��iN`���©M�ν\������i�.Q��D$4���~խ����y���Wa���;Xץax9�,ll����<����"���=E��1�7�(0j�.��Y���}E'L��k
H&�WtCm������dL��u{EW��ku�.���	�#�:$M��q ϬZJ���ڃ�zRp�,��b��Q��1��U�2ۭ/SG0�|B#� ޣ'Ҷ.�f��"���/��O{쩑}���_�Of���-�������ަ9��x+H�-Lޠ�h�[pa��Vv ��|(��Ų�Ʌ���FcjU�	F����	���m��&�B�T�: &�������Q{_uh;�_Ҍ��0�E�WZ�7���~�eF)�wu���p����q��Tr2��L[U���#驽���g��v�GND��u�ӭ�y��Z��u�[�T�2�25h��N-�'�<�I]�M���޳��fK��J��8�(8Y�:D�����n$ӕy�8�3Jgń���d����A�q�@�{��aOᔽz�Τ��H�{wa�����L�d�5�ֆ�z�EK C�����#E�Zu�h��x��� �c�����`��ޠS�`pڤ)���"�A�-\����%*����;Տ�3�&r�!���S�%�Eh�F�W13& d9����0w����\}~�p0t����B8-b����e�������C�����f�d�ӃXn���5��L�j*4������ĄVh#�8n䂒ҮU�|kS#��Rj�Ԗ��W�iV�R(��A�,�=�8;�.~�঍A[W�iso���|j@p�Ez�NC��b7�x۰B!����v�i�=���8�����qY0��� ձ� ���h���~R��ӦQ��e��!*c	��"�ca���gl�a�G8��M�"�YQtuAE�+:=��|2�(d�ڤ	Zp<SG�5�SBE�)�	��I0�<x��Ǌ�OLⷄ���?/{�7R�"h�f�	0����� J5�n-���l�,�u�N�\o|}:ط7շ��S�<��"=w�4||�
��%h���O���������'�!5Шp9����?'���e���<%ď��ކG���B[s+g�Kʁ��=k�f�����c"�M��tDH]
v{���6Ԉ��� �}��^�܌����8�ο�e_�R�[��/Nqx�.�l�K���ϡU2���[S���+ojm���B9�`�L�p�~$�Cx6�����W�5bf}TVW�&"T��'�V�TZX��印5#�3���B�Mj΃e� �F���.�ce6�aCRW_�~�Ϫ��=m!5�����Rɀ��Rwf�B�Q�d|���q� �X���!��M��J��{����Imm�"lZ �eC�A�		2y޿U�פ}�\"#m,;��prA�mq��bo�%~��2�n~��dK�U��q-w^�9a�z�K�oS���^�(�������=+���.��4P�G~DSГ�+J�$n�[?*7Szߡ�T�M�j�L䯿e=q��L[��LV�W����}qc~Y�+���?�|/+VI��.v��|���*l�� c4ϑF�$r~��75��T3uD�����EE@����(�pϊT4SIY%ĩN����"�n9�%��#u(�s@E�?�Bj����1�.ɽ��</�)�bB�m8�<W����x�1��?qmO	�\���WZ���K�6F{�7���J��r�V$/�[E���D�5!�q�hm�r=���Lq���%��FPK���G�T<_*Uu�ִ����9��%\����U�?�:�
Q����߲�mc��bE��O�ɟ0�=��pD?d�w:iX�|�	���>����#�!�P�k�LܔȖ��]K�{��/�K�.�Q.�xp�Ƿ�b��bdf���ɢ �u�!��6�7��u���z}�M�]��"�`&u������F�a%K^�"�&��s0��L`�	P��|��3�g���ۀ!6�Fzt�(���F9�3�_��E�g�&
��+"7��9���o�\���z��b�ޱ{Q���$���ʹ�>|� �-����Ϫh�h�p,�˖V�ä=�K�H=���$�L�GL$k"_W�Y��&��z>zP����X�`Ew��N:��ͨ�ը�;�����K������'�D��▻��	��R,�dn�m�d��=��
���j?e�fPz���~(hSO/�����^��uD���^��~�-��ǝ��Y.�=��BSK�%���Ki��sF����K_Z�$ �] P�~��(��l�ݐ�#��c�t����5FW�Go|�D�U�,ݛ�?���Zu��9���g �Ao�" <`���^�1�h=P\R����J����N����>S��c]<v����mk����Ƴ�����ʡ�^d��A���7�څH��\���^�����d�\�E������j ֑{F�M�g�.n��A� ���̰��q�gsn�4�;��̩>1RH}E�ퟫZxd�q;DՖ~r�rO�|gn��<�_D�9�[���o(��<+���& �Q���s�~7�g���
s�EZ��s�B~ YƄ�^f����g<�G�g�?�gݪ���;2�J=�*���
6~��ó��;��UfER3Z<^"�����`����h�Ѧ�YdA0L��0�Īƌ�(M���[�ք7p���~���GZ5R����,V��7���\�\���z$������S�=�`><}]m��OM&o����b���N<�����Kmx⪼~M�	��/"ό��GXW����[L��W�aW�C��F�'�L�6�g1�]F���ҭ���۪�ч���9��
�q��_�*�L^:��$�$�Љa�K�E+���&�]h.jl>��oä͊�j~!W��DO�w#���u�����Y��){����dT�p���_#8d���X�E@�r$0�h�O̖@�H�iP27%y��K��J^;ڎ��:d�!Im�������eם�Z*Y`��I�a�_B��|fۃ(]r����p��F�X���au����:���}�O9)֛&ڰmD����89���I��6�ǖ���㓗�����D��E�wf��t�o���Mpe�L/����E��mf�T��%��f���0��KQ�~>e}MН.��2���ϟ7����iQ��4�^��ZŊ 8@�'�RR�1ۓw=K�|��g�_�W-��Z�y�&�)K+��p�i�Dz�%�	h�9�,:�͌ޅ�����Y�f��!V��$/�Z0
]Ѥ�q|��p��<�Pvd����dof�{!��;�ډ�E�i���k�!7E�^s&}������S�4���+x;��:��9xtdv;(q�K��u�A�N%���Ԩ�r�]�I�3\���ي���O�ڬ� -藘Z�q�3^��T,��o���y�*��xK#yD��J��S�#��X���-�*7�'<w�M�R�ܠ��R1I��n�h2|@�dE�׎�w�F�'�C��䥇���e�Xr��.69��=x;5X��$u�(qeA���P�ߍ�Ek��4
!ߔ�i�KQv��c0�U~ս~?����5.�&AܤC�δ��\�r��慜���.�r��;~��I��!�6�w�)Ú��Eo!c���̬Ř`���w�P�P���)���*@�*���,%�{4�����x�klO�m�~��T�1���aL��v$!��z�0���'��@�AX�	c�g��K�Ϗ�<	���5[	�pV�����:�/�k�����O��+3��K��anLv�6='"��r74\�`����'��~��tpR���W �/ta�T��Pi��=6�~̀�
���/GG� ."eQt�	Nt���`Ē��.���
�%,�=��h@������'H������������u�S������[1MR����8}��R>GE��]9գY��͜��kvI������GI��Q�<�܁CÃ��:E4~u���ZPj��Ƒ?��2��<�~�W5�F_ux�{�+�-�$��
	�p�7�S��j�������j
�,�i��kr캧yLK/X*[1�u���C�{˟�ܙ�����{����4%�&���8]��&(jbh=�����	�>�w�=nN�=P����9}�#%�����\�t,F�=g�le�	��然���Z^T�)Y&1�)���ܛ&H�h ���?Mk-m�D�WIwB(��^r����4�����4k~��Vc>_GPɑcO�C����ha�%E���ͻa��hC���b?i�G��/�U�vP\����3����O0�ax�������$XL�#�y�T���^|���@���1����C1T�{�_��m�яP%����
B��r�Y]���O�ٽ�شڎ�bg����݄�RG��'#�>�����i���m�\�;q>��Q�j�9�����`m��o�[	HV%��7�$�䟭`+Y��8��0��ekJ릓�;���u2�R/>w�)�u'���f0��F9b\�^V��G?���MNT_���!���U	X����u@����;(�K���;�Ǽ�d�bBqMB��4�`�>a���Ԡ{�]6��pۃU1����Y�DY�W�ɒ~g�<!JQD٫ɺHL:� ����k=i���H�>x������a��ENbJQ���R��{�pV�OLa�����R�8�+�"��;�#x�GL 
���@#�jZ�u"Q��<��&���| �E$�U�.�R��6�"�v�����^��'�/"D�;�$iCw���R֖��i���S��V*R�Rm�@�	Ԏ��/����x!��]󪒰X����<�=�	�̽��f+,3M����y�'�(9'6L�E��q�|Y�#�V��xv�������O=���-�NF}@'ӈē�ɋ���p�皛�ٺ����������_����#�6΂C��
-���,��CD��@o��.�Y�T��{YXv�����Ѝ�"���������WW4�!���Jr��+���`��=
T ��J>m�Q�E
�,�i^I��5.b��R�o��	V�[�rP�)���lk.)�}�s�˗�Zb}��;7%�}�HE�!?y/��jo�8����Ȣ՚����*�A�aWs���{k򼇘��A�����a.J[�Z�/ZX8n���Z&���2@R����vU]����>�c���V�e�g��k)�������6U.�J��W��9���ER(�͞�����2x޸H������^R���aKd�[�|:Ü�`��s&M�j��e�]j��cxZ_�*\ci�ޛ����T�>�'I� ������B릅���S�a�i)�j�+�n&�
.��o5��y���$̆�� ⸒0}�;ol�����S�4�գ�nK�CZ�9m��K�CE$����DBk�ӿ=����Z��"�M(b�c1�N�hPS��i-�3(�(��� �p��l���OEs�`X��t�'&���\�� y�`H������"����y<��QC��^�^�͆b�g1��8�~�A,V*�S���1�Ayw��|L����ܭ�π�m~ڟ�Q��!{�%#�LdN�rW�Zhә6�t���e��p���nu)��p��V���!SxM(� ?i!�#w�����[�P����"C�N�s��la\�`bx���i��������{v�Ի]$�"Dp�P���׷�N(�c�l�Gk,Z˄-I�D��nJ؃6w��B�WIӛ�Ǌ	f����9ʊ����6�`���2��99
J{�%���؍����N�TZ'bbOs�Q�,�|�t��E�Ɛ�yu�F��C�!ӄ"1�n�?��Ng߉57��-7��Y��m�+�3ﯖJ~/��_�G!��e�}����O��%�w�~���S��Q�ęvy��ۗ�6�z�Hޭ����,�}��f�8H|]FB��=~��1p�{���ɨBx���i�`����^�]��o��c�1���٦�b�WޓL�(���׆��I�9` �Kd���BC� �<h��ruM=�]���QDj����tiB��,UV;�?��3	:��+� n��WA�#�y	�(X[u��m!�6�$������nY2ێ�����RA�Xd�/�� v��5� /%�n?�u(g��t|�|7M`�1����o"λ��;�ʸ@�ϩo-�8�+[�6���
�K��-���$��C��� "A��jjЮ��	(*DP��+��5�w�҅h8e^Я�a�[�*<ΈD	��̋Y|׹�#�$��� ��s��(�x�^��k\s��]�c��r'ca�myj���H�#0��yE��J��fy*tb�=��bpe�����yW3��z�Z)��)@'�3�'{Fr�����5Ix�(�A�P�Y��{��-��%B��;AlD������s�g�k�ԛ�m��K��E��n�.B8�S<�&ߔ�4��=ȸ�m��%��#F����*��s϶k�^A��D^E��Kc��,:i��>��&G�M���������g�ڋ�Ѷ��G&~���,3H��!|O���Z�D���� -e������&�X�n%��i�W���O�1�tt&c���L�2^�\?��؍Fr�n�ťt� �_�3מڏ\#��?�ry��	m�D�ԑ~���H��{��r?����le阥���g�Mh��y�C���Ɨ���<
�r$��;�n�b��(�̧\(7w�5���Fm�M��������/������Q�
f qE�*	Ez_�lh���t{z�d�uas��RJ�1(gT�IپYϑ�p�307}̌��Gc�խ�S����|�"��2�Y'��=R�v��7k��dI��� ^��^����V����w�0�+�|�g8AJ�e�'If��c��h�*��+����)&���nZk)�أ:fZ��Ւ5Pm+�:��B���5s��'s-Si/�U�L��({%9��f�] ��׼��a�uW6:O�>06��{���(�d�`o�ܺK� )r�C�Ж��`�)|rYc�|ۢ�}|�Q@E�SS�\���0�c6(b���#��x�<S���R�&��e�&Drl�<b1:!�NȾ������Gk�����+U▵ğ��׾���F�w��A���:+�	�r�Տ��n���	4h���LZ9O��1���yHN�ߙ��~&�RN4�0�y���� �5������LQ�<W�|�Ko��/�Ї ��ˊC��R" ���"�y@y{�S8,��uC��
�������-~�8J9���mm��4�M�'g�@횂��>\����]�K���ڄC���N0�_4��"��9���/��[``�n<x1#�T��J�/��g�

���D|N�BÜ���?��A4��Md�<����̺7n+��ݣ�"d)�1�@1�j\j-��0��5;��8WoVd�N�E[���6d� <�J�K�YG7��7(�k��b}M�W��,���������9�n_j�|D�-/��W{���E�_�"������8�y�9h�� 7$7ߚ��Җ��YE���k��w�I F~���Q�[����71=�m�h����8��?�[����?��I^�?�C����"�����/%�!�r�� <�{w�����%t^o��gfՇ���}ɥ�� y9fD���3�	����͜LP�]`��`�~��GO�;%LCA���B��6��Z^�*4�L|.c����^ⷝDv�@�
�	��B�d��͖��|��>{����L�vF�����2e�zU(��HO�#�(��VB;��>Sc?	Pt��E�C�Ǵ��f��fGd�\�|��y����Ln���C>����YDu��|���b��ɻ��i�]>�1X]�t�5 `�{�tq��7���y,��ؖKқ9���&�+���P��}�bHs��!���̹�Љ%$�Y��W���������Gj��LqhHw���NC:�R�_�暒�O(�*}�f�A�cU:��SL<M�ꧻ�Z���$���48z�fH��v%�(.�uQM��2�����Ɋ=`�]��8.	A��G�/�l�[�����#��f�d�]��J��3,oǤ�K�0Ft:���d�(�r�Ã&�������b}���K�|z	�Z���:�ì!��"�>�\�n�2ए�q�vʞZ���0ig{�$��좋�W=B#��0��o��(��~~t��IB�g=S4�Y;��G��O&��َ-_:�"�=/�ɚ���m��5ﯮS�U $�˩v�2$��R/g��Æ���=<�
���"�����k�!�&��u�V��|촃�@��W/=%���mg$Ga�#�e(E��u��Q��8}��^���U[r�<��?�{���a"�r���I���9XV��b��)M,��1�a��X��At�b�F ��!d�� P�Q�r��u�V�B�Oٜ���SKun�����Q������8�Fp�y�h˳�?����8=�e���c9 �w��.B�Q���?�0ć�!�{��']���/���>�[��p:�9٨��іQ.���2;O���%7Ou�T%��R��7��'�Ѝ����������]'y����ȱ�W�F�3��b้Rq���pT@?���]�R�W��������xg�%�+#�e1����v:4�}Qx����������}��x޺��x����84S���H��z�ׇ��X����'rH�t!���uȑʧʷ�Ѯ�{���G*^���-$&����geL O^oK�෬�{˓�ёLcc�$F9ک��/���'���λ>������e2�v���;����L!�H��h�[�� ~Z5���}����yI�F1���3���^ev���9l�D������Հ�1*���e�P���~�þ�t��|$e=F,J�1�I.�nZ����C����.S-o.����U�R�w��¥@[�����]���cI��jIw�]=��4,!2�ť�c>\�6P����.ެ��(f`�4x����Z9�]��?/KSG��o�ͅmJ1�� P�tZ���&|��Q�t���[z*�%�\x��{����(V/��9
1��[���K��4I�۽6�7\�U�����X����QE�'с��*�5����|nh`�&��Ӣp������"�p�Jr����P}�dhɖ����޿��$���x�Ԛ�6@�D��X�Fz9{�(9'!|�ͿÞt���j��a_^o��`�eW���֕�h�!*_�Pi�����Bsr�+W%V� β��gl1������0Z3p�M�㪆����g��o)�⼐�>ټ���.Y�{�}7yQȾm�G	�x����tp��O����"a�0PU��¶K�7���k�oe ZQ"N6������^��A��/���<��,賣/�H<�
:tf�+^�����i��	�<����J��`��ޯ��|H��X<����v,g�f��j���Nr}D��gt�+��@ur��*���<��*� M�#a�4U�݆����|SH��	�E�=�B��h��M���Q�%v�Po�k�N�8:L2��S��₂r�&��1Ј*ۃ�4�R,�&�|A�WP�M��^֥݉�F)��h�a���<<D��'�8��"���D�w�V����4?
�=�=�(�Q�u���Y���j�����X�H�i�����ǖ:;��0�\X�~@j��w*���:�q�r�D��H����^"}��|� @��F�*���;<�t:W	` N�Y��U_�+����V�q�#d�B��4}�ZD�^�U�侦�(��s�;���r�y���k��Dt*Q�G�2ega_w��DG�?�w=>��۸��x(x�-�c㥔W൥��$l/�֚��l����o�
T}n Qدy}���u}��q���Q2�-�럵2/4抷�RЩ#iq�l��1/�b�	�2����*v3%��aM�
�f�ő�IP���zg�T>��:�4:��&N�,1���ͥ��}�W)��?��@{ۊt,��r"0�Ob��f��z���[:�l�G����_j��܉�H����r�*�_�oc��k��?���Ǖ�K�E���Qy	+l��7}>��so�%�p8l_��m;LQbBx��jt2G\�'kw�b,OJD.T�Ę�|_���U��U&�����Y�na{�r�˗9cC5;��۲�Ё_	�Q��in� M���Z��$����*!6���"�� ��U??�qw����.�PwE�u��2iI*�?�+r��Y	F�\{U��䥮�<��82o���g�s�4���#/s����CX��HA��d{v:<�S)?��-��"�>����f�P�n��wE�m;V���_�3���w�?��UWpi��`Q��H�|KF��TU��2�]�~bς^��&߶bX$����;���!4kf��5��F�rB��g@��zH` ��╹�k�p��2Ա��-���A��P!H�-�εE�������v��:�n��I�l	�03F�����>��(3[O���$d��������L�2'U�7�~pХf��\�/�M�0 A�[��,�r�ʋ_�H*jZeΧx`X��U�>K�֥��,�m�e���Ĭ���9q ��%N�~r�c�f'��7k��������k�/������up��ˊC���uR0%���l��1|�z�Kˉ�!}�y�C�f�9�s�I�HX%���̪��t�"�ˮo��M�d-�>W��h�Hj?�xp��@��_
�c���A���=�O�9�B_�m�B����#{�}i�@�+%������ �&�i\�x�9�(�|��$��9���'6 �U���JS�[�ܠ'��k�VEF6�kחϪ��؂�N�	�$��[�n���BrG�O߿�1�
ٞB�Hf��<!�ߝ����S�A�@������IT��1$!�9�8x�$IP��J'����{�Z��<7P�T~�@G��m�gy��U���)��޶�8��&k,���;*�vի:�"e䚵�쥄�Mǽ_O��� ��"m����R�Cuf��=�wم�%��Pg�R����^�������T�|�l"tN���,�����B�?��o���Q���ެ& ���A���+m�����,e�@7ip�Wⓝm�n��F���n]_G:{����0-�wSd�C�sLU)~�e	��H?(���3�l���Eo8o�}M���c�b�Q��xs�+6aq�k�9�]s3��~`�y���QǪ�s�=�K��"�ņ�N��&:P�#�R����Ԙ�����Y�ȚQ�,{�k��!�5�	5MiX>��ħML�߳"-���ҳ�����kw�R҂�Q�?�+�85p&�����ti�!���� -��Y�O��~vs��ke��lk��P��T-0L���;T�J�V���OԀ.~�ɜ�a���禃�b!��Jr�q��	q��;�%��$Pq4��^X������e�#˦��J�8ϴ��slu�6g���R˴�vxۆؒ҃h���1D\WtM�ЮmT��d�~�������%sẉ;�g������0�!�m�$�m�����ȸ���j�+����ee�n�����2��؞�"Z��w��Y����Cל�ؒ�D󭽆�lZ����Csl,���ܝ�ԡ����S�~w�;a�����1���� o�n�@�ڣeb��/�W�����E��[	��1�i�}2op[�<s��3��i fv�}_��)���i�T&:����0�u-�_?����At�)ˆ��3{��k�R,��Z�2�U3�	� ���>;
���=]�w��
#��%YN�:�.�DPd �NJ1o�Y�E䵬YK���nƵ�DI��W��׉����ӿaB�]Mr󽯒T&(ު��
r��/ɍU���+���ܻ>0��L��%B��T0�?ce�>Q�?�P���0qi|>����`�L��Rr�9�Aj|�-�ܳՂmR�w7�/�������;��y�j)��G8E�c�?�HLn�y���N�<�Q��.�BZ
c.1��򶞈��&�m���ҟQ^��s�g��jT?�::�p*�ȏo7�5����PP2��P�u[�xU�BX���g�0�S��̄.n)�����T�?��t��k]�,md�������h^�Bou����U���%=vf��eQS�����휫��4� O��SUHW,�9�oRDXYtL�0ߨ�K0:��z$X�ZQ��wVqxz��?�~}�@]o-����9�z#����"_��Ө�@�~V�گ�d}"bA����x%C(��*��Vv�O�,�0-�6�H!�#�gh18��5Ϧ��B�8�_��[�i��E�I*eR�v��-����ھuR%k������Ei�岘BC*�ҬO�|����*m���m�wr96>����
r+\�����z�#�>5H0�F�/��v8Ip�P~X��$d�/(&Z�>À?�Zh�sQB�[�*u���$q�tN}+��o�kﮋ��@�tU �y1�L��S��J��*
pA倬y�
dvf������OCQ#�A�>�軫�B��_�j����M`�O�]��(��\��bܿ����/�S�xdCN$��UJ�l{���N"_�f��F
�������G����e�m��˷�8��]Ć���a@�B�[���q�}(�E�ߨ*�w5����O}���Y���4{
L��W|9��v�Sc��t��p>�^���W>�?s�����PL�p�\}�/t ��ݝ��G���ҎC�NB�E���x͕���cn�>Ɇ�_}�N碗(���%W7#�P��u�-8�M�I�CA/Q����/kD����"W�y*�tK��-U��,C���ċ0WGha$'_w���#����Z�5 �y/L��*��M���+j ���:�����`�_镚��O��e�7�{D��3KF�Zt^�F��܁����!�����Ą��N��Cfm>:#[��p ��W�<����Ɖj��z�(�^s@�˲	kD�0�I4ݸu�St'���cV������&SGoZ��-��)������kk�����T��"УQ��dF������� Q�h��;�MH/�\�#�Lj�՗#���UF��j���g��m��t�Jt��;W��F[��v	n��D�;��##kQw��b0��C2�e�ԺW�2�U��#�{��H�Æ�%�Mh���z�?k��#y��8/'��z�ޑ�Q��`)�t����JgV�W��X�r���5�o�����e��pZy�1t�W�D$;��� �ą�ʁd�u�ry��MM���o��㭛�<����bV!Р��¥8�d�92ë�kw���X<��Oc�3�3=��
D�ZWi�^b�YdZ��%!�5�[�
�Q+�����߉����vaXe5S��7�E%��^��-��0��xY�0���Q|���d���NߓX|*�3���\<�X��wT�';L	C���J�cf�����틮h��+�3�7r�����^��ե���DMt0�  ���M4z���o�6���F��+���(���iqx�>��Ʈ�u4F51{�Q`0L�l�Fz�X3e�o����Đ�_���֤CItj�Q@�NZ,��V�w��Ŀ�o��0]�	��C˝��bN$Q�ݡ�[@�k���'��a�"ɽPD~����y@>��N��Ȯ$S	�?�u�
�ޘ!�/���� 1בϞ��U���.}*��F���)2KzS���ɼͨ�M��J6�=tF�76�;#�X���O�`��O�2��7�A��pBYˣq�SlTӵV�/�d�_+0�"�Zҹ_)����W��SH��d��}�w�	�R: �9�;��0穯DYA[���Wt)�4�����;0Б�l�?_F`��|�I��<H�U��SU�-ټ%�Om軝q��� ����+)�ǖ�n-����|�w���_*bţ8yw.T�CC��-:=f���:b'��i2����"���z�n6�������}�z6t��)p�V�T�Q	�ݑ��!9һ3��K�a.xE�2Sz��l�j ��I���+ ��v�3�ξ������&a~�1���oTv��%�)��LB����L羒v:�⭛C��h�%x�K���82|{�F��O��:k�?R���l�R��V�;/T�(�T������!c��miw���1O��֩p��)n���G�Ù��<G'gu
�������ŵ�Z�����s�/ Bc�[՘�����;Y�	TwXt�Ɣ�7���8ǣjg���,�'n��4�'q�T.�]
uQ�F��u _������2.UK(S��MQ�d텡^�l��f;P�n.��x$��h�J�V8�� �9wΤ��I�r�e�q�W���,��uj�"gY�
��$h���v�l�ɖ��r�L�C�a7������>����h�ΫΜpM:$ʚ�^�<�#�Ԑ"�|^�^�FR��m��K�]��a�/O����꽷����4���8��mk�x-9m�+��ܦ$xs.Gl(��	���*�o��\n���k*7�3�"��#���LD���e��C��o��vE��a,�p�-ֳj�XX������d���Oё�͓E_��8�e�V�	�������v.fƁ�� A��d3��9��wi1!3�:�)��$�%�����K��}	N��Ǝ#���, �B��v)$l�з�nM�ƛ��t�z�V?a#v��Õ/��b�+��뉲�[./���8�;���ŭ������YSQ.�b���w������I�=iƄ͙\��B'9�������_�,�H�U�������7J
�8q�F\-du�R�)А6�8;�X�QV���kx*���I���E��_�� �x��3xο9��P�&z��1,u��
b�bP��4=AJpt�0��g����lM� ~2H2n�Y��;�u���u�SD?t��C��C�c Р-@�"�$�k"�w�F��9J�'{�*���tQ���}�����jB79��_���,a���sŜ�r\x��Qs�p����r9뱳������{S@�z �ō�g�Ӗ7$�9EM���jhR��c��O���\���h[�(�#O�{iK�G�g�c�"b����q��9z;K�;^#s�ͳ�\�N���v���MG� ��R8q��K�/�l��יL7���հA#Sv�4��D��i�ޗ;�����o7�e�[`�j ���$q�B�Y�x��j̽p�ђ�f,]i���~�AY�oM������P�I��[�暔;���������v�'�92�����0�Kd��iF�9�� "D���ʹ9����R�#6���������c̈́C/�	�2�ur:�II32i�F˹���\@�ֻ���GUE ���mw\���b!�-� 	��mw��a� u������)F�-N��"W0ަ3�bki�K��t��>[Y"O�SR��s/H�D����)��L���T��0	�5_���4sQUv#�/��k�qpC�ڎQx\M��a�>D�b��
�U䡲�Q	��3������Cg��8�� �{x��'�I� �ݚ H��a��"�f|����`���9	bdS���t4����p�P�rڝ(�2���YnuQ�+��'�
A�ߠ7V,Y�v���۞t���=��jq��6�2���yd�l���R�?�������ML���ܢ[�)*�����0��-����Z#�dY߃�������{�J%bQ_�8㛬%4s�<��t�$R-�A�[���P��TU2r4ܵ(k_��JdK����>����{sS�`��6���8rnU��T�Zƶ"�4\��R�4C�>�ir�f��ʝ,�{O�ޏ5ZA��孩)�%_a�i���v)6�����9��.s��-;ec|�Z�o�b���>�{��q�*3p����	��]�#�����
=���ms}��l|!*����>�o��Ѯ��fQ��� ��tX�F�hKS�l��L��np!;SH�<��{�n�e�8���4�X?�0��ZlVr��H���/[�O�J�q-�CO��
�m�4}u�Ȝ��cOe�X*Y�{�`c3ܘ�~��=���	���!�#o��V璃���
	��� R���t�L6&c�:d�v���i�u�%�j�<��{�Ms<������4$����R�$ �{���
���w�Ɩ��*�`���N_���:�MV�a���p}�����'7tHL�[�<��T]�ALexak廸å�����l�/%*�-c�(@Ȫ�a�a
��W!(��v�d*i����w���R��Ԋ7�R�,�r�W ��T M���5��G�^?HX��?*v�q�����)� Z�QV(N���  �N�FH����2@�`�?%+O�~901}s��EL��m�]J��/	�.L��97���i��h�� A�p�m)�׽�Ь�����A[�.mT�X�i��Ej�V��pDT<�-�xٌg�Ko��N�yB�EqH���ҫ�-�����ȫ3�_?}�9�(N���ݣ��h�	B �qn�k
��>8�k�����?H}��j�ˤ_��oa�{�s
e� 0�\�?��.iM��}ZN�"��1p����%]�H0e!>?� L��{��A	C�Bɽ�֏�=�=qc��h��g�K/��h(�c�����>��o)ʡ1+�Zǅ&������k���A5�h���I
��7�񗏻<<u���O �ҝ���@�|e:�	�$� �$�pL�G�L����l��������k���53���K7-@�d�����}�2��X
#������5{v��>3}J"�A?��~�e�[A?g婭���6�J� aL��u�uV"kg�_7�7���,���<�pJ�D��V��$�"��/
)�U�S.A]a������Pܝ�Ͽ�_X��KK��cѻ��Fsi��\l �d~έ��v��ʅ�	�3���PĹ�M{
d��ڡ�������O�c�횢O��`V��1�|�~}^:��ώ9t�wL@��u�}Nw!׌s�f�徠�TE^��B��SV g�n�u�g# �]��f���c���nw�^�5%5�g_���6�79��V�(������B��D6���Ȝ���F�Ɗ���A�>����C��lL@����"Uq	4���)���V��"�v9guG�ej��e�qn��2)��%>�D�f�#�)���#����u�:������Ǻ��.�_�Gۻ�@K7��6��[���L s��N	�|�T�f�p~�^�g?(�_塉��4WNy��U,#pV���m�b����������
V�g_�X���%F�%.�Vv�iB�{�p����+\���93�Ey4wmfN�~����z�^[>m��60��Y�<>O\uv^�ú�ˍ?F�n�M�� � �<�mc;�2�u=)��>=��;@�qV3Q�9w����^���G�8�YX��/n��K��#�!6c<|�ΎWџ�j����h�s"ɫu�	�&
�����Ϗ�5Łe#��n�\������C]�PL]U�wid]�F:�@�]hqV��T�6��h�Hd��-��ܓ��I���p_<&�J\b�K���K1{ʎn�m�w�wN_��T�9�V18��E��@�2����u�e��;�$@��Jfk>�˩� ����jV������$� &� �r�ed�<�+���8�*I_M�x����S\h@�3)Vb�`�����)�����A��K�9_���~I�C_�f�`I�.�M�x@�!��薚g��M;����!%w`3��w�=�[]�uI�8-���G�LX��������V}���}q
�o�q�����g�K���j`��p��e����S"岩��
�\@�*_���$�߅t���5��$�j��Z
����?:��;֯K����3�q�˄@5^o08�*� 
��J֡��=����VPd۩�+βW�B���Д�6R/��5�k�C"��p:�ΰ����kY��fv���Ox�c�!7�-�u5��٨3~��P !қ�Z��}"
85&9���j�w�u3¹2��r94��-�r�b��Y���"ԙB�`�ԛ�	^ƟW�ݑv��㥭+�'�Xܹ
Ly��$/TO�����F�iףp��h�_-S6 *�v��\
6�Tx�F	ro��	���K�-��)	GF�~�
��q6��A��_)�^�?Y.~��pLʘ^���1�)fQ1�b��;I|N���ԛ����)G*�G��P���ǅ�g��J�'#)x����P��Do"�'��gĶI0b��Q������*,fx�1�~c�a�T4\��' ��R���+��U}D(j�Z6 d�}����=�u��q��5x��Ҙ�~$n ���-�+>m���h֋�I�a�W����Bkl�Nר���e�5�5��ǇU�es��8�����?n%"v`5�����y���)lY	�por􊫽�P�#�=�S�>�P����Ǭ�	g���ć��6��2����t�ԛ�:�m2&պ�_f9��,��g�g���ft����,c1�\W�������otY�g|����d�̗�OV��ev 	�rR����G�l[XR�놁��95ð(	^U���9��V1�4n�?�lx�����F���?n��QG�����?���ܧ�e���^�������g��?�l���88s�aò-iJ���l�B}�̜�� ��7���s��,n@P��pM4��H���>�}��ˇ8>�p���Q�Z��5�|7��
�D��c�N�xԐ�W%O/ƪ��唚� :��GtP�Y���h{�f]f�~��+u.=)G(�Y������������N㧹�rϝ��Q	������4�
?�i��s�����R�X#P��o^K܊�nDs�V�Lt�=��� M����S^'x��a�gr\�qE�hnxk��KT��pn����f&{���G �'{�l����L~�ha�,�x^:9�v�H Bx�h�A���w�%�b�my�����Jv_K��+�����fVc+�=b�0V�a\��Q6�F���hH#m�H����G}����<���G�b'2����Q����G� �t�z��&��7����~��q����es��ြ����3���G)�����
c�?{�af���%�>��Y�����ލ���6Q����^k�-�\'�	�D��{�����`��F���0<��U�fvH�J���W.Z�8�q�����Ν��}�`[@>|=��j.�&�L�>_���4��*j��9�8� �p�5>���A��J��j����S��}�ib����+=m�ut�4-.�����12�(�=u�CS�@/ͼ���ȕoT���ެ�'1��'�q����kQI�,����?8$������?��?T�0��JF>���)6&�<��A��;𱪒U^�:#9尿�FG0f���ڢ�9%R�A!]aD���V*c��i�X�L�H�26�~�2ki�����?��2G@���n�u�Yю���y��� �&@���1�-�ϱo-�g־��=��j���ʚ��c��]��Xb6����sF��E�/!PX��sVu1
�|�����*Jk���V�H���+�;^D��y�"��'�tR%I�wC
-�S�x�Zmj6N#��p)�i�g�@����N|�R��u(Ƅ����+nXm�WSO��cL$ۉ0��"B�\F�tpc�tt�o.�b�18�8r*�
9l�d�Ѥ�d"xX�uU0�w�́�b�&?�豸�<�9U�Rx뇯������?.�Qrs��A��Z�wu�y�Bѽ�:���'F�C��d;f���hgQ�}���H��*����!B��H��s��.g@��/�ʾY;�C�l�hr���������z��A1`��Y`�-����lߥF-Wa�$���0���QfK��"��0�C�!PD�k��}F�M5]�H�_��ȿ��ҍ4H4�c֊Zo���vK5�VF�����>��Z+sJ���$-X(���Ϙ��P��j�s޴u�1B\��O�!E�~�+1����@��ȡ��\������n�������{�bN��R"��	k��w��WGD�	j����?0ʙ��ճ��W#f��ޟ9�}DC6y�q��A�jfӝ�FEoо!�]:$�~�f��$'�0d�� "��A����n�72��x�<3A��w$gҢ��Wn;�,,�X��f7�WDcx��[�R�=��A����l9�mE�F^C��os��ac�䚑��xkd��o6�v��hW�1+̧������r\�ro�0�{օé;�)�댡`,~��"������HNgL���G�!��c�=��&鬱��,��o�e�S�,Js���2R�1D]�G Y�j�4p�������4K;�)&ă���!Q�!�����C�J�A�p%T�Mx�H�0&�l=	q�_L4|�����=gO��ScSа8��Zђ!�5�T+���4�����CW�7�!����rw���P��?#���r=�B��Aȿ-2p9%Y
���%
eV��#
��	V��M���{��]�w�li�qJ���,>����0��к�ܷt��s���˭�$�=w�uI�}�(���_x~�.[���&�g���nvSK=:���E��$�-�u�q��|�x%l��R����T<W�����}.ݧ	���W��'
Q˾��ݟ��#yv�im��|��8Y��JD�*[���`�֕a�:�2Dg��������ivP�f���Jg���gh��ȥR3W'�zo&ݔax�\��P����B��p�*z+�G���x�����jQ9m�|�ɵ�]�Ez;� Fd��>2��r�����Ɉ=�Ȩe<��\��ĝH$)������m�Q�# �Ǖ��t���/7:�Ғh[�ֆ�i�:�I�jFN��P_.F��ոA�L��:�%��g�Y0S��m��Gy�y�H�yZ�n�|kΈ�vw�a>z,PB7�g���'3'�{م��!to���Wk��N*d�r���?Z�������Y7DH}����9_`:� wo��ߝ��R��m��2����D�$����ZB}2@f��k�\\uԢ���E�rM�N�Ui2�a������Y��sW��8E��(�����?�g��pxz�-����V :�~��>����4J��h0�͔�Tj�ڒ�XQ�iZf8��v��T@�'�\t�d+�����iv�.���i`�cܘ92�$�ȥ��5=�A�9[|l�a�6���t[�\su�~�����SCj0�Ut3[��(�f�3������p����S�+J��,۳�j�'n�cn��:���)E�Tː�.���v���GWEU���!WX��y�a�ɗ��-��I������?%�$,o<o�f=ׂ�����c%�E`Z�R�ٕ�g$��g���lz�UN��)^4���;N�Mv!��E�:%J?LcZ�������0�D(<G
�>K$�Ö��*����0IJ]�	��ww��JP�����Z~*Q��Z5Ol���+F�@���;JѸ�=jId��K#�aa$��tg����DLY�j�>p�Ј�����Y�8�0܏r�b��z5;��o�Zk��I:~+zīV��,��%E���~Y˔Pa�+֖���4��s��1�IB�K~����^�6e��sJg�����y�	Y"9clG=�7�4��� }F1����D5�m�|}P����E����Q�j
�ܲ���z�TT6��w�rS����k/l"��J!o�Y�^����bA��E����e�����껱����8��"��_�q��*"�U%�0,/����A�d�$��̌7�eFn�ء&6���R�#N=�[���X��l�i�p�E��V5$l&K��W6�$p���k�DfP���*{�j4#G�#��c���ӁC`�mA��Є6]��u�#�����T�!�NC�s��dM̗% ��V��-.�f�1F�z��QiF�C�=\��f]$��˻���+��,B�I5@���(�;���\�7x*��P�ldBᯮ�my��!�@��E���k�j�3;D`��󆤝R�li�%�\�䙣��Ǽl���DFbE��!�5�U�J�f�}�ԫ�;uݦ�r�=`�E�ld��Q8����Iv��x��\�b��-�'n��\��q/(�0O���5��\s��#��?9y��OJZ�Nf�}Dﾇ���5�Mh�-uK"�]��A<��,�+hJ�cr��y�Tu��$��d���ku����tq�9���9�Zu9�~��JD��r�J�0w>�Gӧ���e�K��f
WN�@���:�(�~m85��#"B���xnĹ�d��b{��v
m^�#�C�V������ѠG�Gt'����Y�7Z*:��7����gH�$9W}��l��H0 N�˸���jt�*��P��w��ή�Ұ��Ϯ�-2N����ތ@r����_�ߞlԹES��;h~��ʜ�*���'�U���c h�:�A�1���? fO�/u�G|EK>Y���Ыh�߽�ϩ��%�)���P��?��G�9�o�`�rO[�
b�<0��܄��(Ȕ���vFc%��Ő�r��S��K�X��n�t@�>��ĶG��2��3jy�*@E�����DS�J�CB�c��l��F���0?��5�Aoc�"0�cל��9�YXZ���� X�������+3�8Qe�as���61��LKg�e�@�Ֆ�����)P!��v��H�!2�p���F��D��q�+$�WFe��NV�.���:��a������}�]�!n��]�p���]��<�o���a���׏�o����G���.j6xf��e`
��&�sE��+�Y��[�yG�T�ӱ�
W���[?�|A���T���iڸ��1���!��]׊p�~ͤ�j�ϭ�?u�T�E}��a��S"�N�^�%���9����fn��F�	��|���?2�ܯ.�Ә��m1�������'.���47.7b�I������!)�m09�S.'ģ�����uYl}�{����T	��J�?��+.���㷡B�ȯ�pp)3�:���m| }J�o5���N�M 0��������Z���]�ͩ=�58�P$쟈ȗyN-�'/��t���#��lxU7���2�k���O7��Cv�j�Ȟ�h�g˒.�;|V�~�ʮ�����+/f-���Z8b�Hz0��zg�$|��>H~�"L ��,�����G��.���=8Y�e,�p���s�?9�V�vރ]u`����>�!���٥�B|˶��EtH�Ps8у4x�T't�_�-PK�W)8��۾u�
��!��|z���	t����E��N����2ׂ�G=�z
�nrw��x}��vlg5cc\_Xh�#��>��ӱ��d^�j)��r H�^#Li��|ˢ���� ��F��V��	�����ͳ�P�\��Uޗ�ƙ�`�"� �h9b�_�Tu�|[����i/�ʝ��};�4wWw�tXŀ�PHfY�H��OM�P��ġf9Ǳ�*h�h3���܃o��\�᤟�w�&��I�PQ���kkA�OY+�Un������_U��a����}#�����$�z�IA�	]^�O�Ag����X� �Uř�\�d��xz�9�D��ƿ�����ʶ���I��e"c���(����Ӛ�H�h%"�D-�J���k�>PX�I����R�!�nj��C��u��  8׎�xr�.'���~"�	,����~iiO�W��2@c�iԶ������x��P��=��^ω1O�S���5���o_�ZC���މH֝�)�l�]��"���7J�}�i�yW݈f�
�s�������Pq����9�UݛïP2� ýF�-Ѳ:"�f8�:T5jޓ��W�_`}�b�m*��e�1�OC�� ��>�P]y���qy�.9�9�W�[@���\�U;Q�9Ȝ�Rb�EX��G�1u ��~�04N�Y��q�bZ��6>	*����DJ_��@��]�G�jy�K�"�����L -�?1:^��J�&��Eߛt
�	|q	r�81���D2����pY�-���d�C�ۤ@{g���<�z���~X�\�����R���}.Q�oڲ��c��G�O�I�V���;_b��۹W�xc�ot�������,�dz(��"�A��D��%|�ޱI�g:B�#e��O�Al-�@�X]T��V�$>��PX��㥒��@-�e����\-@�~��}���	{}����	���g|Bc�Upg�˦���;��O5�aF�����Wgv+�R�eq�j��!
����
,�=g>�96
>vp����y�,��a� �O$�����8�n�c��M݅��a��Y�y����w�WVܰ�=
k���뻭����B����._��+�8~�wT��n�rI��zO�)����
���/� x���yUp6>�@�n�Ur��M��&� �<�b�~��d�����O~�,T���[�f6M�W�%Ev���̟�vNt�䏥'���Fm��*�,�nt�^�T�쮟�"���c��:seP�4�=�S�IΞl�߰��&�0����H�]��^�K�U��OO��b��|˓�_�������֟�1��Z�q&^a� �]��$��EP3���X�G�;VfӜk�l����� ܖ�	�-��V�RT���?��x#��҆�{��MC��⦯�oH�S��0s$��E�a�qw��A�>m�0�j8�����w~������vQ�ZHh��;?'M]����]Z�"t!���b�<�i�(Ĺ�"��)@���t��E	�f�k�̨�FV1�}>�:�{{ ����Ջ0�]���\7�,K�\@d�[��%��t_��U�X��2!lE���尸�ތ�.�2�
Գ'�푴)OL���>�i���e�
�\�:�xLq`�'U
��S�^h�6�oN�]��:U��࿹ȧe�^���5����t�Xʌ&�qg�n8����x�z��-� �f���0�&~R9?i���3T�e�j��D���f��<�`V�C��Ә���Ẋ�*�g]�Vp�e�u�=��x�,&`'�P%:���,�ٿE.YLj 9'Σ�"X�r��=o�4$�'�G����8p�@	ɼ2Y��	iL���6�EQ��{�//����n�KP;�r+�"��C���ℐ�.�t7V�z��)R� Z�xj��5=v�=���U���x��;��-��T������ ��	�ѫ�X�:lf�\�A_��_�h��=��-G�T���j����7��!��Z����K�K���kŜk�T=��b���C�+�R]�U�i����Ռ#����\?Yb���n����#���K?��`ȕ��0�y�R���	��0�a����7�N�[~4����֧���҂*u[�T�jPY�b�"k*0�T��r��`
�3b���tF�p�~L~�$}��$����C��r�ˌJhA���|=�����Buw��$�;��
����&�Z�v��(���	�$c����&��e0�d�$ed���7���xQ�=j�@3P�j�K7<L�(�J*�h�5eė��<MǞ��N�SR�>���c���+�;�-��7�9��c]H�Q)��$bj���|�)�f��n���y���Ӳ�f�5��{R�ʲ˼�u����-E�=�`�-�+���MG�d�:TC�L�QB9�p��v90�۽��;���?3��:�Tװ2ǯ�t�Щ���_%� ��*)Þ�
�e�C\%�ك{b��V��E1I���Q�UE������d��*b���2֟2�JXVl&;���B�S���ߴW;T����}j[=�_�2��f臘�I�%WГj���;���ЎJ��U�V�I78�xF0\ߕ����.��s��O�Y^v\��J��"$��s�q�X�xԳ�#|z�xv(��	H�@_�<v�b#h��*�����p�����!�V�����\��K"�����f_tfl��r�3��&l��8ӶBB�_�ej��r���iUJQ7Cti�9L,�P��S<������v=�q������W#p;# K�&r�FM�#_���d|�x��^,+2���w⎮p�/���n�L0>ЄCs+�B*����APY�����t&\��D���Y{v���u@��[^�L`d}0�����ׯ�XTUpn�r'֪�x�ܦI�o���	��*��5Ěq�O�GM�����xȇ_��,�@ �ru�����Z@*�]���ZͯO_J����^����ia?#���z,]��X�<��T���T���A�������߁Ғ���D�W:xW:ߛ�W��%v�-|--���