��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jåا{�\�u�?߷�dn@6�zf��r������;�&��0����n�R���m0v���o��O���v�w��-�Zq���A��못ת�u#H���d'�D(��ru���@�#Մ��.��xN���(,��'MV*Ln;����-X�RNbL�0����V��h��}B������/����IKS'��t+�2���X��m�k�rl�Dv�E���l%IĠ_���$i��CX�$[H���ߗ�ͥ���sy�RȂ�A|֎�������tjU���eGp�� ���4.Q En�tD���Ŧ�t�""a5���sxɲ�ښ��q���!�Vj���9�WD�J�A!�=$���vMVƇ%~���7!ҷ_���f��Y���i��rDg7�U򃒡i��s���M9f{� �y�����D���SA��2����_'�r@�J��'i�K�I0/(/�Q�������;�tI8Z�V<b��>��!F�����3j�,����m!�+!��Q�=��ȈN��U��q�T�͇����������95�ø	�?�R��d��D��t
*��@�&�Tj����W
-	v����Q�nx��Fw�Li��>�,Mv2�2����� ���^����)���aw�1��y�X~EYr�ӆS�2�V�<m쓔0y=J�AQ���i�O4^Ԕ�'��x��F�ᤘ"�?���P��jV�R$�!�6N�il29�9ήf3/6ސ696�k�o�,8UQ������*���.�M�[Bx�[�_�����)��LLcd�y+U����bp��S�b�|�c*��k4w����e��_�w���*sV�C0�Ž�G�jƕ����=ԋx�ᙏ�b�O˙�"F�5w���*O�]r3&N�n�2d"E�<v(G�I�sG���X_`_=6�|n.��xS|�8b��%���S$��&\����25���%�`��@�Ɂ��B!����?�j3'�C�U���7���㖞��,�8�D�/ƚ��*�FKcd�S�Eۈ0��_�V(�Q�h����n�l����i��#�jDQH���ʲ��y�$i��P�����Fv�&o+��X�h�ݢ����ۛ���W8�l����K�������E�8�?��'D�V��9��^>¾��G�P_��m�6$-8��o&L��vfs{�OU
d̉>Z��8GrW�,�k͠k���a�4�x�b=�&'�QLY�n���~ʓ��s�����nq���GYi�b5�~��'�i3��Y>w$�#K�������LՀ�(�"�t�:
�/�vV�q�{���A� ��WV�O4��B��|��K��k�Y7
F�V�o�z}�Y��7:��>"_G�%���$�vt6��`�c�y�3˒���#\��g��h2��V{�宜�c��j5��sBt��)�^�ƚ�+�ߩV�t��(��0~;>5[g)��])nM���0��)�	�
;O\�8v�l2c���~��UQ҄�����+��b���%`�.#��F��"��_�<E+�D�P �����˩?~ۚ��s���y�p�a%ѲUp�~��v���%�5 z2J]]c0Xݓ���Ch�1�B�-��61E�R	�է�׸�U1Ѭ�ˇ!_	�Շ�.�U�*}��+�7˃�����yplj޼(�P'P7(:'q\?o�;��R�n��^}�����&�q���6X�SY�Ó��~b���Y�z?3�a�BBH5�:���m�C�9ʢ]g�W��R�l��lCo� �K�ji���1o0PoB��:=T�����8�~�o���U�i|��]1����0
(���E�H%��0�SfK�=Z!����D�A����8��kC<6A:��M��U�nU"$I�lu���&��J=Rf�''�i٠�|��;*��.��I͹�<�<"sPy�~Eta�c�y���uc]a����N�����AJ�P�X�;Z�������TsF/V_���C�J3#�U݄�Y��ɦ# ���^���k��K���ԇ��'�j�Ѕ��8Xoj���E??�������]�G�p�˧o��jC��L}}��\(��La� ���n�4�O�]����GF�BA��
�Ґ�:�%�ƨq��sv�Iڞ�>T��u�y�ț��5zBN��#a�������nt�冶�ć�}P��� M�%����~p��@8�EB�?Ry!	��:�=wnΙ���U��蠰����B{��Q�Z���D6v¤�ݺ�v����^h_l����Fk��S�P��B4�&�i�a�@q��`�=���e��}��e���h27�t��Y�8�o����V8�#;�D�x"�:Mj�E�k ̠�N�ۨ{E��:jTZ��z��cϺ�����8߿W��u�.3�#�TZI�G� ]���E��2Z��8*��{*��0��뀽e��eONٱ���f4^�@�A��Z���g�r����muyp���[>������]{JV���f�4������{�U-���V8O)�j�P�@����cR����
^$�Ԓ	�;.tt���k"97�>�CUn�u�e X�.����ݢͅ�������ں��E75V������?wN`Y�;�I[��%�t_(�?�5���s��C
pdAO �fhӹ�L���4*&�+�uߪ���7j���z�����Y�R��d��z=�����^�z�1s�d��࿯��2Q�5�:��c�	�M{AȻNS唗$���`�b[�[F�`u0=�p0��A}��é!|��(��0��)�?���]�{5����֐�U��%�Խҩ	�*�Y��>a@z�D,5��|��Db�D���h]�8��u&�FC��h0�OÁ�DW�'�5��'6�rW'�2;"����P�r���K�Un
=&�8�@�lmB"o�Kƴ�x�b�ݺ��&��ʾ\Ϧ�%F*v")Ց/���3�S�eV�_��SN�ȴMwUX��<�����+Nƫ��3�U�-�U�ӽ]>yv`��a�qJOz���t�ѣ-0@�^Z�{�C��S讓�N�F 8@ۺ�;�w��˔����3g�1�ԑ-�n4M��`��I
�T���r�lD8L�\�}���9�K��!HX�阈����X����Y��jPt����WϊvoP�-�b���oB���i��$3�=�ש�X����{d贽�b˶��w����!ɯuگXe1`�e���莹S�%1ʊ�'��گ,(53S[�24�Ԣ�~V<��� ���#_�T�m�E2V��h��D�=��h��褚LFR�O��(j6�QIfɲ����������%"	4�rA"]q���x	W�@���ɼ����tJbN���NSH�ϲ�&69t7=���	��Uc+C.Q�hi�L��@E��E#=q%zI[Kl8`s&;x�mU��������������᰸8%tpDԻ.��Ǔ���\v?����L�6
���"�Ѧ�tl����'b|ۃI�?Y��db���`j��'Ir  d�,N�	W�c�0�qm^�=ϢZ�VGo��fݬ�>�ƾ�7�9�ꑅ�j@�7r5�o�i��Y�,�-硹|OT�!ib���{�c^4��U{Fؓ��򓛉�}B_4��#N̖�-ٖU����FY�_hpvP�h�:$���+<2�[�؊���c^X�E}�B�s��sx	u߯�<����e�rBt~#R����`����{#ŕ���`��������UѢ�.��orL�1����}/[���ƴ�_�[�v�T\���a?LD�($l�$;������P�{:sF��rdQT^׈��(�����^I�Y�n�?"�z�Oq���>}ȄA$���/x�����;6�������o�1��S|��$��N�mL|����pd��Lz�F�"�`�e}d��B�6m�R��(����:� ��]5�������I6A����c�e�ټ�u�h�R[��|-��M���'/!�dߪ��3ŷM�Mo���\�3��?<v�b�$�."�C���޲��p}���.����BGO��R�g�.��-~����iD�̅�!�Y���*�Սlm�ףxp�w�#P�����T������L�[Ld/Kֻm~�^���
�������w��H���
��;�w����\ȳ0z<��t�e����6��0� �)��7�F�0��A�?�5�l\�d�:��sj������|�9~m3{M<	���Ji���\�Z��(�����k�޿2��z�[�M�l.p�?�4�g�<�� �+r��#^rQ�Pc��v0�J+=Vu>��(^b*�(H�^}2��TA7���/ :	��5^J"4#y����9���I��1{[�a��i� �	'�w�+g�����d�h�z�_=H��Md�z�o�8��w����9��-`��q���"�_@h�OT�B�����ϫ`U����,N��Ͱ(����?L��J�C(��C'C���Wa����2�_�
���<�|��< C+�uj�d�rF"���w�+�!���F��t�����=tjK�,3s~a�����*�ƪ��Rq掬qV�?�Җכ�#6T���6�̌��Z'����t9x&1�N�U4��P,s0��]��w���}Oy��O�f�5�����%;�T�aE���b)b���'}�����kl�����aU�~�8�ʐ�Ύ���7)�� �g���%�y�R�%��	�T1�~ڊ^��O�Z*���\��������GZ쒮U��гȱ/6��(�N���Ƚ᛿�� �q_��<�!����e%��)r��`b��e����\�Yk�� �jp~��L����ywn���y�y��j=�{<�f�hPD�B�{<U�!��^��5���~X�'��������Ė������J�����np=��S�R������e���0>��m��[�	F�l�	��n��,k�ߊs�e�X4)��!� �:(`�H��-�ɘ$B]���k&Gj��LEAh���V�����g��Ӡ�,+��ԫ�"���1�.���F �j � �j��ч��Oe�!���@)�T��6ɒ0��V��}ș�FM-s���xd�ߦ�ԍX`nJ�+�.�v�
B�g8e�h�kہa�TK�aͺ	2��%]�܃�|��X+8���-�̖ܣ���^5ס�*�9K%~Aa��	 Z&
ݒ�0�����1���� ��Me��1K���<����r�=��?�}�O��l.=`D�SRȀB�2U�}�S�	
L��I�ޔ8#FZ���FvxF#�Җ�YԭϬV�_�_0���-H�$�k�d���PX�v�=���������g*�u�;�����o~�;zA(j��Þ衡�����/I�����-X�t�yX��ʥ	/�{�_�>?h:�ҷ"&dI��e U)��-��*3��.��;�q���;�8"��&@K�@d`pq7�01�W��F����Q{$]��w��G7����L7\��f�_���Z��	
Ok�Kj1���(�V�&Ť��b�B��GX���H+�4�E����`g�Ζ��3��������!x/L��)!|��x�{��*�E�L�iZ��2���S�1���?d��]�������)c@��ˮ+>� ��"����b1u��'=��J#3�lA>�CB�iFDR���I��`�w�Bb�y��[ q3�[��@���$�㙾�'�E�8���Uv ��H1Ԍ^�(��ڗ+N���q��urߟ�-0G+W��5��F��f������IPC�i U�N��'���!�?��r�l.L?�p����3�&��S���\�w�UK91���H�-N42yi�k5dO���#E�<���z[��������;�Ǿ��].Ujx+y>B�i�M/v۽ފ����z#{�(&`�G��=G�W�p�nXmX�V=�4pU�ɟ���2Ջ����2e��I|�s�Ne�;�6h���nڡ����g�x����1yz�'#;��s�7;{��
��-��J���c9N.3ITf"����rR��@�_��J����g�o��,:�O�<��YVƆ�*G+�o�'!���|`��;t{	D@����̧)"��L�#Ŝo4ƢO�nS c�|

*�P�� �o���{���T�^/w���86]�����'���[w�?&�5Bn��j��>��?��M�9U��@��ʹ|P���FH+�@�>�hg�����7��:�a"�w��p�& |v�'���1b\!=[G�_Ւ�����0}�o)Ϛ33�t��6}m>�1���z�Fl�#�[���c&�`��Vƣ��l-\m��z��iCM�ୣ��v��A���������77�飻�o_���V͸J�R�ܽ�ʀ��A^1q�#�.��e�ha27l���������o�9tpE��7-��0d��?S#X�
�/�>%���Ұ�I?�93�]^\�HS)�+��]�;��4U��fCy�w%�x���Y�	�d�u?�6vc��Y��g�B'���ZC��)�y�4���3$rfE��]��fw
Ӟ�� ��?r��&�1�n�V;f$�9��w�J�|&�&96�Q�,r�O'!|,�h��� �mZ�hdOZ?|����0��	0x>��>:�X�j����CͱN����n�{����}������%\�E��#����i$���>�n�	�`�J�^Q	�َi�R��َìmVp��A�ˠ<Eq7�o� �+]O�s ��;�j�S��[�vf��<�,3�i�~G� ��<��1���P�k�	���L�^7dD�C��Uj�Z��O��E��:�f��a	�P�f�O�La�H�~���6#h�替�P�P������b0]eG@��>w\w��$YZ)�Z����9��\���rJ����|������/�OK9�5b|
���%�
�u��V��U�g��ȍ���#���`�c��`�6$<�z�,�fkD�
�,P�S�
!�q}~�l��{�T��]���e��-a�o	O����a�>S���&�4`� H�7���y�M+����~�.;��:��R�cw����	M��7��K� tS�Y���x���&���)���x�4���@��4�M5xZ�/�U�'���5J���>v�ؔ�æ��A�P�|R>?y�Q3L}�L�B�í�޲A?��3$&:��{?F霩MJ�����D9s��T���+�^�O�M�H;�yc���z�!��R5��3-~WB��h�k���F�U�����Y?�%*H���3���w�� ��F}���)zE��vtg��#���n���D��e�rt4���؉��z[ԝ�����R�t1O���ȟ�C�}KTc�L�|J� <�	��r�-7h�E�)����e�)l�b)x1(h��
����l�g�L7Eԃ?�W�&�����N�g�i3V�+���L�,uD�BE��B$GzU񥗸�8���\�# �ߛ	�-`�cA�Cm��[i���/�o#��7My���E1�p:R:.6i̐��Vr���)s�x�5v���-��;�S	h�#�m��"����mv�u��\�3��2Cr�m�y�4f���̦�}5F�83~����9Il*�ߺb�M���񍤡^?�-��ۜ��XS�$Ƌ�5I?��{ozF ���j��ř��ēe��.`����vg']5B�� %��gx���->&��; ��OS�%�>R�� ��|�;v�"!�4?�kR9'I�ݖjyO:��� ���p�9`] Fe$�=���ק����Pę��Cnc�~D;���,V��7�}�%�ߓ4q���Z;�L_m[�q�M�hL�XzVS�����֝J-0Bw�YtH+C0��#L�������KH(:�>SI��Y��������^�D������F��v�`$�~��q�M%Un�I#��`�R�1�f[r�������u���6ʔ&�'�����ǎ 	,P\�Pq�cJ���HLD��'��7�~d�/l�WV}S����b�v�3ո�?Fr��[u�����$�Y��^�3�i�z6˶we5�/��;��r�r�>)@�Uh7��T�Av�f��,4p��l��o�%�Ư�����Jt���

f==3�Ʃ�Y��VLbU+�B��,v��C���x##�~���D��x��m���j����n�dj>��_F&4�43����d�OU��f����;:1+~��#i�܆�����l�d	��ƛ������vk�`�HK79*!/�CZ5xץw�EJF	���#'5���:_���X��;��:�o% [� ��{%Dl����]�[�T�7[F+��`q�M�X�&�����50�@���q���OY TPf>Ph����o�-
a*��1Q���]�-zYi�����l�t�W�=�n�ҍa���Н&��I-�T���ho�$�����HD��ܜcSړF���;oZ�T�~�b��Bm4��u���%�y�����<R�]0:��py>[m�B��y����\�� D�K�zj���d~8�������J9WsP�}�E���
���BW�P�Bf��b Q:V����ku��*w���ث]���V��J���mQj�I1sfs�ӑ�L"i+jGM|��"��k��R��^��^�&��B��C$mJ��Fo֚%a�1�C��( 4m����6A�@}5/7�!c�x���5��Q+���M�69��j �7��)UV��m_��LF�ڮQC'/�5ն�sVQ�;_�V�nς<M;�Nf�ѿZ�1�U�n��yb�8�tis�'FJ�W>xT��뮌37�'Z&�:�R������*�!�~������{ ?���7�D|�1�*B$T�=�V�3�n�^h*� -�0|Κ�s.@xԚvfJs���|�=��B]%% y�v���Ng^���>�%O���%p���=�ܒ��!�����q�2������
�2��ϱ��-S��xY7�J8��lT[�kk+b^�������n�!`��>��'Q_|���v:2�~���۩�N�>�`�M��&�|x�K�xt�SNn\n��U��)_�����ݯP��x3~E��"J�Y:�Qi��wX�)�:L��s�5�d�o\\��7��#i�vR#���u��Rv���<��*�!]@�s�<y�u��J��Ou�Z�d���F�A�o=�x��QE��.���0 ��0M_л;���Ql��un ��[��z�,I肆6�����i��;d����u��G�����VÝ:C��U>׊�+.J2~����y����1��\yE�h���v��W���/��{o����k��[���cݑ���p.Ra��#�%��p�ᴦP�
���f�� d`����Q��u�Bɩ�kx�&�m؆��S�s��4íP Oo8��*�ئ ̏��yv�#�DAU�!Y�@����Yٶ�AQ荵[��W*�ϑ�7��h���*'�B����S�'��ˣ�ׁI��|��>�F���6��5���y��gg�2�Q�|�����;u֩��>��q�Vp���dO
A����Ƕ<V>��h?�?�6��Qd\*=#ݤ�tG80�9���K���#|zZ�׬b{^0[�u���G�ٛ�� �;h�',Hb<((�5,����&�IC�H\�e�&L���9Va��G��w3U��=��X�[�2��d{�DV�Q�y�
���CՈ궎}��*��&X:G)<t����ŷf�I]���Ua�cO� �[�o���0?�d�Ĉ�'�/�CLNw��u3dl�������
V䠝Z��"���U��Q�j�x�⏬�Jd
�`�v1�NS��;�J����|6�|��XѭO�"ʟ��ّ�e�0�,ؘ�&�Wݜ6,c�c�4[l��" K��G��!�%�����j ��l=HxbH�~.Ȍ���Ş���tK��*"��Y�ƅm��&T���Ȟ���tR
"����ac�a`�boU�s��_F �!3��b����_Y��5��*�|���;�-"Q��vCJft��xb�t�w����G��u~�X]�sy~�K
���x��3�˙,�*@3~FLqa��\
p@�4Ո���~��#9j%�&^�ݛ���K*m,��2�2#���T�V�3�� :�'>�|�A�\.hf0G)�'���&�+�CF�νߙ�o�}�`���D�3%?����g�t�$6^�K�.U��#��?��oq'�R�Uh@�hx<���R�a��q�<��@)j��"�K\Ͳ��w���S��U����	2H��2��RQ[��USʪ�x��!¶	���i��$�]N������ǧx*�P��Y̗��9j'�RL̡S?4�B��V��cg�6�ܬ��5��*3�i�h��w��2g8�]XU�U�9�OW$<��$w���ה�o��&�ofm�-. �Q��A��;�M��D�����6/�(#	0ܕ;��U���+�At�d4 �R9t�D�i����`&��6�r|C
ؐEs�h�ؚC$�E��Q����n��3IٕDv��F���y#��I)����+3�Z�e1JZ��*th���v�4�S�+�k*���̴��������A9���gL�;)Z��=�7�Ẏ?u��H��N$�����u��_���2�J�o���[wȫ.ʘӰm��<�P���E89l=9h���U/cs�Z(jA-�������Q	xR<�7��2��4Q�9!�J�>A[�����H�I��<�Ӿ�`�����Ty���R^��|����O�h�ܡ�V�A�c�e͚\I����FK*ߴE���YP=���M�HE_u�Ѩ ����%myb�V��k�ۍ��fl�����f��Uji�ǒ~{:��N<
�;�|�Q�<�>o��BL^�r���F��w����ɴ�u��9��3
�R�"*8�SQ��x�0gd�W}	����k�Z�w9�6g���Us!'�����GL��G˄��1/C1�pl �M9�Zr�wf���g�Ly"�M	J��Vs�C\S?ˣ�ݬ���`Q����}1�6����'ȳ�P��?K������Rz�5N8���:
:V�2T'�;�[������5����ب�ċ`�Ϳ=�C1#� c�����]c��CW�x�/�(�>����X[G��
����j� kE4
���-^���A�IL���M�Gt~�dT�a�O� R�o9�ƺL����сa^�k�Lj�;{����r�"���r��։�lC�ԸX�T�O�)� 辢�Lq����%��fS�?�b�8-��P���ޑ���<~X��&������T�Ħ������~�˥�ŎY��%����������;�ʶ�9���Y�u{��#��'�V�0]bn�������� h�t��(�Zq�d�Ƴv��\J���p�>�w�
yf��(��
���&��$�`��*�J�'���(����w-_��gc��1���WѢ�L1)@vP�M���Ử]�m`۲T�����;.��>@��*{�:���y�IQ�p��	f��F�i��Ype�Y�%�r����Qؤ(g����r�&��p�V4���8�a�+$�)랮��Rs���SEoN����l��$����kmaR(l�]�!���� �t#N�`.�-���F�/x��P[��?U���E
t.�]s���af�	�՚�������O����s�C%v`2��'��M���^g�u�Q�A���Ph8K	"OD�>��F���w�U�̮/
���l�`[(�t�"�yX�(��m�e�[�I��{/idøA +���1eL��$����������ϋ)��7^,�*��<
D~	���Xe<_�z2�S�aɵ"��l���ߥ�n���GOtG��t�%ɐ��7׃Kd�����\��T�a�*������
���Ǵ�"
P�b\w���3���BE�e!t�(���o ��p� �r���������m@Msg���g��vP}ǒ� *�W��wS<�d��BV-  2Hi�=(=mcN��y��\FŤ�9���]����'M���\j9��H����G��2J�nUzj�&�S)���_��sgeN;�%��3�����5[�R��oP�L��H,�����,����o8}�LPŅ��}�X0�Pivx.��0p�p�38睮�S�zâ}�a�&v����1��5[~.J�:	���@vX����X�%g\I�Wvr4m�%m��=%$.By딴��v��f���G6��/}��HE��e0G�ZE,w��P�K���4ݲS���5��ߖ���N\�����LG��X"�L�|1�������o݁��(Jg����k�.M�6.���]ps} ��H�s����o[�}�s�G"^�F[z�X�Bg
��r�Ge���2/�+G_���1��^IrC@����)�G�W?iI��#�$LA�U�+R����~�=
�VK�^�8�M�,M��[>GA��A�4��\I��ވp٤�����)�|n��y	��/�Ww�������)��Χ,����:�ܩ����l��!����-}Q������/W�t�7C����(���"3ǅy��w���@�,!i�_���,��x���9$�>>�7�%��f;.���&��J�)56�>��J�����R��k�P�.�� �z_�!?.�̏]�Rj��W|�XyX*SKazA��ƀ�d0�ԀB>NCq�̤�lxė��k�8���,����ф3�C=CFF���l%o�yuF�F�~P�>>j�љ��_`�|�ۯ|��.��{u�D@Me������x�fYw�!N਒8��h-+�[Ћ ���D( �uǕ���ϠD��TQ!����у�Y��M���$b�-19@�~x`�gb �y u��r����5�
+��ɺ�]<�q����l��,%��4ܥe�N���o�l(�54Jl?����� ���=S�qP�L!I�4a�nNc§�E��/���CxmK@�os�S2�A5�>�G.Β(A&f��@��"as��G���!��L,N�d�k7+~YQ�bP�}C�|��UG�3��V���kc���jN���z��fn���<��r0���������|ء"֦��v��39N�c1����X(i��Sإ�H+�b4p3k���.��*�i���-��n%�9`«�w���I3�_x	�)^��(�����"O&e�g^%6�X��@Kl̥ h��m+���{���
��X�.h���O�ab��]i����8r�L��W�����J;��¦��_u*����Ŵ"�sTR	]6Ref��h�ޣX�L��e�Ί�b�%��H��>9��?q���x%s{yG�`���Q�0���G�h�Bic@]BbJ�>R���%�($�\#20�Jm��̅��bϩ(|���{m8�,�j�Z��n��񌏧�$��;V��O��@9Ǭ�j��DH,���)"rJq*�k�6>M�uv=�324�Nj��KH3*�� �U����n�"�t�D���:^v�#d���a~$T������S�9�|ir�������Ԋ�\��<�l�ā(L?���	�-+��Ij�h��L��i�?�"릶�F@�k�S>�x�"Z��5܀����V��I�ِ1~��?2D���۬m���Kk����cX��('�'�;�X�*��i6�e
���)68��-[�4��}+d�� �
5����X� Yz^#�>��qT�1�ڜޜ��yT#�ˣfJ����
� �7��'sN�X�W�ˣA�n������H�0>�0���y
zt#LJ������3�	�;��=��?B��-T��}8J�|n6�)O�XpOL�)��U5r�f��|P��B]m�k	Y����y�It�az*JH��ٱ��C��Leq��_���۱�qC�=���s�5G�G��a�iU�����ʅ�:�����r���-�qn�Ek�C�LI7n�B�7���59�.���椨��E�M�T��0�U��h�D���b�Dr��@gƊD�`�A�`+!a�*Ǜ�P�܃\i�mމ6	�PLwl��b�*f�X�Y�qG���g�I|�\�q#��6����5�����c�ht�ښn3)�������Ж��Cy:{���vj����0��|�Y��8<�.Brٸ�D��iԠ�Ӂ7a
ϵXi��W�`$2zm���[W~�&8pl�������j(4���[����O�[�EBP"���z4���Ԫ�~��D��WYh�TN�ʥ�J��t/�a���+m��}�1���z��<�@2�Nu.N�4�}1��e!F�:!�N��k�=l��/�h%V�h��㗅"�1�Z�O�ek<.�iγ�y}�+q�kL�"��0���x"��T�����$��빆I3sI�+�Pq�K��_��Z羈�x-�
A{h�\�m�iPT���ٲ�wd�����?ZOf8�d���:�?���
�E� S��wfmx�g]�q��g�h`Cj��$7G|2a��7�\�/�!y�c��<����q6 �A�Ѳk���|��$�ˋL}��YrT�ޢ>B;#[UL��R������Hk��V>^�½&T`�_�jD���� �2�7��u���Z���.�@"um��#��$��k��aW%���.�����+��r�pM-��o����n�q�\��Z���(���}˽4z���i3��������B��m�7�6�+�n�����Ά�vO:z�1����pX�{�;a/��-�`�S>���H�u_��$��$L�x�a�X����1�͆��nt����>��Ҿ
������G��,�34r;a^
�|�6�/+���f	�%"C��zz+ș��mg�g��9(֏.�tnV�:E�*�~E������G���x�e_[��g��%"J��UB�̝���3���z�aB�e1G��B6�-^��K��Ex}��V�S���ΏSO�n��v��E�	�m5�٣5b$x�2՚%�D�ݼ��f��s�����-����:���F��2
��
�_��?|�UG���@��mE�5�:u�/]B���R�4TD]!�;������#6�G<i.k�C�͔=d&ٟ}��~ay�%��c�!��ce�n]AU,���B�%|E��-nc�q�$�EK	ӏdb�m�vlt�7���XqZ�izuq�F��!*u�[���S�)�<{�`��ѹ��5*�e�	���ߦ�Kw�����켖с����<K�01(����K��Dq�`[� �/=�0��<V��
!����[΃NOo�[�#�H�k���λ|�����N�J.�2�P���ͷ�ы��v��T�W��m\\�k��|gN#sj��j����wE��'�e{5sb���8�#<�y� �!0_6�M�����1� x�N��Tm�v#']��Z�B���Nc�oO>NgzF�:XʢًK-�zn0�D��Y��Hd�`����NYJ��o�p(�L-�Z��)3�ñ���I�E@u�	�>���W�f�r����G��w2��N�%O�3��5wh�+�kg1k]����Px�&�Fe1dI�鼛��Ϧ^�Ze4���ǣ��G��U_�U�"���\��K�/����Ԍ92�\|��:�KOG7/q�y�����h���P�F�R�5�p��2+��5�׳�9�Sx3�W�r�Y�Z�N͠� �Sc߇7m1^����i�������͕���U���o��vE�]�Y�?��C�D�=�����Yum�*M�t�=k%�i��n�zU�p?�����`���F�|!Ӳ+�4�ߺn�?
��,��m'��Hw_x��r��,�^��ǂ�)3<)N��,�qb����1tQ���-�A|���:��7��l�
����V^��[�����6� �}�}�yT��Rۡ'm��LBpJW�����^���u�<�]S��P���d%;n<�D����C*���b_�!b%5yZ�"S��~O���g#���MV)8/Z�w�����5S���9w��F�Zܔ�������nep��F�s W�o��b̃uؗt��j��ᦶ �%W�oĠ7�|����2����6I��Ȝ � 55�q�ݠ��oP>s�M�1��-�RD�-.�;���,�.^��gэ؂�ӿ�E�"�Ѱ�r����e��	ԇ�L�.�2C<X�:�I�1Xޟ�k�hx��أP���ۃ~�ý�*;,��0R��	��
j_����%�bAE�R�!���&����.*��Y�|�7�2`Yh�J;˒=J���uGb��X���^H\=؟�|'
'��iL��1�%ʠ���X����{[.T#ϛ�ǳ?:Qo����0#��a\2��Mէ1��݄�E�4:�# ��Q�z�"v�~��MqG4�7��m���� ��ԨN��Q|M�'��m�t�� M�}�o]�}:�J���I]6�q�EӞ���(#9�(�V,���h1cs���/o�Ǜf��ܠ�h�x�߯�f�Я)���f;n��#֫5��7����8��%��M�?�ÎG�ĥ�,��#tLn+�p�=�.T�9����)s����G���EN�
�M`�V����d~j��Oj��L��I�+�(��o7z�;.�
�! zYwW$+�ɢ#D�ĥ!�e�p3��d[gn����?lI2�4<|��ͪQR�&��)���;��o!,��J��-���F9�l�T�E��sr�MeTݹ��c�*� �?��O<{��M�6�����s�[G����h8~)�T��sE�
�Ͳ���[7#��{,�����`p(�S���	n���
�H���u7@M������P�YfG�d�_�����l���^���'�t��j��f��U�bFPbJ�dH��WXCht������};�g�����j0�T�s �>�9�����G���Xsl�Y��1�V�͋{{4ۻ�(*'���;kB̚�B������!��c#cj�����}�� ������=���Y�W�y���$L�%%j��T��ص�W����^�F��]q�I��6B���.���}8�ש�*��B`N�Kf��2�*)�kK,W����ry)��<cPe���7ߐl��Z�Tm�S\ }եn3�lq���J�)�frG�D*���^#�3�9vM��A� U���Isݭ��HR�����K3�j��ϥ���ʌN2k��lR��#6>�Z��{�����UZ����Eis�_�.�Υg�HQW7x���hK��@�G�%���Ev��v��,��un��/ka�#��8�B����H�f��u��ԓ��k�����I��p����7�|�WQ�������x�P{A&�����W����|K����s�8r���Y��!��~d��#l�x��#G �?ȧZ�"5Ĕ�?�{��0����0�l��H����RA5��O<��^��o����P��%�=h]���6z���ݔ��3��\�����#F���p0���yX%ytQ�;����e�K'��p���9v���-��u��5_C�&����� YLU���@ۅ�!� �K0�B�?K���o��%��f���z�*p����^���jB5�5�֏��e�-#F�K���;g��aGnd-5�`@Q��JL�B�B�s7r�	�b�/H�Ԫw��Q4�}Nin��8���c+��44��A�������G��h�x�	t�}�[6��<TL���H�
QP��w�5���)���+Ea3����RY�{��d��&�1�P� �Ȏ�1��o*M�Z�(��J����8ok�H����(��4)�1�n0��'�$L:[,���'��~�?�I�|�:
+d_�mp$L���J?�w`�lM*��ڗGDY3=�\'&t}�Lgl㌻uAO�CGyW޾%���~��pM�r��iɍ���+4�e_q{����Z�[U�ۻ�C߰�,�EZ�=����Q��)���a2^2���\:��f���FSmba�,�W�����aJt��q2;���R�=�o��[�������`�5��X�ߺB�����+��t�X��v�,����a�ItW%��f��� <�vb�{�A�mhE�T`af���%w�I'�)�Ca���I|9/`����M��y� _��������'w͏�K�[��8��y[�A�Vrw<[��P�!�*-��:�Ns(��r�N3�1�Sh��� ?���uma�Qq��rԾ�W+�lԷ8J�Nl�C��\�}Vg��N��^=1��}�Fi�
����
?<S���Y��.\4vu���{�s��*�座�j�u��?�Ƌ��ze��$e�}?�`��WeC��1�K�ߌ��6䶝|��&)�9Hō�5�m�u��.e{),F�)o!b6��ܫ����?������}��_��=��	&r�X���3��Ź�pP�[�ơW���Y/<{�7�UYK�Hw�+����k �u��X�/��ίI���l
�C(����m܅̤����bI_x �U���^�NPS5dNp�V�	��ݦk�VN��l^-�hJ;m�:ǘ3�W4CѦ�y��5;a���94���G�0-�KQ���}b�ZL
D�VE�$����w��Q�l.��s��4�O9Rvu�O]:�g[qԙ�F������-���T�=R;L��-�R�ՠh���\$s7��;�������|�op7P�5�ܥ+�d5ր���+-��-���mw���^rF���e���OgD#�W�)ԱbP�r�3�T��}��k����WTF%Y�W��� ֏���|����Ry#�G�e��.Z\}�r�Vʹ�[x��j�A�g�����SS���\��Ix�u�i�|��A��c,��n�r���r�*^�>zwk(#e~H���ʹwT���} ��*֕f<���&%Ǭ�IpO�$esPĵKv]�l�¢;��te��ĲU���Q�8�Z�¯������f��&����BTm����o�t�d"@��	���L���˺��ga(b�4S��b�D��0УU�D�K�FGC���k:ӛ	����0S*=4�_� q��@�8�N�~q��8Q�	���M0��ke
��QG�0�^O�I��&��v�/�}���5q�ڸ��Iƕ׸�7� K���Kw8'�h>9�2�^#�1ˎ��76/���j=�J�.�{��ņ�n��ee�ɯ�1��r[��<����"kf�����"R��H:ˋG�*>��I�s`�����iFɔL��T7��{��e�Ⱦ����	���ң�h�WhY�p,����<Jf�C���A��� �)E9�o�x/��fC�R��� ]��iś�H8Bp�oA��B�f [��\J�p@�J@xi|��,�d���j���LKz���=�Dק2���vo�	��q��.�ŏ�_p�LH���K��ɳ�:i!�Y�R_'��y�p��'X��T�L(=��+Ȣ
���Uʸjg�R���gW����Q~߼���jy�8�)��HY�6E���U�?�{兿�xG0�H�'���5�% w��a,��MN��-��J����G.�8&���	� S(������׳�i���\�?��n���^[��Xc�j��I��k���f6�'Fq�m,�Fω8��)e2TUp�p*�$��ʿ��+��X�oɟ�\�����8�*�űA]��$��K���j��y�$T*
,�xz@��'�vCe3�t�JG��@���(�eע��<���#��U״(��� 5`�2�jg4J?�a�����Y��\L*sn�ٶ�6
K�����-�ʴ"�B�_�R���:����t�F<�
+�WY�>B$!�ϓ�̃���{R�dY˒�inC 1�$��*~?��_�*��%����C��E���0���]�)��3�յj���2&�A��-�J>j��=K�5��~�-�O�:����<]9�J%c��*��f�Jxiwƶ��e���	�EH���rms�+�tx�FR�ʙ2s[gpe�Lb�T��G�mh�1/� XP��[��т0PD�����P�MT6z��ǻb>x�6�>�?WB�c�qN��җ�L�Tǩ�ӯ<Vh��9��u�wj�	n"|Q�9h��c�G��_��T�ʶ�g�])�h�rM�cv�-���3H0XꡅD77�6����4�R#����t4y�Y=��u��&��ú������@E��[!:1�+r�/�^�҆�D.&��F�)wG��C�k?���� a`�Կ�ibsX�#_Z�m�*����oAQKO�O~|=F��&��7�tM"׬qP�sR|3z�
��CAl�=����!��2�e�������l���׽�惙��ƀ��2��`�G�4}��ph$;�Wy����Xn|�����vn��*�}#�X0<yZ j�c�W���?�ET5�!j�2/�ѷnM�Z��w�4cuQ��>��\&�+{�[��"����o}I����%3#��Z���4������K��ʐ����sE-`�4�������9;�7e�˛]<�u�e&|��^��0�Y�P��u������Q� i����)�T�)Q�G��[o���b��P��l��~���4��7��&�O��VR�/�W*�6�t���F�:C�QZd� q�hljGe-�R0߅��$�oiR�Ƈ� �������D����V@���f�ɟő)0g��t	{����l.t8 p��j_Y�����X7d�����2��	o���I4��Y��7��Rld8j��	4�A���C��}���tXR�j�w�.?[�Wg���ޘ��;��h��)��9d20���jo�B4�2Ӌ�d@�d![��8z��r�4p���SJ��{慱�-��w��r�/��qv����8�E�X�uR��7���N'#�
�xr��Q��,4�<�%/<o��	�P<w#y�.�K�`v����p���k��3��t���ź��v�������������9�u]��x4J�5�3��"d�5�"�]��Fi��)~5X�>v�t��
U6��G�zݬ/0�P��r��	��%� ����Rp��Q�qn�ap z��S+�9\�#)�j��|f����$�+��#R����c�8�30�P{D�j!Ѿ�p�w)���F,��-����Q�o��iƝ�r���
�:����B�L�:���{� �����lד{ZyK��=hP�y��3+�4.z4RW7�� �K����Y������5f�'/��@|�ͫז����j�@w�6���A7K����0ٰ5C+��r3��&�_�&N�P���Q�����3>XkI��>��:w��[����%Rg0Fc��ɊD�
�Y��E)a�Q����'�y��m���ȳF3&B��#��9O��)ȵ�'͑�>��~���2i.[� y�g�Y,mƁԯ�{"�b�ɟ�� �;�z,7��ߛk�G�l�Ӗ>�M o�d�ZB��[��X���}6}��	R?�����
[~��б:[��^��+�S�x*)��v$f�^{8A��j�RF�z&}��A� �[�dP��8��{��c�s��5+q�5�a�����daKvl�0���A�7�C:/���,{ݭ��Җ���V���!������?��K�1t����[-~F�x�1��x��Y�?g� �����V@�$��bۊp �@@ �������V���E��\���U�-nu�l����aرa� a'�u
��|�KE��=A��<]�7�Ȣ�;Q�S�ϋ�)��Tn�D��Ϡ�� hU=71��W!���"|���4Ff�] ���#G�Ю�W�+�Ɂ�]�I-�'���%A�Q�C�:ʶ�wYܓ�Q�l}�/٩P^*��ro{^�N�{3��?�0N�%�L���b<(�w��=��X�پ�&���8~vG��u�B���R���1g�q��+�J����+)	ݼ�>��Ϲx�0����^�X;G�e=ڴ�F���;Ɩ���Foq���YTS��%	�?��z)�抉͌�du�G/%�vp%#�L".�zyl�)��g(z�ι�����+`�-�,T������h�q7p!Y����ž�މvY�����i;��k0��U0K���z���E+Et.��"���8
!i��[���_)|����>���)�O�045��������Tq�� �Q�9�Gj���B��=Z�gܫ�N�SI\9a =�M����Pl�n7��u�t��a�q�&Ƴ���gE��'~{N������XT��Z�#(���9
 Ғ
�G����j��Y ��|����ޜ�˷�-Jt��D�MǢ��Bұ�m�,h�Ú��L���e��w�$��.�oU�\o�<��C&�2�ԙ�M���O=F�AN`{��;�%l�pA���e#;$jVM�݊�&�i��&N8X�'@�
W�2|WU�d�v���&i�l.�4�W������@�K�yL��IU�zQ��J��ܟZ�JfL�-��
�Պv�䮫�����+���.	���K)���댝��g6�,o�����O�q	�D-��\�t��J�f}�V�4Oi�3�;���)o�~瓰�U�\Ni|��bq�k��R�h5ǔ�	��n����r�En�[_�[���>���-K!zu�����j�"!���Xp��!W��ߥj�f­��r�<�`�~w���8�K�P�~S(M��Yž�@���5G��B�t�XŚ���~�Ԍ�q�DQs�]i)�\#�Ogn�~��6��ْ�X�Z�����@����p'�����0H�Q;��f8�E��z���m�LC�M�jџ�?��h¼<���H���aH���d�1�PDKAJh9�{G%�x�S�8��,�ޔ�,���y��h����~R�
b��Q��Z��o$�`��_.� Ӓ0����[&�z���V�,NX����?�8�[���'�E*��yX���
&ol_�)r#�"�$[dn��_�|dv�[Q�HL��,Wx�lbY\P��-R���}�_O���6kMPs��GLu7���.��$����JZ�N���?�=�yw�,6�n��u��>�>6jɅ�w���=��l�"S<��:��F�	����(�է���1���G�X�`*>�]���=��9��~�	�?��\���2b�A[kG掭Ԡ�񍚬��#�rʖ�����TzY�L�+�eEh�_h&�5)v���	��&�-�豦�������[Y-�^��b�����	Ǝ�=%�T� a�"��D�gG��X�O��0ph�Se������(�p������� �}Gs7+<��"y���ʃ���e̘۬�N���|����)��B�C�?�+�ng��J�nn@���5��U�ɢ?��o^kU�0}[����7q/����Bߋ��7%K�|R�HݼJ���n�{�/��o����eK��R���	�}LIUWJ�g�@Rlm�/�y�X���ݘ���p�������4�aO�d���d���'z�=�B���Hzы�s<�k �i�z�M��愽ޠ��Y2K&ؤ�oV���%��Nh׌K�	��(�n���2������m�+e����l��6bNg(��foE.,�����d�J@���!�n�KMO���;6>��[ +k�[����'�[RL�����܍���,փ���{!,��L���a�D1�2V7�ge�"eT,_���?���k��E�!�i�����&D�g�ɲ���5�,��g��D(��_gº\
	X����B�N$o��uy��������4Xǡ��G�(h�f<dK�b���]z�Ԝra�v��R���;R�� .c��� �񢂓iӸ��kݟ�kE�\q1�f7��Y�pW���f�aϏI���op�.;g�V
���Ҳ�M�֧/gT�	�o2�j~���&6�F���#�w�G�6.)��1	�*���R���}z1(M`8�}1����\*juC��V��?Fo���P��C�E|7zgW^��,�uv��i�������t,���^,'�:���H��JX\�M�M���Nr��ua�YtB-S��ِ�vN6R5yD CWmHA���nj?^h��
c.+��I�r�p��٪MR���Kc-kO�T�D7ţh�ȅnx�)��T��Z%$��D�f���f���4�&g�wW�YwX�U�/�v�pm�atf8���-pzH:�h�m>aE���߸�f�:�V|ؗg}��Rϒ�«څ�}m\_YЖ=��X��p���.ОK囐O��CES���6�S�C��{��bo��->��R����#� )�t������LR�����+�:VX�����2��sl>��a*�# ���A�͕|�8B�93L�J�?񗋿��ț)?��;���YYq�3}�CW��w�,6�}��J}���;�}��D��U��$��0n��j�jm�d��A�6 z�h�^��ը� <	�a��#��;�Q|�����.r�2�C>T8�K�R��xD(�9�*�!��~��ӹ1;S�o���j�-��9:�i�-u�9Hn��؍9O�;�O���˗@Þ鳶R
@�W��3.�5r
U�/����,\Jtg���,OW$��G�͒TT~dy�e�#s�Y��͇����0��t=7�	ɇz����y�o���l��=k4]��/�[�/�"u�W��:NB����.�Fmζ��J���竡)@���^� "k�hfno�NB&��P����ڧ��A@��u�T��`�<ab���!����w"���2����Ϛi�UK��8�գ��~U��DH���b;_��c$��թ�#��p>��[�c���FشԴ��Ҍ�b���s�EGY���)��;�� B�r��r�	��Xg�}�����B$�(�Q�YYQo�_nc�U�ՈV���D'�9�Y_]"#�����Ox��
�f������Ν!]�k�!�ÿ<���|�;��i���U��
�em�!4��=Qb���E��~X�����Ex�k'�i*���5�~�����s�?�ZśS�h�\��U�u�����)�[�ǣ��6����r`2��ҫW#�RER-r��!�Ԛ�f��U<��(~A��̗�������׼�)����R�y��Bj�I;��Է��Ԑ����F�7��,47�lѬD��-���^��<����	߱�٠Y���	>LJ�3��YiM������d u���*7B¼N��3���n%l!y�\l�ic�0�&^�?�#T�ݓ�˼ �`+��A�+�UA	@���l��~�}�7�W9J�)I�q�y��3x�@ٖ
��=?�/-�P�����WרA�_��G���ZA�5m]����L�|��q��&.�q5��U�^(l�ÄF�'Y�N�]�O���2��n8g$�ӆu/<�-#����� |8���iZ�o�ACq�V��O��&a���{���n����ٽ���u"�Qڥ�,�e���E8V�%N�����ϼ��c_�
� �|��׃ ͽ�wK� tr��ݐ2�(HT�~�b��8�s�8�iE}w4�OY��T0�NZ�k�-*�1^i�d$94	E��u���;z�6x�D�d��<��'���%�\ @x`��|O����4}���p�ޯz� dw�����:q�˽E}�:k+�kh�p��@KH3\r�}�"�i}��FH�^�D���y!�7���ͮoJ����2�_��tl�ߗ��R�2�g- ����k����<)n�JR`�����!io�P����	1�7���˃�����B�+�l�۶��/�Ѻr��y�� "���npۛ}i�W�f�(���s�,�%�sA4�!�|�$�^m%n��<bc�:$!��jH�!��~��٨:�U٣YO�<���]�`�I�q�ʦ�[��N?�dE����,�r��[1:7	j�Pq|8�w~9JQԶin3t�r4c'���gJ�q5Y��w���o7�T*y��ڍ#YBm�E�z����a��G�"�&rgp� �I�ZrW�	�Y߇>HZs[��k��e2�<�ww9M¢	�pTɶ]m���P� g�g�Ee�o!v7��@�ƯN�O�-�Ȇ�j<;d�<�"�jt����2�W��s'W�����i�Y|d����?Lȍ��w���u�U��?��}fj�jp[������A'��o�Hi�*؇k�v�$�p��,�i�n7G Bc�P����(���N��>�[�3���IE��y���Տh���y4��j��%'J4�w�"�ð���S^Q����h"s�ٯ 25���^׿�_Hrk�4�r)2.�F�/]��������a��-gJH
�Q�\15(f�|���Id� jYYVq���ԨM���9b1#�;�4����.޹�s)J�|���?*�|��0,�L��>����9k�m&^ˋӎn,a~�6���p�3S�<� ������E���M��+v5�+Ӣl��[��&O%-�v�bh	�r�F�#�pF:�#�u|W�
TV�ncɽ*`�Y�C�{�s�t�y�?.�[S*b{�ݰF��IMq(v�C�9�:��u�}\h��ה3D�%��J��a��j��h�$��1�#9X6���:$#d�^�����U�yTy����/�s��.vw�0J���RX}�����Q6^Ǚ���!�=����
Ⓖƺ��|Nnbc>�8E��5gb�J,3Ѧ=�'�U�\�P'�He�/�xs�{�9�������eǌ7���qt����R2��jf���s���s4%,,�
�=�kI-W���:�Bq����2Bї��ȴ�j-��^�(�`;�Glk������`�Ɠ��<]�^~��)��s�H���R_*���,��V_,�͂���ta׊����K�[�|�w�|aD�92 c�g�޼ܰH^��a$:Na��X�ܥ,s.-c�q$N�C%�@λ:q'S�3E.�ws�t���Zg���b�v>eU���z��c�9�}��j���p�b`,�`фO �%a2�wy��&�tt[��,\Hba���&�p�v�`�lڸ"�s|�"���	H��%gDN[M�X�. p��x/T�:����u�����\�J-qO�=/?�-"��3'�r{�qȡ���E@�)W0;��5���O+�h�U,�����	�PG�(ѻm�0���B{����>T��l}EjgE��'�1�ճ��ް'T �� �q�wPñ�7`�3='��#F��������ZY[Dw�����F�L��U+
�/J��@	b��Ӝ��܈0J�!\ǅ��yK�B�}�Y��/:,�L��*eeʼ��9R{z����%��H�!�~��Lt���i8-���L������B�oY��$�$��1�N��;�^v�z�G~���%�ѐ�"!�'�2/�Q�WxCɓ,��Eh�LA ����x:�ed������}X-ť(�)sB�]�g�����_Vb�HV�!*XK{�>���,�U�Y7��$i�{;��*�[�c�_��{�]��w!�ހ��`y@�D��ͰA1�mg��DE�O���'haf\&]<Ava��;�{�.2���8��lm�������/X��'T>�C8@����� el���,�@vU{��������w�&�`�I�mP�df�{,E�t`���WۉW���Y�sd�q�-�|�gհ�
�$��
GzbMV�"U�Plw;��U�ͅ�/��#~�Yk�� �����;pom\mӵD�es���=;o�n*���_���
\J{V�,��ur��ʥ�U?�J��������#_��