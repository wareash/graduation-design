��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jåا{�\�u�?߷�dn@6�zf��r������;��r)]����c��`Sz��/��09���b�Xb�>ޒ�����e��4�t�y=��M�c����zT\g�HE���mԉT(	'~д#�
�3�#a�Ɍ�*��s�LE�����<b�S��Z�k"B��x��63�	� ��������'A�ԯ4����*�u	��;Ck�$.�́ʗ#��h3q��E?t�=�,[U���+s��:�/H}Z��X=��E}�c�n�8�8�FJ�y�*rh�r�G��y�m�!c˳]���=�I&.c�߰F��]I'�A6�-?��\�.Lz�eg��40����؏�����xM�%�V;鉎T7E�����O$'�}���5����&�@v�;dsc�h�;�C�X>�	,�leChك%���8i�H�9ԡZ�a��:��Z��Fc�O����(��4�-mY�oQ&i�R��4/�a��%Wv����5y4�Ȃ���@\��x����/���3�N�Z|u�l����5�	���#��qxYuh�M4�ɿ�u1�+u.������~2'i,R�H�ZB\ڔ��ƕ1{2��o���i�����˽8M�r1�e�[��/DI[x��^���ةK�������"J�P����b�n775��;�v��-%��t���,�YE��	Ҧv���I���Z"�1£�;0�vb�K��g�
�"Z���G��uQL?��e�����趈�hE��k&A���(_�d2DZ��?�|��@ƱO�Tzͧ.���k*y�K�Kª�cL7w����C�� d����򷯜�O���Tz_�꺝�s��r������0_���\>�h��]8���u�^�P�E;�YA�7��~HU0�jsv���O�b�G�k&�"�������s��ܞ~���|'�<��-G5N�+��ϣXQ�\�؜�l.A��Y����j��z�^��d�3Ӎ�96r�.p��wz=���i<�U�����jÙS�B���Ȯ�d:��>T�=�[��M&���@�WKɲ�;	�����?P|4&�a��H>�V�$4��>��a�t�)ɹ<w����b��<��:-��G������õ�p*:=��B�Ie@t�xD���4��.�g�R�2������O�FZ�*��&~%���Z�^�;~�79ng�.��gK��j'n�̔��֦�9��Z%o��y>�~x �	K�Ӑb���r'
��U�Y��������h��m���	.R�J67sv_��)�qC��zaC�(?���*x"ŷ�Q<.g"��<m�`���$��j�[������蚁PZ�߸N�����g�z���
iH�kK'���9�YO?gP}/[u����c8!��6Ѱr㧦<��*�fH�<B�;}x�Nr�+�#���[`�>x�z����y�U����^۲�/����w�&h8��~}�S>��Gj�f6���v�F ��U�;�a��
~¢�������k���'+�If]^�2SS�1�9��0 [�QN�#�ʫo䄀t�Ql��~���u>�|�ɻl���b ll�i��ͼ:5���\͂����VhR��7�B�D{��ߛG+��|�x$$${Nnܸ�խhY��	��Aꬆ�.�^�?�*��]�]��� �U���}h:���B]@�	��n�#'v��KZ�6��Q��3��G�G�P�v�:9R�,�1�x�cG[�Ź5�8����y��HZ:!{�	��M\Rt� ��;�ٺjv�@��E@��O�xFew��@u�2' �F�/�,��p�)� 8�&������U��#���]���#tW�Z���f���P��o�14g�����B�v���W�t�e�c�.J�㣷jEA�9u[�1\���.�d���`���/E �t�@X�4�ӆ��\c�Ґ���de��G�p��.�5��Xf�b�S0e�Km�����As�KګZfڅ� ��4g�G�l�K����y�4�����"	:X���� ���:��d��^�sQL���M�6��CrȠ����>8_��6Vmw�.�`�Hr��sWm�M�=1[q*�����5=�@��-��)V��W#_���/�ak+���+;:R�z#Պ	�5�����Q��b�#�C���{l�g����K���w
�*����lߺ���=cAz�lC0r'%h���/R���U�����I�ؖMP?4�Z������b����{N��^�+�Ni�ӝ��a���C�߽����9���t������e��
�C[/3���l��QI���ܘ}��e���[����i�R'wBjC�_��m��Ս>�mn���>��J�{r	b%�G��{�iL�ʢ,�/�m�2uj���CX����Wc-a����`njzv3w ��|��Z���_լ���ri��ĺ0Ӓ1FtM��ku�ٯ�}�>g�ܗ��e�A1��"�A����|�ZB7��a>l4č1r9�-pgK?���(��g!a���̭(�ݎZs�A�&�����Q�h�3R�@񧟪�`�^G ^P�~��\�e3�}�WL�����e=1�{_.�A�v��lk,�h�xu�-3m���N�Uc��V��)��lb��9����.1[+p~mOG�6�U
n
��b��a��S���� ��	�9mwA���s_?�֘U�I�Ȧ�,�6 qv4?=�	w�ma��ȏtF�t_�?")������i֥#�g�q�0��W�x��s�rk2�4�0��D�)�y�6Ͳ��.�0C2*��7~�-e&��0j�E���Nv3�ΊA&<9�C"C趀)n�f?����y#�0q�j߾�=8��A,A�P���)x�ET�[�>N��@=CI82x_V��Y�D�����^_�KM"�'�;���L6͡�F��+'@�0lq#������N}u��P�Ae��^~S����= {��)p�g�nnk�l���ɰ�T㤛�Y�5��?,U���	z����F� �J���Ӆ1/��w�ץnQ%�)�3���("5�L��9?�d�ql �t�w�_�"u�{���3�	$&(���#;��q�����'͏!�8���J�,4�Q�&��vX�p2z�eָ�zY(.~1���9�"��V��U)I�0��޷��"AAH9
q��`]�6�����G*�-����g�-�'p�6�k�棓��7�&�¹y��q��*J��˶>�x��h������ź�d�����;~������M�> � @GK�OX��"�v���7JmZ��Ր�1E�f��q�y3'�V�] x�\�g��ey�	}%��J(}Q�����5A�3L�&�3v�.���,�_
o��U��Q|���QB�c������I�gw�7$n!�	����T�������s��#Vd���M�)�\y�K�_?πD���OBA�+��[��թ�IE1Xy�h-��i�$��X�0��U�:����LX�<<�V�VU���>�Z_E�3�
}�S�,�
n��$�8�m��2�E�G���Cŋ��5&@�3G36�㚭`@���q9�s�uB��b�~��!h�׸��b�O�q�Rqx�G�)�����f�!(��z�[�(�t���?�������h�"��on���� P@�.e"y�σ�H����!vܠ#������� ��*}�X)�3��Ǌ
�ۃV����k�~��{�͘a>���,�f�H��)��g�Q9 �c���y,���Z��VlD��n��U��/{0D��r��W�DgXO�y�U�]�d����X:��jRyˊZ��w�[���6���}-��mn�������v�P�Í�mk<,�7	�=�dEL�6�ϟT� �$�&q I�<G̻��U�^M�'��� �'k,�6�Yu|s�0����M��f���������4ݟ+�ѭ����٥�~��,rg��"�6R��/�fBLS��^��i���e76Bh6����[�ث�|Sw�P�7��zha�����قx�Ɍ�	hR���r�n��!~B�������|C{Qв��|�e�F�0�\_��6b�C��k��g�_�1�^�&n�o3���h��Kq��"����u���<�Bݖ�RI��j�[\^�BO�t�e�c�)�X���x ���{jL�W��ZԖvo�VPG�jm���U�	:#Q�O�g��i��I�ݴ������E����+��Ж*-�ֹ�����������nzp�[K.�6��UkF`_�*���(q3���A֔�$�=Ԙ�������ON�G�[0+�>���	�m3	6�^!�6ژ#X�F�
)Gi��ۛ>|S�.�+���#y5�:�G!���A��꼎j˫�H���8����ur ^ m=�����"��f��yE`KoG��Ӡ�K�e�A'�4<O��:k� r�'�vc�P	�z0JoA^UV�P������ʟ<��v��b;aQ	�ȶ={{(��qp)�^�Yk���А���yU���p2�&��c�B�i�Ο�w�f��X��SA��I�*��?hB�N�#�`�������)f� �L�y���ɖ3�9�_��#��h�/�~O	�����
���h����޾;=ӎ3:[7�d_�C���0��3Q�{a�����t�$M�>Eo�Sz����E/��Se`>��z2��M�t �P�*5���5��O�4)C�eC�j�6�vZ�IS��Hcd�y��@���7꿛|A�bZ"��9���3���z<���v�JT����)�U}ה����>�9��{E�.�j��_ �كKQݳq1D��7�j���u*���P}W%u+�ZO�D^�5�K��j.���Z�K�S��~N�H�Buޏ��'�@(4�=S�"����\|�Od8��P̬�vJ�����S��-3��0�N���me�}(E�<����E��gJ�,S٫��u��]���V����m���5<�_��|֌���%�^P�9��B�&JvU�gB@Ph��kH.�_�瑕_��9z*�þ�/�h`���hG*�-UD���Y7�z= (ձF�2��<A��`�"���͊!�������g��w�.�!�y�(6�����Ѡ���-z��v@�r�T\2�qn�`�y���h�]�nh�rj��+����L��=�����?������h��Z[��d=j�l����~@�b�f#����Q;����\�;���<)�7ӿ����\|�{��+ٔU=�����V��e-�nN�> +m�v�����ʒ��x�Ԣ�2������D�E��j@¡hs ��+�`�+c�~�u����Lò�,xLg�N�e�,!_Ǭ���'Z�n�&)��Ѩ��)�gl��u�����ꛊ!���Yo�!��~�C0��g@�_*D��u�^��������<)�b�`��GT��mE+_�C}Wa���jD+�N�������:��.�䂩z!����{NW�!C���a������(�ͯb�8���y��4�18�[#���`8$��~E,�I�)� �ր$\�^�}x�$���LO�)�4�m�+'�^�8�a�!:�-�
��Wp�++��HsB��jV�(`��$*���xz����S���5R��{m�6�<+>E�1�埦�J�ԂQ�t����gqO�`{<�GlG�!+B�j�GQ�]�������b�ӮN����m��p6	a{s�m�y���ؙG�P�����T��,-����ֲͩ	�N	>�����>P=1r̍��E���b?���Y���Sǟ_��aܪfI1&A]����*�Ha�_T��0,�/�D�mr�^���.�`�0�u��}�k2GF�1ց�oX\�T���euR��N���L�Es["7kj\��)'q�X�`�_�cTLW��Ux���!F�M��X|1���y���J�I�X���ӭX�+�omiz�����{��X�j���)�����l$b��r���v�� �a��Υ���\����c/�����%+�BpC���V����7{�CS����]s��I&�����ᶲ��1�
�?rS2�`�$HY����C�������Z����=��)�_`�oj���:�Ζz��GsU�B6�H�b�
?:���%�Y�ڙ�Hc]�'s�r_.�o�]�1�nd���U�&������'k��H|�V��8�������$?����{1�2����Mک�� =��:��.�w�*�k�a�r��*P��K,iŽ�n�pPJD�Ӥ���pP�.��)���P�%��r�B���B�{���w������_+ZA#Q�_�{���C��'V�f%8R̳ྐ��%�c�<�Fe��`��=���9�u�g�9�NH�,���^l%���ax�g�������\Gھs��dH��4Ǎ��U������Z�:1�y��|���fא�#�m<v���]Ԥxb����r>�gO�Z�,3�:NG&`T�(O!�4��d��I���"|g����\B�9YC�6@�\;o3R��]o�Ns=�X[n�X`aK�����Vw�n�[T�&�J�t_W��ň5�&�99b���^^T?(ƴ�i����'&I��?�	'At�	c�6��2vl�aX����`���}�C���c���6�T��ǧ��²�B�Mڕ�J�D��V8'�T���r�FUs���	�8%��	4&�pY4��q���)1Ƶ3��Zur�����6x��/�r�`�l���7��`��	9��I	��t�۱Bz�/���E	��U?�3�,}+���X�Vm�u�8��i��(�q�g��j���:Wh8=�f���	E>x��G{���!�oǇk��7R(mG���$����}#K�ܞ�H������ |o7��T��"�r����@�q~W��-�i7W�~��#����WN7�C�-Ajּ�Q�Y��uxȆ�7'�T%���v����'K���e<�����`�����!�{��
��p �B5��rn5L�;f0���5��Np���}$�