��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jåا{�\�u�?߷�dn@6�zf��r������;��1��B���7$)Zf�ʿԖT.i����Y=ұ��ȵ���,�<�9�Z��{�`�V"u	�t9��ϱ�G*i3�ܽy�hq�T��������0'rލA��y�?�,�=f��FD�8���X*	���|#��N�9(���ְI�`��CwQH�d���P����u�v�f���G4dr�$Y:r���z�&�_�1�m!�x5�9�X�;���b���x�<o >�7�{�m�>O�Wq(BA�3���)�/m*��ظa���E��2�ɢ�-ڿ���ea�>ߋ�'�o����w�i�KY�3�����P̞OX<�ބ5P�6��0{��
 R�Esn{���|C�;wb&�;��9kC	ĕ�G
�<7;/^ T���+]X`ݝi�	lԃ_��լ�L���o/�o�Z�G�&��O����a��h	���!������6�4�:��x?|�%r�:�D��h;F�qt�;�9d|0�}��"�>2E<�?�D�L���n�^���i�=O�U}	�������}�W(����<&� 0(��P��t?��8���Zm �'�R�����������l�Ö��/Q�N�X9:���<q��c�'�|RX�ڢd֧�)om`ɶ�d��C��)ĺw�g]!�-G�zwJ����_��K���`�,�����n�92���v0��/�+ޭ�	�tr����N�w|o�/��L]q9��O�>�*#:s.��>"W-$�ײ��;wfcf�\��N4�+nR�A�[�#�~�_��O�n�O��ȧ��{�B?�pZaJ,�8mM��L��P䍦�ⷀ�R<�HH�L���N^>��SJ�SAa%4���{!^O����2��¥�B����^i*�x�L��
�=���J��~�J/�L\���q{`X��5��[��^���nl�[�bh�sV��%�RȽ�#G`N�ke_M�Oz��(8�-�A䷗�r�IW���a��-�I��{�h�����Z�"�|�����c(�k.�0b�����ۢ(�h�pu@�=h_m����$�Oe�G+�Ҡ�m>k[��:�t׆$��ˮ5��FD���VN1z�0	Q�X���%�"�}��w��}��Ӑ1^Hht� "�G��E����LOJ(���oؗb[�R������rG��G��V��X�v0[� h�T#�M$Z�5�S�qǣ��k\;�Ň���Qql�����k:������� ��zp�=%�R
�F��g�&�ff�#�}i��s�ֶ�`#{4�ñ:�\Vhy�5�h�7Z$.�F<Exb)&���_|�"0h��$��	&�u�ϼ������k�?���<Y��I��&32p��Hv�6��J��4�U�υ/xO7��l��p�B=�2��řQ+��x��;����b7qyؼ�O�	ɢK{d�UE��9W�ӯ����^�*�	G��b��#.fa���Q.pt!��xJ�ց�K-=.H��+�G��1��$}����CdY�eD�}���mÁm��nH5\�ʳ��PL����l|�!��>����Z#�=Uռ2rC��jxk��6�W��ٞ��:ߋ^���5 �����^��3E���|�*tb�:����f�%c�I����p6��'�p6�Cl���}UZcc5y#E%��8�Ꜵ��C ����x��}!"�F�#,Nމ��q}l��2}ׯ�B L��'����~>�d�d�X��#��F"�'�n���.3fM�K��Q]������/��
�f1���~�.����1�N�w	�iEAt�,9J:9pw h�u�^k1j���G���-э��2]Q^��|��M2��i�~�Ď8r�vi'���5>��ƺ�Wkʵ@���NQ'�
ɀ�PT��6
���A�Ǽ���dԖ��S�V%�7�H�Ԁ���ܯ9į-k�]���:�>F�ʬ(�Z8*�М���6�u�����0p�CFq��I+M���6�c�	�d��q�]n#�>:�6��:�<Y � 4#`_��9%	����s`]��l`�<4��p�b�z���P]&���3E��d�	���Y�G0�'�]�W���N��r�c"�]K̂�n�.P/@��F�x�}�l�h�ka[3��b����Q�����4�t�,sϹ%!	پ{��bz��S�`ד�Z7�-���L�Y������t���)�a=�x_��Mؓ{h���/U�z{�,a3�"�Jsp�Hb�T����it����{���O:��Oj�O�0����H�j���}��������~"]���p�hJB��HEM;8f����!3����_*ܡ���ǣ��TN�e2���R�3P=[;gga6k-0`�-*kEk��0U'I��R�)Z�m�WG����B����#0!1=�<������PV�t�/� i�[ѫw�d�t�oL�b�4�o!�p���R-.��l�%0���M�d� (r�YV`)!/�NY]�2L!�w%Lq{r '��m�pU�Yf.��>���'�:!�D���X$�y���P+T��k�z���L�e����Dv�i�f�g7����7���Cuvo�b�-�6�߫O���P�h�<�`��[%�&at1���BS�oӨ'u��t<�ׯ�aI��鞷���~���i��sυ`^o��;�Z-����Ȫ�c��t���'��J�Mu��=Z��I�0lsK��'�"��5�A^��e�$F"RjN����M�Ec~�Eᣫ�A�[]��cx-�ډ;�Z�6BoUN���|�u�?��K�?R��U�e]?(t�~�;�E�
��PR��1�TUs&��̩�_D�Z���Y���=��ӌ�v��F��4(II#.>	p��S���3��-���������#�$�?�+ �dA��}c�ֻNyI�a-��
��W,��4I��2k�ጹ+�7�F��bl�-R��[�m����̏��p0��*��ph������������4g����2I�sض!�@ht���Et�{��l�Ѻ���ˊϣ�X&]������kiʴ.�Dj��k�<���Ml������6=N����&�J�=�t��7��𙷯v�F��ۚ3P�$�`OxDo�~}��������w��S�53��15�/Uc�k�
!�$|fLT4s�꣍N�Dن�ǖ,;܀��q�-6Y��%ؖ���B�{o�Hٜ�3� �����]D�tt��B��%LKb�u�!^���=ۻn�1��3� �l��ѹW��w#x���6�%�lbG�"�ա��Y��f܎�&(�h��FT�+Ϭs�g�X�&�Z�@	C���������Vl�.;��9t��[��'�#���4aO�ґ=G9�1�+��9������8P:Z�V�5�W?'��\�ӣ%�d�
�z��W��������~�S�P���0PC�,^7A�ՠ������N�M`���O�D|�vF)0�#���b���;�DpǌI��x�rL�i>����@ol�3�n�4<�,���ī���Z�?�q�4��U^-ҿHu�i-�@�����~�;:-y�o��3�R�O��9�g{�1��>�Hzf	�q��SZ����r7�'p�ϭ@�bǅ�s��N11^�`B�_A�\�h?!�����;��H��f��c�;t��$�.b���w��@5�F�\���[Gڡ��l��	h�KǫivF�D��R"�z������y�c������ay�BQ��g��ˣ?�� �#�p���>9}A�42$m�ǹg��y�9��X�)h�*&��
�� $�+��y�`�|�+�
y�Z��JR�i�h*�	o���|�� q��^	��+O�@�QU�Zud��ٞ$�y�X�~:&\Ω�6/���͂{T����"ez��f��ϟ.<�~��M��@�H+ynx �;4��ECZ��57֫6#&㮬����,�^8��Oō�����zc�������]��@VaJ$8�����2\��M��֟u���:#]$�9W��П�
@0�W8�T���W�Y��ƫ��)L�J�!�f�G�JO��@V�F�Ur���ת�0��qx��~�w�|@ǖ��u��*k'�WT���mp�(�MX"�Z��њ��o�V�I�v��h�G�n�uL4ݰZ�^�{���I�F'��k�h�3�ǤA`>
Lz���݉6D�Q8��U i�Ƞ�:/.yu��sL��e�ɨ���"�����Ǉ�޶�����)�eY���բʁ�r��+�� ,\�z���ˋGLF�9�!�Bh�l�.0�����H�����	�a�,�v�]����?�ֹ{m��F�_�*R��U��G=;�	/kD�]�1 t�*D�S1��{�w\FO���Vg<s�hL��b�t��\��'d�Fz�So��m�^��)P�jQ眍�j�*�3Q-/cL�67�|Q჊����q��dc�RS�Pٕ��q=�m�{ٍI*K�*��<�(Wgu�&&D�Hsx0d_�����,��?���y�����������������m癈(\p�Jw�9�n������<Z߬��B����%~h�%>tߊy㇗5i��'K�B6�?#� 7e��9���b�M�_�D����7���8�]���&��w������o��6}E-�>���	Y�\��V��q930��L�A�ˌ�3�x�9��T{G��>�w