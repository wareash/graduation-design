��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jåا{�\�u�?߷�dn@6�zf��r������;�amb�����_�P�TO��(����,��㵸0+d��`-vc�5YX~h�s$��4���:�X����V�$�����n.lE�h(�Jق����h\�P�s�7|р������2�l��G�G!�'��O~���+���F!�-�~�*�_> �[[�����N{A�O_�Jfޤ��gQ9C�N#��2��[q�R��'EYeE�y��<C E���ǟ���ñ{��Ǻ����9���p�̎�:��i�O=�JgpwU�I�U�Jɵ�/�&�9J�j�w�.A����ە�G ��Wd����RB�ɹ]�s�}��5���w���p��=����W��t�D~�->���S�Nۭ'"S��p֢� Sp�Z?`�Ӆ�L�8|Pb+f�VNe	�Ž��z�Ŋ��%��NM�4e��p�,g���d�;
�Q�Y��{DwT "{���+\>�<5@\��{�P�3V��E�N�=>��uL���,Eb`��LZ�C�)KV�z��;�(^=�|���[ݹ0�h�ڢV�OQ�A��j|������	�ڐ#~>�m�\�T�`�H��ː)+1��Z�x�>��"�6"���ڪ��<�s[�����l=1���y�ۛ���1�L��r�ͷ���,{=b�fh\D��
wc��P��q�&��f�$I��˭�i���� �-" �s!��{;Ù�ڣ��%.*��
�mQ�=�w��i��[�w���a7@�Љoh5O�
�	��l����[�0-���Fwg���O�d����v��j�f�7�}ͨMx�ޒ�I���[B��`s���w�%��k�l��oG���@��9o%�f/���lv1���p��R���= e߆\7-2���
�'�R�X��N���h�>z�Rư�10̀�e	��{v�����\�e��í+BRw?Q�d��˥��R;F*JR�[���C,�	�'Ǌ�ߝ��BۏC����%8��"��j�6dvt[�d>`��f�������}�ş:�vy���׸^f��x\�@N@ʧݵ��Z԰�;����Գ]~�6H���Q�AeД��n$x�]4�В¹�ݸ���s���ٕx�HQZ��@{�l�c]�n4E[@���弣 �TX�v�����#���,����ԫ:�'�jQw=9%��/w4]l�0�@���M�u�{r�g<Lz��;ae��c��K�FvN=b��'�������-DDW[�qk��O�օ+�-M�(�����>�^�Ƥ>�;�W�95�0<o�>~�s��=d��;��F��t���V��ad"�hr�d�q�ͦS7�}�8�c^�qc��r����|Z˽X�g��Y��8��6��F�$t�Ӕ��V��z��a�2^>zx���X(�x��^^y�/��S�H6��\�8��S�	J!���$�[����:eW��W�RQ�x���n���T��¤=�F}<A Xަre$ӆ����@�/�]��;c��y>u�r���6��z`(ت˲.��5I�}==f�C�tM��D���_�#��Ԣ�:�t���d��%��>�z,�*�y笘�S?�ퟨ��s���Fj8OWy�G��k'��������F��>�c�|��T��Pt�=p���pޅ�P��C%�0���4N���q�5^�i�IF�LZ@ �G~^x����u��T��Rl����r�!1C܎�l��nr/�y޵L�zka��E_x���DH����M%r���������c��e]�"�^�4����$�*_s���
aM�s�f5IH�x�C�!$�E�%��0�Y�U��3������a�?-�sN��3(��M�z��Q�à���2�JH#��ǿ�	�$)yJ�����\���kR�T�'�v6X�� Lq�(�.���i�щ% VˤqIU_ʆ׳F1՞��nX܁z�E�.'��,f	���s\�����b]�ό�9(�S��m�q��;��_�i=����{m���X�Q��`�B�k6JcrM	��un��z#f�����n�kkG������F#���4_��J[����ԫU�`C��W����"�B���˼�a�6B�*���)�ㅏ3�ͅ�����>e�] 0��H@X����8��x��M��t������#ܞs����c=�H�=�Z��u9�6���IϠ�?��6��ldW<��:�~�VS�6I��œ|E0��Mݻ�l˪��sf`M5Z@���%H��%ج�:��Ţ���*�M2�R ���hK�f|Ԕ[��c7�ޣ�I�Y�	��/U;A��2De�d#/q'1��R�Bw��!15y1՝��nd�B;�vf�� �m�j�]�H�Y0�f�N����%����c�C��D�C���2ɽd�F���
>��,xz����rKh�8�I&#��
�˶�訉o 4;���O;��S@�] ���CR�d���H�洮Q���ޮr��3�&vrXS�3�'ʛ�'���ߗsw�|]N3[�ec2���_qJ��rt���[(�0��l[
\�]Z5w�"U���?�e��$\�E�����%(�k�1rT����Y�֧�~��IG�s���&ЊqY+&}姑�e�HP�PӤ�&����G�Fb����@�Al� ��[�:���?��6W*.�p�l��n��,փ��ȧ����
.�Nfݹ6/�վ��+Ԯ�3|N�م��6I�M�%_ǵ�P����K�����N{o�1�� �u����İ�S��>P�����n����Uv���&���Vb���y׻>��d0�4�f�(�������$��]�Hŭ��a�����ۻ��1'�Җ�l��A�S#�5�"��:{LN}��kY�t�O	PΠ�B��P�{?A+$�
3.�a�S��wh�l���N��Z�S�J�z��WҮ���3�X����%�f\eZ?B�K��*Oܴ�-���=�!�Y� �,�\����b>ӑ)�����EV�$�؄����Se��fH�5�`�"�ӢH� L�v� 2�dW��F��~�7a,4�%���\Y?N��P��Z���sU�k� ��3.��r�RJ*ŭ T�k݁�2�f��C��߁���E�����f�x�c�Z����~�[�Qr�wQ�-��f?���U	l���̀��h�����8c������:"8�ٷ���ª6v_��D�q¦���d+��ά�w줃o5�Nb�nR�M��G��-��h�Q�+�u˂!u`��} i<�k�]�y� U޺���P���k#�!+���߉�b�8����=Bm�y�S��s�W �;�*�?�؛���2Œ�^�����T9��t{������B.�LP�����2�%��ClV� ��,0m?��uZD�I�o� �F���*�@�g{9`�@`#O����5����{�0>k8$xC�{P3?�~�J&�{�C��ɉ���GhǍ=�H�Z�F�g!��w�th�f㔝���[�����oZ
����d��X�6O�xF��%��SԌ�+7��BE��,���^�YD�T�Y���3V�G{F��Dnاee�Z��Ÿ����-\cf;��F��C�P�9�(*�΅�)E3B�VB�=����iB p��a�{�:*nUd��?d
�c^�ʋ6d���,5�Om�QҢ�?�zW�0L/�S�\o�i���g^$���Y����Yt�H�v���c��+Ɓ��꫊�6��D��y�;��G�6e�Li	��<�*��Ń&^<x�k֛�LK�hQA��Sy5���"#�������!�_�"�k\�~� ؐ� t��ۺ���� ��D5b��2CD7�n��P�n�Z�a�����6�p��H�`$��c���n����H��Q���A��������/郼��B�/�{�X0�FHD"�s��P�i5�D�%��r.D��79?B��N�������-)�R�������Nc���OR8�o�t%��|p��<��s�q�;���]B5Xh\�kfZ�(��PP"�Bwe��0���n�i�:�E�?%��ӎ� c����۲zK���`h,������4O��w��ж��[R�l"w�@�����X)�&ա�?�M�5��� N���l3��#����EӼ�-���ֆA�K�i)�ސ���ĿZ_R�^���wQzxԚ��:V�25�@98`Z$�pe�W��/� �<.�]
�D�E\Lc�	��~�/��i�i��>,����[�{m��(��6���oOe2wl�%Z�#x�_�C1��_ل����~ڵ;H��S���|�'~JRJ���b*�y�C�!ge�T*l�9���b��B��VZ�TD�lMH��Iy��	�sȤl۴�5F�b*0Vs�6�$�2�x4�P���L9Ņz���(i
 9>e��w'��4+1ՓQ�w_f9�d���U)a�8�4�b4aJ��Jĵ��q�u�����y�s	���Whc�$l�'�n*����S��N,��,�pk���3/�V��x�e7�\%t�_���1�Hs{q�������W\�j!i�q�<�vp��:Y˹��!L�S�B�iV;hlR!?4_� �ޮL�I��i4ph[��8���M��}�A��	�����+��g#f�p�c���F����{��$�:��@�t-g4�_�L��B��f��c����i�;Y�$��%��/64����3|�a�|�N���S����Hך)�5�w>�����X�R�tu ����ǭ9ó)����&����>AG,��i,4C�J�Y�7�cw�5EJ�|M�G��9��a|,E�Bv�Kߞ�x�`�22��1MŅO>��3!�+�35 ]5� �8����Đ��W;�,�,̤�(E�:(V�?�l�c����me����`�f�hB�?,�-�\*?G?��i8.����08m���>SE��9U�қ�W�Iq6�GF卽s�U����V5/�7��'�;dc�%�	r^i���֘�K:�!�Q�-\��4A��E$����:`�P�erPy�;^ޞv�o�گv��O5V�u���I��B�&r�-�� ����_���H�
-��������	Įc;g�_;�4���*G5A�T�IЦ�W�*��1���J�v-�<��F��y��]1��8%�c@���$���Y7�ҤM��"W`n�<�vb�X�.x�#��c�kͬ��0=H�2��� V�G�����D=���$x�]0��%c%�K��y��̀�c?��Ʋ�:�_q��7mc��-�������q��xm� �Os8墛�M{.���L�\Lu��C��(�MkS�7aqq�9�7nڳ�r�� V���3����À��'?�e��4[1|��#�͞R∂]<�@=飻O�c~�eX���~�]yM`0nM���A��s�w�`�����撛�ظ��m�0JhFȹ�%��>��l��ޯ'W��n:]� ��z��� M�py5?c��9��&m聫����״�@
n�кR,p$ne�
���%�EZP=uԔ
� ��G�t% �Q��|E)�b4x�@�8��#
%��)]b�!���R����a)�S��_�؉��Z�[��&�&��KÒ�[">�1��[�C�D�b*�V�K\_QB~��>�e��̮�*(f����"������X�EN�}���@z�γT������B���s�cF��21g��t[�v�Hޓ�6�OB���y��U?|�j]|��NB��s5VN}�5�;M����1V�vy���Κ�����!�~1%P�^��zE�� �����&���b��B�Sc��bB#�Zx�����״~��녜�oZ�H@�Hp\�|/���	��GǊk �p�5d���Z���T7�L�?�P�!&ʖ�Vh����2כYڲ�������N]+E��谅
/�^i����ލ|ߜ����^��Xߺ+Hڽ�v.��%}����י�j_I@2،�1F[��1X-h0!�/O�ʈ�9Q�+�<����NϹ�>�_���`�.u�tT/^O�% wCs���.އAM���50�� ɚ��PD���4�y����0��] �sܷ�n/o�t�����m��~��yl�<.��pѢԱ&A+��=���2\�K��3�ڕH�}��b�4E��P�"�{�--/	��4E@��ҷ�Q�����Ml��O1�l�$��p��q(�j�v�WA�o�R$����	����u�iN���;�8�[���}m;���;�_���Y�IЀ�g}�.���U4e�.�|�a�i�?�!ud
�����keI��&o-%"�R���Q]K R�,���G���ibL�^��}>��T��i���)*C:A	kECG�g�ʐ��~���=32�85__���Ua��� D�0����:�����G e�Cb�,g��G	Iʑ��y@;�Y�7��:����@��=.��~��L�@_0��|z�d��r�@F��B�������޲U	�t/^#�%}���:RfȽ�HC��],6ke��?2�#s���	I s����Ii�r�X��O��>��!��-'+�������p�@ �B^�j���2�T� k���o`
�7h�5+�5w�Q8r[��A]�_\%ET%\4�!Ѯ��'��2�|���i3{��Y����@C�g/�qw6�yAz��6,=W��]��O	zys�jES^q2yx�=	 M�������~�#�>�ch�o�{Q4g��F����p�&\k�}m�pA�3�7'�{�Z��㈃o��V�[Y�F�R�^T��Fc���}o+�q-5O<�,FW���UlJժ�'��8��� N���F̝�4��
�*�h�륏�B#��z�C9����(
��S2 4�B���E�>�|١2R�x~b������a���q(���~����)�+E\*m����b�/�PE�����g,{xwF���$*2�9�pZ�Hr�������,%�ʴC��xD��FVio�����tܕdo�/�]�|Tb���*nxd�%�R�����;����DkG/2����L���΢���.;��� ";�۶8[�7_4'�����L�� ��1uN���X�w��y������MA��0
y7�g�������Ɗ�ӥ�~<Gi�u���[�v	0 !U�ua���;xb2�/b'?�=��B!��q� �:�4l�A�5�&��v���_+��s��m��yY��&�%i��,�)��Y�f�tY&�p<B@�˘Y����9�A5a<X{^��ǩ��hP�'ةƔ�M�F���#儶@�*&Q�h��i�B�	,���AJE%��f��~M2��Ǆ�]�X��y��3��㌧4�%/m_�fNb�$[;��3��4����ܞ�r6�
�B�z����UBDb;�YAT�9gV���i����j�SF*Q�=y���RN��[�ֿ�}J�d#]�s�Z�`PĔ��T��ea�<��>C�����0Yw�Q�t��H��D��qM8+���+c�&8�x�����f�JFi��"��1q[ee�8��	�D�*��lw�jJ�p�b��N�Z��z�7X�6�N�B�~��Ԋ�����P#a眞�>�x���3g�%e��:c;q9\�iz �Hyd; �@�ߧM�o\��|
M��R9줈.):8ћF�z�~ΰ���t��e�Xb�^���%�Sm���w"�'?��.K�-��;^'����	�iG4TaMq,_��(���0^�drl#hI	k�(I������ix�42�(X�)r�S��@��nۊr��~GFP�A_��Y��\'��uR���鐟ST~�?��1J��HM�Q�D�Z�j�n��l�a(F�������P�an��#4�8m�>X�k�V߅�����ߒ\=�о�/q�$�m>.��:�Je76�|�N�!�ꥷĉ⦳D'��<w�)l�������={@!0�<|�"b*v���_����cq�J�;W�(�������4��:�6�:h�ݑ�i0m�B����w8h����x�m���'兔��������8$�_�?֤XFV���7rX�/�OWW�Vb�y�9	I}-��R>P���e`�����Ax�����bl;��*vڗơ���H��rW�%*���U3��a��>�'��2sJ{V� Q�cWoUc��-L��N��R8�=ueZ����~������Z+��S���'F���7����l�C� �*�b�>ݭlY�?Օ��P_zk�����,�rf�'�![�� ?㗀��(P��p,(���O�ʻl�/�"��}�o�d�4-:��d�Ê�=��Y�~���>#��Z@x�8E��Z�{�aV�\�e_��%��c�:�?\!�h.>���zw�R��C~���|�'"3�I��[��l�����:��e@	�`כ��V3Z4�k.��e@�f�3��?�K�Yr�	�iMn��B��<I߈2� ����dU2�C%��,]+K���#�����L&�{l��iڜ�;�V?�����`��Lvf�Z��c�V�����f���ڧ��=���.viTX�}�}�]-�NYX�)%A� �z�1�u�vf��X�e���B������SOF�0G{;)?z�� {!5
���d��5��|�!F�W����+�hY��ɻ�7�[�!����_)���<�u��b�]��E��ed�Q�tBt�,<7����g���i"	q��!�N���34��L�rcv�G�w��Μ�)� ��L�{��-��$���_�<�fj�>Y4�4кX�bZ~{C=��2�	u�d�j:=�{�*85�aG���\5ka<���?�Yo]�_6�+G��u�n����Еˍ2�_5���D�_#�Y����C<�OԤb���_�[�dq�jЦS�i)�`r�+5v�z��[�Nl��LY���L	�dh�J/�O��C\UM��"��M����7�iȶ?p�M3XY;٫�������m����ǃ�d�ר�
L�4�V=)L�~�{K�`*�X*��%�PՇB+�Y����	 Ό�^ꚩ
�n�����0��W���%�D��SeX-w@�_M�����4�mԫ9}h��+�s�����&A��$ѭ�p�����|�������{¢��j���)9����>a��K���o�dKDI�X����R����DA��z3rOܪy)QIDƺZ=rB�n��)3$��؃�4��!����NŪ�ù/�V�}�F@��8QA����2�bG�h�2�HkS�m &[0�����_��.�3o�vuBv��lT��>⻞2?�:1��r�\9���!�,)k:�?���I��'���2�LRE�^�"�-_��&_X�,U2;�����B���ѸU����_�i�������5#.�������i���,fN�Q����?*�f�7U�m��ӷ�[:�;�'.F��{���[.C ^�D�>�Е�pO*Zel����F����� ��y��nP�e;J-v/���o���%|S�4�RI���]���6V�r3�/D������ܿʦ��M-�8@q��!	U�5�D��|9�>���0��ϺB��fT�uH���qNw�E�� �3#[N:����i��葁 �&I�����\ǁ���۸�}Q�V��Q@�
�8Yϝb�XA�WR�d����	Ɍh��U��5P���A�'�^R��!�ѻ�V|�(5������������;���f B�6���u��IH,�}K�����|�Q�(�K�h�	�z�:���7Tk�����y��G�6��u��f��r)D6�0�2s�R�8�^��x�����X�B�������)�N$*����A1ˠ)v�mi������Mw�}����ӭܛ~��M��&��)H\�@IG���u�^*m�nC	�S׷����-ɿ��C���-��&�h8���������sĄD�����Y��,=+��RYB����6��&��M67�lثyyV�+2�>ϓ�Pe����ߗ\K�P)f=�V8Q������r���٭��W2{�p(��^�@��Q�^C'���{B��N���V�N=82��B�
�ɦ�`M�쑫'�D$�Cw537��}���4V�|�7z�fZh5u�;[�
�s�A��%�]M�bk��q�E}��iG��0��}���
7�(N7˓���5$�f�h��C���a���;�i�0�0�����wb/�����?<K�	iB�'G��H�`]N��WߖC�������}�|� �_�k�A�@'hb�#Y+�m0K�8	=����2Y�{�&~pe�n�|�3��]����%�����l��)�^�n;�b���a�`	�J�t4�@`o�Rg{�&�s�4XR�u�/w��.��,}D�8���2��JG�-&񛵷㕾��|D)w��Ag&�`y|�<��2���a#dڂ�M�Ķ"~���}�Px������Ъ��\Jݴ됧F�" G2����𼗙��r����p��a��45?HA+R_�GmШT���&uIܴ��W�����V�-��=��>i[P_�����W��G��$�� �ʏt(��h��U�G�{0�!�?# q�:��U�.���[M5���,�z}� �q������ܐc��\���.E�#;�I��a�?��/JQU+�%ɔ�s�>�;s���yؐ�t�����9�$GBm�Ƚ��S
f��S!=���I�N6��?Uqw�H$�[zb��$o?�[8�l��f��gi����+G��<T�6��O�{�"�D��@bg��'p��أz�����m�W8���|�K���?�F���r�����1���h��P\r����SE��k�"���+qjD���1�&y[6������w�P��gAGk��#�M�w�-j��9����sf�pQԚ��Y-B ���6b�c�Κ�.���浚ᚆ,�hb[;��w���X�=$�>�|T�D�U%���~m
���ԓk�a��ӫ+�c�Sto�`ǉ�����c�2N�f%!o��/0�*���y�˄@	���m$.֓>��ns��۩/3m�9�w�u!��\'6�	-))�&�nݭ����R�r1���f0{{��P;�	��	l�P�)4����g�Fn���9{ ^ױI��Z
�6]�"�9�Q�E�'R~)RJ��S�Ve-��ͷC	J�?6Ċ'6[�b>�)b�J\�!���W�ZȌ���0�#�(��N@�^�4cV�~��b-�L.��Vi���X����J83�X�E�t�{%��cm�P'�s��>=��S�o"�k����AE����_����2�R���oko�|E3ы�jȶ�YB!t���B��4�~��A�)`���er`F��q��%� ~�9=GpƵaj�+�>�¯t�50�u
��Twe[�q�01~���~󍧁�ϙ?���ٗq�+�|�����OoH����P���ş�;\����9?�����M�ۣ��=v�՝�_��`{�-��]��t~{�s�Җ��5�L��7��Tg�����Mܶ!��Z���A�gwGz�5A�o�^��%��Oj	��v}�B�]#��6�����J��?mu�1ց��d�E�z��&�BtzO\d�I{c/�W=z�ú9R�ؓr$�7�;�ü�[W�؀g'P��/	�}�w�? yDU�6}����ش��
nN����[u��� îj�@� #�T���qZejPpD����؜zz�[��j�T�Rsg� ?�Y\4�]eA��Ze;c�8V�{�oJk�P�٤�k�W�B�|c�a�� F'_��|�����Ʌ'�"�/=�Rč�q��V�Pt���u(�N�U!��Sa�:�`����jw}��;hb�kpv�|�(�܇VN�̻����Bor���J�c>����c-I#������x&0Ž�^QyԠc�r�H9�&�{3	-+
&�|���(-�u�Jj2&Ts!Zs���[}Ѥx�|j�&�J�e"���hf�#ݡA�ځ�\J�$#���+��H����Ǣ�J�H��By���:;I����n
F~d]W1s��Ƀ�^����yʱ������E��ȾB����\)���hU�d��� �X���T�>ٵܲj�A@V	u�`�}"��8}>�~������r�8�����<��(F�w,\���9��4��*\_���3<"V$ ˩,(�X�D�^�͠$�#*�c*��v��,�z�\�3�R�Y����@���~A-A�j�,��Re0T7y�SL|�U<�k�DPjR�Xk�A����˘y�N�Bd¾@~�֋�C0�t�����4�Kcv&XuE�Y��3�Sc�y.Q:���}���W�8�f�j�[�Bl���_">r���[��,"����v���x�/
p��9K�vـA^};�y�@=���&i��Pƫ�y#��B��n��=*���1�DE�_�֩;���L�o�a:��US������d�C` a��o��f:�P�0����-��9�1�	+DZ��t�nAQ0�O��ad�'�����M�Ha�~�N���'WG@�x���?r7=	L*�2@V��V���l�g>s�L�`ڋd��m��Pjp!T�;'���H��O)�h��ia4e̼�L����-PK�qx"r�C(~o�(6�wg����ڹ���T���Z$a��yv�/�;�tw�c���)wHrW��v�Iԇ���`Vb#2�N�����Ɩ��~fZ��xW��9�e�W�!�}����d"6�T�ܾۤ�	��>7FKN����i�Oԭ�A� C^e�iC`��J6J�_3��$&�R��a_w��pM������fw]�w��'�wbM��ަ��I� ��/pA��y��W��"]d�u�3\r_+�C��n�sMM�x&5��n�����S"�b�9���\L-V��pn�����Uw�W�R�	{��>sr�&�{y-�m�wTkF����f ����kQ����˧�(�u��v(��C;�I�-&�|^�F�.�N�
���$=�y&�G�����0����nxb��mt��S�ح�&�$JP��P�cfoko9��Bث�V��r;$E�?��r�I��r�͘�\Ij�?�G��on��>�N�&`ۯMJ���z$��ݻ����Z \G�q>[T�ĵUp�C%O���n�?�����,6��� #F��W|�[���Y�/�!�u9G2*`�N�R�`���m��/~ӲB^�;+�q����:z���J:� ��9�����,$5N5�l�J����fJo=���D��#`k�.�|��U�*��W���tdа¢���c����pf�u��R'����n�+ǝ�tj�ʠ���>�Mr��1�>���u�S7���9o.��dQu.*�sq����T�������C���*4�ǘ���L�%�j���Z��ޤ�T"�	���U*�^b�[���gP�Y��R��[�#,����|%>Z�G�[b�º�{�X�yt���ӯpfz����7�[=<���-�J'�I|O�a?����&��&S�0f��"��`���e�GNr��3K=�.��i����#7|;�x�M%�o�������ܐF���[�-m��sS�1��1�,a7h#�CJh_��3�EB��>�J�P�ˊ�g�\F�+F,��_с�.�P�zظ��?�,yy�Y�c�/��������Z�٣S��ձ��D�F�d��8���+SʌG0(�f�l`�l��$�Jz�����oK���s����#&����u�Hd�' �ɼ�T�Q�<�޹��ʹ� v��<�Į�vw���c(�:ؗ1��G��H��ܭ��R!e�L+�0�� ���&aw^�ˑ���Tɺ��`�ba�����~NW��p;�}�l�0Ծ"�
�H?t����
���L���A:�d�8�5�K+B��FZ΢v�d��Z?f��%�9>)~��������L���e�
|�����<.$�z�|_��.�x=��s��93�%��T�.���#b��
ZniK5�0S#�Of�Y�;�|�a��LLZ��P>�+qF�k�ƃ�[�"��m�]�ˏ���zV=�ኒt��nH�b&�i���[0(ҡ�Z$3I�97���M$��)���̫˪�,�& �����?�%�pE�Xl�v�-ϙr��"��|=;�!{�k���5���'��������[Vp��KB�]�8	�!/�͖wT�)����C���a}��l���?5������= ��ɬ�5��ɛ#�Ϥ�}��@N�!P�g�*��o̔fF������g�>��"%^Ӯ���<�&�S����y���CoY/|����-�0a���v�M�ؚƤ��k����K�1 8��w���ՋT�@C��2���6��0>v���Ot�����^ۡ��A]�<���0#�P�l�{�:;����.��˱|���o�t��^�1��l3���ٕɱ/�=��@pquǨb]��R}>8y�������n��iK APsjC�t�'��''!�4��iM5Q��0� ��ON<8�<
Y��u�;w�G�4��&Nx#��G�1v��z���o�zf��+�,ǉʛ�~1��ݖ[�U�H���P'l=v����7���*.$\o_�T���G�n�J2.�~$]*|���_=�؇^����Y��U�d&���(gZ1E8��w�@�x|Lec)�K?�?�I�k�_'&|��̕�/��W���q̫�\�����`%šJ�_�- ��]��a|yWy��%�!:!�5%Ĭ3���e�AU�#$±���V��!m�Fs���18D7������>��5��N�Ε�	V޺Xۢ�/T�S��^l$)��d�SP�E���D`����f:Z1��P��\5�PZ�m:腯ևl�J#^���/�k���{Ӂ�AT.�YD*cJz���9)=b�%E;U�R�F������<Wx+��� nd(�U�8�c����Z�o^itػ��H8|珃<�! �a�f�3R��K|I��}{�.k ��n&��Hp����j�h�-�0���)A��N�]�R��#@�w+u������0B<Jr�!1��������O$��h��1�F7�lM�1ջ�=�3㣚c�BΊ*��8i�:Ѷ��&Gf>�p%�ӱ��;���%>�sK���XL�h����Z#]����"τ�7�a�4#"�)"����]V!M�1эh� ~֫ꗗ`:h>^�Eqg��[n�!>�`�ʧ��Տ�,�� �Z%���:Pi:�.�ӭ�aӁ7�h���h��iUpvo����ѩ  �1>�� K�{�:�����v��?��<���2��f"��^�2q�|!(_Jр� �T�	&��~23R��9 �ʻd�H���{Z+�r��n\���i9��^@w��k���ՁҾ.��56�:2�D�%�蜁؄�]ڋO����2��_�G��}�98 �f3Ӹ	���h5�	 D
1���63�G�̭R�~��@�Tkp�D�=]���jn���T���0c�5
����EO�Ty��Z5q^���nl��ΧY>�������)��ċa�eP�~}�8ɂ�0��3ōJϞhr�	S�F�l�6����K(���[��P+G`D���Ur%I�<�b+�د���\YN�}"qS��R�Bs�<�\�Đ��޷�K˞t�i�)�F�iBŌT)��
~��KE�ؚ�xA���U�w.���p4�9�h�w^�p��>��? ��-?�>���`��J��B����&��4������F��y~�ӘA� ���RR琗��\��ED]�v�[6��M�����p���}��0����t{$U'�%qb�q)���6�������y��c�\?8ez�� ���k��T�F�!
�=%�f�IL�FT�[�P�Z��Ql��P�%P���x��(�ka�H<� Bxu���;�'cG��&�6�ZG�&�nt�O=~�M&��_���<t�F)i{mFھA�b��αg�2�5Z��O�	�(e�(�d�HW�~�X"��;�>xV� ]�d�~�e!��ࡶCh�ҙ��z�b��������A�stՍ����(�`𜏉B�Fb"L��?�Ć��Ayң=�i�������d�D��H6ᛠL�Të����h�jNq ������X!�l���v��D����R��}��5�9 ���I�E�93�9���-�Q�;JX��9�X�<k\�CD���s3p�g_����1�k
3n�q菍֢�jT���aDB�Cpx�gb0N��s�ا���:�M�����"�����wTW�"��'#�0�����u�_�������bz�b�+f:�B�FB�?�s�}9��v6��5q�g��U�yeaE�n�Ӥ�ѥ���Iz � �:�lM[�9>1��u-B�8���F�)kT!�!�P�G�%g��8�X���,�"̹�
�4Cg��MY��Ev7@���o5M��u<�EcKN1¹ݡ����vgPq��?zt"Y^�6�mȍxa_��yr�	���d�]pinTм���n�����*��r��'�A�A���鮖80]�I���d��5���y݂>�(�\���J���N���
�t�_(��ԧJ"�;�ۨf�¸Y�U���n%����f��H�݂�E��<b�P''��f�[y��L��أJ�ӯX�ι�*~l[*:�>��d��z�c�	<���F@q� *fz ���* `�sM��tG���	��״�����wy��W'f\f������X���C��d|����PW!-��'@-��(�]�źC"d+!\�H%f�	l>�q�RYu��m�xj����ʆ���̇���;�%������O���r��	�+�Zf��z1��B��N����9S��SH]@?{��U����q�FX����ʪ��W�X�/�����D������©� ��xY%�J�:ni��J�f���8)G+�
*I�����:-�-��Zɟ��t���L�e���98�;�}3�u����oGN�*.�r���9��U �q�G�$�h#8�	Gv�9�HxJ�UFD����#Y��ކ��*�������v!&�L7�&�(�K��m�\I��w�/��P&�ܒ'������u��R��� �~)��� � 0Ub�_����������Ϧb��ݤ�֎7(�kmxa��&GRzX(�����i�+�������@�d�:{]�G3�91�>x��%�����Y��E8]���� Ng�-J�e����W!;5Vu�qj���B)|������F1��ǰ��K�J�3����l�� =cP/ Tvn����R���0�]���G�'��m�<@A�.��qu�1�G��w$^M���8:��WՄʙ���$֡|j�q�u	�>�%.R�/U��:�P���jƭ�;"UU����!_�53!�b+����;�,��{��q1X��մ�#�Z |�	mБfһmx�,��g�j�<h1x�=��$#0FM�`i�9P��a�⻖e>�<��<��U��:��������vG��H�����W�.�8)��|�e�����\���m�H�/&�Xp��8K~�7���F��;�Dyࣼ�9ͣJ���b�3�����UY�l�.[�:�?�a����I���$" ȃ{Yܿ���ǎ�g������R��X� Я��a����B	 �0l��T�Fq k�t9ɵ�~�7�d��v�9���7S.�qPtn���̆���ʾn<���%�	�a>���D�9���9��-�.3��IA�h����uCQ�Q]7҇{\: ��/���E>���?�n�E[K�`EڐI�GY�h:2	�l���F��2sJ9� 2T�o%y�����Э�6D�6}6���f;t��{uX�~��{�(��A��1�}��%rw7(�C���q&
���7�Wn8�
��Ml_���^|����u��/b��M�U1�����δ��b��tZ��K������A �7�:e���D�����u�<Q<t�,7E�ꗹ,����	���bf|�t��V��N=3~ ���DQ���A��q��$�8L%{��;8^Ed��r
C݌lcsMl�-檿l�R�y��9�ο|p��*OQ#���LX�rHX=%T��Z�+;x�#��ʂLtއ�����V�p�9�����ߚe��xY����кhQ��^㭿�uP��0ׅ@X�^��K%�-+�;�2�u�[iUdatX+]���c�����rh����OZ��[
?��ߴW���"����L>0�Aǰ��~��8������>l�!�:r�#��]�\�X�8i�=b�����Û�M�`wh>X�����f�����ds24��ݳ��B	+q_�¹�<@<9�,����4�0�wxfe�6kGE:a��h[���B��L�K�����I�\�(%���Y � \���?��bA*�1SD�$A"<Yc�dF���(�i=��ɛ��^��]�g�~o�z�:Ү��}���KP�����>I��%%L u+�$$I�ݣR�>$Pؒ����ж�d���&M8ҙ�EN
���+S��Gc����c�`2wJ�J*#�H���/�zo)@z���k�Յ���S%�r�ǟw#�i��=JFGŔG�$��X?��Ԝ��O!�u���d��^�[F�౒3��X�E�w���^�ѷv��Ѿ�J�?�4�E���ɹ�Y���#V����,��'x=�t�{��2F�U/X�s�:��5��2�l2�B����?��x�����Գ�F�.��ω���ḡ�Ȯ��޹�ĝXc�JW�S���	��"�G>��)�PR�GȔѠG�������Ó�ⴊ{�G;(�vu�u%e�/���&%5����EtP���K�,hlu;	�S0�:�K��:���n+~C Srcޡ�)�L�Б}d��H��F����������ZA߈L`��4h18n��&l=�'�cM4��	��9�����$,쒽ʎ�>����~�x�f^����߂���g�4�Ћ����=0� �~�&G/n~���bW��@�����m�ㆄ�[�0��q�\�[�.�7�=$�y�Qd��7�س$���Y���+yD��H�f6Cw�Ò�<�_�����ʂ��Bj�{�ah%��\��!X 'w�!F�=uU���h�����yn����:�aimU5��t���d[	����w<zr��o���T4�c;ե����]�f��=I��E�N�;)�o���񯶒�o��x^`����;ʙ�y�a�ݒ`A���1k�=��H���д�06�Gþ�����_���(�\/�o�\�q+��>f�\�u���w:W�=N�Ʀ3e��F����e@��4�;C<�D��8�A�s�=��y��ڔ��A|�mj@q-~�����B�rS�������A��ϰ3�U�M:��(jt�tX�q�1eu�J�i�T^�����G��{/�f�w�OrO���m�2�	�ʵ�f�-��zX[�t$ze�b}� iA�p%��@��)
scP��U�4Ë��yb�w�;bQ*BK�Eȴ%ir��~��T���U(:a~�8c�p�Q��5��LLYbE�Wc�w�i$�vL�8�B��@��={~3��l'�1��)h�Kw�2���C.<���?�������N;s�]�X����*%�����y5k���|4P��(�OA8�JfYՕ��Ѻ���Id�	�)�����7/y~ ��	n��f\p֭�Jl���_Yj�F.��R�ʚB���ڸ��P�I[1�i�h�N�����H�!ا�3��#T;�P*�8����X�����h%ΠZ���z�&�슒��S�\��5[����n�|?&31n)�%�����F�usR�v�d�%��7u��I'�1U1<�K(2��ȴ|�":����H+���4�o��@2>�7YcI<�IPFW�#�?����k���f(�!E��!>��>톆���\�yxv�5%Nk}�dn'���o���{A�XH�UG�w����Y 彅����T<�NdA�<�o�I�GbI�#��b�ǻ/���*���:zL���hH���/W����Yq����o\�Y�W���αz�#�m?�&	O�J^�4w^ò������SC;�2���R��D��eTH�Mv:\]��C;}B���KF�nt/���t�>�e0�Fl���ZRw�7y����Z9|'#&��n�����q��B��bT����=��R|�#O�ߥaK�9d/�Z��� tz la��1�x*>���)�+�)�F&�h���~�&C5�!l�Lb}�Z*?�e�&L�{����S����ºYN��z�(��f�)�����DZ,�O?��T����[(�̺a�&��N9`�$뾝�Z�N��� U��;u0q���瓡#z�%`��P��V*V5���1eb��N����|lE�E���]<͛�B'Y��LgZ��(g�c�[8�3�%pI,y/e<��d�p�_��w��1�w�:=0����Z���!�~���V&*{�,Rpu
��> r#��G��	�ٖ���m8\�:D+�	Τ��?fd'q����cJ�*�i���@���$N��9���4h3�_װc���\� ƚ�ό�"�?{��9��rt�/Z���C�t��"(��M��R��L��)�L�D~�c���mT�t�S�RG��}�!�r2���&����Q`��Y���l��D�kLD��8�} ����N@)+n�2����Z�q�h�H+%_e�-_�r(2�T%uYvQ���SPH�
K���O�(��y�qK�AR�}ի)=Ol�	S�?�vr�'X�fO�e�-sڮ��,��5V?	�C6n]G_����PmIՉ��-�<\!�zY�Q؇�!�ѳ_k\J��@��R8�&��=�l��;/i���.����5&B1��P�Ya�$�
�	N:�M�J��+ݶ4�a��Bu�4��i�ǘ�_O�#��n�fr޹�P[o��\1;��f�&R�: �F:Gv)7��~��O<�ȹO�tg�0�r�);MPɳ�8�2uJ�:f�25T���J���^�V�))���H}�_��\�YJJ�}��#R��=EX�a�P��W���
�xX�[�O.$������#&�x�S�q}����x@P�@�^�4ӈE���`qjC��јѬ��
\I3g�A��Zu~��}�/  �`��@Hl�1x�0S��: �"|g'Ri����u���Ҹ��,�)
텛��W�dF�ѐi�����^��i!d���=&U���Οl e�(�����_"����^�r��^鉂�����k��,����]����!<��;}J�v}�X|y	Zy���?����?]�b��)���@v�&\����2:t�o3��k��!�ݠ��a��E�	��i.��p���$���@o����Ӏ]�)���kU���/xY}�*@����u��C��n�'C��?{�,o������ԍ��L�{��z�:�wVdGQp'8��"�ޅ��؇�Lm X45u����D[��������C�E$E�(B�g7�χB��;� �6�F��oO� j�[�ϊ�e�Rv� �J�8��I43�yw/�L[��TϾ.����N��P�`�����ҫ-c�3{��9�y�44��w'g��yi�猟�/�3��?)��D2���4���]��3(H����TǗ�[�\�4x؆��$z��;�tu�	�I*�hI&ph�C�7�-�n��fT+��a�6F�oin(��ӭ#���s�;e���ȸ<���r[ 2Ԁ� �����g�2����K����L�����!2$�u�+�f؉�0�&�.oRE\'��TN��o	��{�yimx�]�����^��w����^%uNt�O`x�u�"f�ʳw�Ju���y.X3������*�*�:nl�˞E"��ų+,JQ���@ϑ�t��IQd�,-��/�r¸P�է*��DL^�^���|�Nt�vsilKZ'��f=l�3�qWh��q�Jԕ��?䉑G��gY�j��g��E}��s/�1���<�%ަqL�^���l�M�!�����Q��kߡ�1��^�j_e��BW�*3��Z��V�pU�J�R�qx"It�Q�Z��4^���)ޡ��?��)t����e���PU�F���' �������u�/�L+D������i�q.��]Sc]6 ��&���	v*��+��L�SH̜�8�?��h����f�IV(��K�����˷w�?�Z�щ��\��ǘDG�Tə��r�N��͢���-���өt�$���C{ol_ʤ1X�g��AgY�Rzl5i`7Ad�*���V�L*V(����Чb+����'+�W�}J@�q\&8�r���:`z���\���ӓ�i�fU���B�DEƴ�u��gl�L��)���������A+4��ͷ)g� |mc�Dj1���G+1����2g�R����h't )&�#�B�9�<����x������0�5��cd>�%�ξn5B�_��c���9�~{_9���P�¿�8�����'�d�ۿ��Oۖj ����_�^���}�H� P�2w��O���]���@2��s:Cҋ\�Q�5v?���[�
�ivH��o�aE��u�xC_!g���yx�M�(!��
�釣���A� �G�A���_�St��%��VDeR��W+��Jȟ?��Yj�W��<��G��)���Bw���u�/#i��� *�cLCX��P�fv��N�e�&T�b{Ǐ\���52�l��38���`�����=�24ј�Jx�� �����d��W�R�����RR�|��/�&�z�]�A��($2<����a�t�G{9�YN]���o��[���
�'`��m[���?/��Y��h��⊜C�p4�y��	��f�BZ7/�vE,M����_�~(M�B�%= .�)�����-Z��`T����3�=ˆT�_�#4L��ƅt�A��+'��F����E����;鋛
5c? A�k�����u�k��Wײ|��F��~��F��=�8l�m�]��Z�]����9S�n�w�Sx#�8%���Ps0�̆F��_ʣZ/2r��f����@����N�i�l�U��5?����[���ﯥʐ��aNVG������*3Ȼ몆��!�j먩|"���*�l�Ձ<���[�4�Wt��[��Q�q�\PG44��v���P
�+�R̨X|��Jɪ9���z�j0��1ga�kXzo��n�ivF#��l�ʀjh��Rz�@�jw���~T�0�ճ5���ߴ�ڿy�?��fr�$V���ǅ��q%�څi݈�jZ���)��A��)f�AD)z���+���cZ}O�خNnS�d8���4�bb��f�1OyT
a��l��j����_������݋;Ԟ�%g9�F�KtaғP�]y�7\l�{K�u��>*o��!�{B�r��f
�x��4W������� e�M(�d�$낃�-"�� �ዼq0�=V؝�Ѹ�S�Pw<���0�c{V������(�fltw��s ��Z��Y�"����_��U�p���4�AX��W &\������l�3Α2h���j���\�.���i7�P������ge|��1@�0�r�M!���+K#0A%��3��ϲ儡��w=p#���ۻ�ڶ�UR�
��E�����A�N��������и)Z'���y�{�@�C^K!1�i�Zg '�]�U2Ƃ�|�KM�V/���.����۶��nRV�($��\�����+K�K��J���E����<���y�y ;��@���N	��bCS>B�H�kW*�>�E�!@RD[M��F�E�m����>]_�]���QB&�L�EK��{����sm��cCL�Dĵ�d�CJ�na��6Ly:؟%d^r�9��.#r.�]Қp`��k��c�ޛ�#P�X2QYh�n�,�K%��#�C%5`O~FV&���Y�JiGh'8��'ޜ�ȏ�O�- A��4R�m.����S8����В�)���<ۭE� ��V�c�-��W��.B|��`@�jr�nq�+�DY�Q��%|O�)��,wB,{��*Xx�>�M��!KH��ـz-[S�i�	��������6V��!"���Vx�EI/ǀ�H&���n�6Z����\�Ӷ�fP�7������Ӊ�#+��s{��׭]ڰj�0��*=\�H=I!����;=YH	�}�Y*l}y��y��I!�[�ʝ�U=���q�󋣰�$��ǂ*��(�3D
φ��-����1Kp"�G����_/M�0.�W	{}��q��c�a�Ҡ�e����"
܏�����\� Q�ܰX �.<ǋ,T:[�,�&O�Bj9u�_h�ǡ�6&A�	�I�k�
?��&���E�>L_�>q%"l�:�@i�)�n����0u4!�'T�;D�S��K�u��q���o�V/���>����/�$U؁%g9�{@��r��������v�M�����\V�0� �||>�6}9$�}�ļ̮�BՈB�㼚���@���X���Wf謩�H��A���)��X�k��V����lӡ�l�&H%b���9�=q�?蟿��
 ɰ���̙PD���������t��9׉�������!'�(/��,G���R���E�����q ���/�G@5TT�#�DCҶ�x0�`��[�]�#/ø�~&FSԚ7�o@� P-�VDX�S*�T�
q��^��>2,os����W,�;����/�r&��� Z��ol/F.�!/G*�J�\�n�>�5�PC�%��3����qQ��N��o�	����N�x�������M|t/����w�����F�y�O]�wW��ѽ|�I	�Bb��2��еn�3���y�f_�|S�=S��/Z["����4�A-Cgaޤ�;Y
W�/����F��~M�~W���?m�\B��2�'Nn�v3��_mOJ7�p��������������p�Psh��mR���u���p�����"�s�+���.M��ш5�B�&�2�Ҷ�݈Es^ܡ;��n���&�)� ���{v�I��E=�CΎ�i7��0�F���&'/�Ҍ���t�J*�%x�ͻsq�67�C.�u���4���i������a��o�j����
ł����/L@� �F$Sȶߕj
D�u�_tgҬ�:�ݵ��v�6��G��_n�����q�J�F���y�B�����i�Y�,�Q$��d�xC��d�R;)-A*"� �\rϮ��tj�:"n��gK0���%�B��v||��fɫ��8�tw�k��Ca�/���,MuUS��3� �P��7�z0o�g��P1]0W���c���z�i2̟��,�59�<��23h8aE��Q!�7TF�l���E�U��k����K�{�c_}jA�j�#��X(����]�����.��>n5��E�5Ga֓!V�׶�<@�헝������S�,�_��솊X��� X]�4�)��&Ŧ�G��E�E6p�\�-)I�zC�L[*�۰�&V�I6�p	��;�#�ݚ��W;J_����fmU�廪
yyp%}
Ҥ(������6���>I/q����NrD��(7�W�շ�F��JO�O~d�k"e��Rٰ����w]����+�	ln��Iۂ�H[��M]�O��7eX�`��S)��9����d�*�j}a�v�����0x�8��=�K���E�Xt�n~���
����Gbq�8�+=�T���(��9/՗z�
Ĳ�2�s �������ul�כ�^��ł�� ����:���9@ff���	������a&3~�$�-J����7a�`-�f��S�+�%���%pi��]�Ǜ1�i�R@�{�/o-��{H��_����>Y�p�k����$�@���6}��⹟�L�)5�w?��Ȅ�Y�%��v%�k�i��F'�+��[��(�Y�����(�~�z12�F(�� �J33"K�5Z��E*�K�'h�/����u�W�x�K�x<_X��7YD��Fe�ZNI�Ӂ̍���j�%�腓���D�����Ld�H�r8{��]��>YG�>���	�6��d��}
�\��ޅI&&D��!*{D��� �a�l
�[;S��8M�}�Ѯ(����F���&fn׎&?){�e/^,�T�M���%��u���4n�""r}C���y��+��K,I���ڇ,m��CNh��rp��S�&���v~VI�,L~�z�O���T�e��.���� R#姈�E�r^de{�ua�z����N�6웟�
� �,�C�"��C�ˉ�AF�������a��#��X_�@��
��`�}�:���7cR�:A]*֕/�p=8ގ+�X^'X��Xbc�R�ϒԢ��^�����k|׹��x$b�P�觩ߵ�4�Dl��гB�`���|!W�D����}{�XS���XJ�SxV�C�U��c���2�
�8��q�(�Y�i�#,,x��b%�S�ԝI:3t&��>ᤥ��[SA�U m/��F���>Y�d�1��p?2_p� ����^	�2�. ?V���ޓ}�ߧ���0Z�z|m�s*���}�����{Oq�����=t#lN�S*�1UÿP�J��Ci6��Ԯ=^4�>�Mh���.�BN�_t��+���W|ٟ��,�ލK�G�r�q�E���XT�8Ղ�&
�����ȭ��EҐZOڎ�9Ϥ�F�%4�������xE4H�F�5?Ri5,������Q����l�;�	����x]NS�·!k�K��/�)��ܛ�W�d1&
Rj���'2��dHo�� �7�_�S�3*#E/��[7f�?өe�C�i��.k�����
�գ ��`G�
?z�|�d�wh&oo��A���n!ęP��EP�h�n$j��q$��r��� ǀ����y��WM�N�&�
�bEJ�ґ�uJ��S��7���B����UZG��*�"�'C� %7){�\�roE�0��;�IL�'l�@iͤ/�8��d��z�s�xC	R��r&�d+�UQL�� �Uܷd���qwS�5ج`����� ր̄�f�l"�)�K�����E6\���a���g�-h��ǌ��%����Dz�[�m����u4��N�3,�i�LN�P������\.���%�1���q��= h��O�Ŧ��C�@���k��?�#��6	LվɾrV�N;�e�]�V���.�q!tLu�PP�E��_rVcO�4Zٹ���Cz�w��Ihn22�nV�e�ǋ���!��M����TWb�����a�=	�.��ɬ��Β@�DoI_7v\���F��%�J��b}S܆��Ȅ3�:V�:�/�vH�g�p��8`�LwUo��ĿE0�޵�<C�N�J"֠��������ӫ�̷����x������)�zsbo�w	s7 O9\JA��*,�yWJ83���FTг6�٣�*�uk'�>;���b�߽-\Ч�b(�o��/޷1U#���x8h%���<�.L�O� �N��{&�Z�[�����u�(	��C�W�3H>�����i�W7�~��*�W`v.8�Rl�f��#��pp�B���]igg��+R��O�гJ���86�!U�\�m���N�sE��Pw�FO��RGN|!���Y�����BJ]{�
Q�+�I���M�n��P
2�S��v�U��R.yl���(�k`5�i��\}(���4 �鲇:4��w-�������1���p:��x�l�~Β�����0��76�9Ö} ~��5�N(LCz^����g.H�ufaQ�%���8�����ֲ�w�`�kvȭP��D�mz��*nal�C��hX��i���߹�Hͮ�z��{@BJm,���p3�Y��ƕsyl��ǖ�0�:D/䓫�;�|-r��M��:�K���^�С�v#$��pӐ���� +��sIc���0Z�3&�s$���+�v.��߸]�`���>j�s����^+Ď�֨�8
#2y��_A����*�|F�ByӾ�M�����<P&1��3�Y�ūK.����g��|�Ϫ��{�n����Ʊ���}�6ٜ��n�ɽ����кa���8��z�VO]�^�Zқ�J�?Rƽ�`+����8w;4��1d�b[g��RnK��0��>�2N��7��4N�o���s���#e@W�S�.�xf�S@�����k�p*|B�
;	�s��-C���`k�%�4��d�d���2B����l�'�[����m��NJ��,js�w��'��a5E��=U4΋/�(�x�1���&�f�A�����2mCʆŲ�&~m�/�������k�S5��G	��Ja�탻Z)A�0:-`Q9�I��!��4�Y��{1� ��냍ֹ?t�Oq��6����3b@@�&ݴ�_�Br�_�6��ׄ��f�}�Ҧ�Q���k(���#	e�M�{_�]���y���b�Т8²Ke�[J�3�FLnf��;B�C�t��W`��j��u)v��߿3�Ɂ������X4q%B�! ��<w��_�Eđ'5��_L�c���D5��-�y
�X�����_=���a��w��In���O(?fo�I����0��]����>>�>F�q�h�t��ܢD�w�ED��C+�䬗�c��ZPUI`�LU��Pe�=�[z+9m[��7�^��Ӗ��]����:��&�MP<����=E5�-���ֈ���5$=����dz�������F���Ӭf"�u�}���	�����H���2�QԒ˫�։4V����8���,�),����Ű<�%�8�JK$�I����Tx[�n�7~��/5Slc���^e��2�<�k����=�4��oR�T?/E����6�������Od)=�����=k�$LX��̓E�2�z��ה���e����M%"%3���U0Zo�;W�[/�5��JlO�D�tZij���M�'*s�5�~�`L��4��=�w�	ݮ7ڼa�l"�E:���IF�;���r(hUc�zO-�F}��B X�@�<�Ɗu0Kr�d�W�?�p�W}�����)�ڱ&'a�Uf�c�.˛Sʌ�cy >�WFD��!���y�Uڕ�ȍ�܏� 2������1�����t=��$E���"�60��J��'ؤGԦ�3���"����[ ��6p�=�j?n�J��i����yG�m�;�O�E���p�lY���u�E�d`�S��Q܉�h%2��Ԏh�U�ݲ������y2=5w�)dɌ�v���,�S���:��\�v޼�|F6�˦�]�<,���/��w�qe�Ψ�\�|2	��B��]���U7�)�7�a����IHl0���S^�Y�׈K��]����0��#�Ԯ
貽��bLrβ���G��޽2��$�8�����o5a~TRG{D�iaњ�Eb�(�di��j���4�9�smF����WH��b�1K���*VO�7��o~W�@+�����-��|`G-+��3f�
}i��?��[@�GG�Lg,��vj���VU&/��|��<1}QVz�P��yt �H�b[��v��F�3���NVb�Q7�lWO37&VK�Y/��l���2���gU�EB��O����U�(~'�����#F;?�������l���	FkO��M�8��%^��u-g�R�=���Œe������"*.���O����!?.f����N7���������x:!.�w��(eQ��Ǒ�!���
ԓ�bq�r]���1�h�
��C��0�x��c��
�N~j�n�e5g1�n>�=O��G����c)�-p�aq]�cg��7�I����Kxq~^�0�	��2\0-̭�pd³s��Â�֥��"�i�D'���W��a�u�mL�k��˽��W��1[Y�>6� �|b8�g�d�:�ܞhQ�j��$������`8k.�G��jOk0���E�eR6�Mwn<��u5��1���6�9U���Ny�"`���!�I��H1���-0T��u�.�$���E�ۓ�τП��M���<�4]@T{��Y��'G{�2�|@�u�Ŭ)
e�J����}��3�n|�89�Zզ3���W���侼A�4�SE-߈�P��Ɣ[b��&�n }[�<@��yI�-����KK�˷a��:�,x�c�$�=?�̚WM����>���I��nvfh��X#T��[IFU�+*b�z�޹�@��,��=�:�����a�=o�[<;��^��ݺV�T	��P��&��-�_�Kkisu2�����#�֖���:R�����M��@)�ǿ�a�'�O�̀�r�D�.r�8g�w=r�\~j1sc�{OV����y��W��Ee��A����㺽�@z���V���-މ���ץ�Y���\�m�4��,#P�8����p��� Q��r� e��T��s�֮݅��(��x�Y}<�E�e}9ae������DH+�8��to�DX�4P�L��ꌃ���+��s�mu���A�9�FŸS?��{�xt��:�Zb]\�D�m���Z��M��T��;h׊�N�p�ꊋ��ŅJx�L�^����Zj4��.��8$�#
E[q	�0f�=3�O�=٣8�c��a1��/Ns��m���� �,IB�pQ ?8��Ĕ���I2N#3r޿�ހ+��F�~�e���b��i��՗U?� ������ɌS��F��QI��x� ���`��6�	ȝx>Ю�P������Z`�A���E(o�o�AI�)�w�R�q��/s7�"�bv����&�D[EP^��uN�����6�5��9��9��%{(��E�߫�̍b2��y~�����=f��R"~�>~|�o�R����Z��&ึ������K�]��<��d|����ݯ0����J0���Hg�f8�A�h��̨�;�����  ������@LT��QL�եVm���w�oT�t_r6�z�:d~%�^���'�yK�+R��!��J�h�� ��b������G�I���b`vY곬��qmE�NR�B��K��eE,gt��1,�T�"E=M�t:�����q����[�������$���V�Ҵ�`���x���Y�lˎ�9 ��Əw��f@�D5'�Pce�	��؉�Qn�[@m5䑼�3����1C�����n�;��3���S�l���\���ްɣ�Mq�r
o&q@��Z}s����}������)a����cwB�	��l�5I9���<p�4E}��?�������h1�y=/���hvDi���XV,B64�ye����'����E"o�z&�]���J$y�n�U� �4�aK=��8{4p5�NY��Z��fݾ��-�<�Ӈ�C6�b����P�C�D��Cv>u"TSL�*7�ڋ�٧R�'����30��r���
 KaUx yԢ�|t�����2���UV�9z�l�=�9��~�yi��j��vMDI�'�6�)/�]	���&�s�}*�v��53�����;u�f��#�r}��\m`�����։�^�e���_�'_ƶ�-�ă�ХS>���3��j3҈m�s��,�[Q�rߊu��B��Q��eZq*����c?��U�іU�����\�Z�u#��!����@*�+�^;S�/A7��bƌu�b�379i�ע*���m��8�d?�z���UiVc�doJ�>pV��g�ҍWD�4!<��^��o+����sK�{f� 0v��(�40�Q���;N�n��㽩��!��]U ��a���ٯ�MG��F����C|�P��U	��T�!%��tA�**��:���=�|jE�f�Tӝ{��l¿"�.C$n��G4�fٿ��ցjEc��7D6�P�D|vR��mH$~����un�Zs���6a ��+�˚�A���!'�No0	�m�d0��h_�E� -uf�K�_����x�/�Yo���>��Ѱ�.Ȱo�)ß�y�k
)R�~ӭ�������a+6{�o*Q!��_e~�s�_�r�]c/��t�27ڽ�9AW89EJ��5�y����Zm�O��w��㷃~hH��t1��LF���q��|�x�;=ϡ�4�B���E杳_ VQ�^��"l����	�OszQ�\��D���`m;P;���y��G�&����Sk���7[{㧙�"��pB3��Ւ�"��U�r�!K�#b�1�̞/� q�t��31P�RkDI�Û~�74BH�쨐OF-�l��\�P�vp���C�qz��Y�ˏ
���8|�\9��.8��x�eј�ᡋ����ْ���
8:R*Ł��d���l��6<�ݤ38�v�z�$p����d�h˵Q<\��?���-�X0g��6!?瓱�{32յ�U�R�1mZK1iѪ�X�a���Y�{�S,hC�H���Hlc��ę-�x�"��?Y�v���A�d�Î��^5�~���
B��
���W���f��h�R+D�.���${��h	�+d^Oжؚ.+���i����+*���aK[�o������;��Ʒ\X�=�x��H[@lw5�fn��MY�-_�(A����.Ɨ ��x��C�\(�����?g-[��@���=�4�S�̾Ŭ�v9�P����X�¬��AT��Vח;6�4+5�4�V�8y`��Rt<� }�
�^g��j�n��M%3F3+h�L�����7�Xt�5����׽uv��.7��(�(#�wz�����f�
Uۿ��,��H�XN��$`%�<B;�4���e���G��"�.:��Zy�s{�u�ȇ͵�'�ך�.��>j+� T�ZFn�O4�ޟ�=�����M���-:F �K��i�~��X���F<�j-�kib����'%9��.���m���l����}O���1�v�� ��!ݯ��C
�ΰYрxxc��r ��o?�"��k�F�J�t ��C�*v��O.tY�S�-�3��9q� �'�@���})��kgJD*�
�E�m���ʇ�4����G�-�`����G�UdVS�����։��-���W�C������c�N[���{�%���b-ũD!g�JD���ݬ��� ��L���2�����+�J@��f �ٴ�;ț/�	�Ofnd8fi�����U��a>�%l\W��6l�
k݁�rѡ� G�� +�Z8t?�@=��/�i^��"#��UNO?���\ns�/<��_�R�At(\H_A��U�ʆ'���EY!��m��ZpZ1`��:�>Qh���8,j:�~,�TR˛���N����1�>�'M ��<�{Fg[!v���9�4�#T�9��#�#������:3[���J��.�=Cj� E�>.8%.�i�-Hp�<�
M����`���	��ۭ�bl���8K.v�6�g�Pݨ3��6����.0�Kg�Zm<\�۪��Ѭ�� sB��v�ʁ������L(�I(O+v#m�3~'<P��Ya/����NN�;�����U-���l��I7+bc�'�؏>Qo�UU�,�̠��Z�QE�������h��ʈ�e�}�β` s�O��Q�]5o87���iM��p�p��D�%Gs�B�CxM��y&���)������|7eԪ:'��ohD��+�ۺk���i��8�<��<�O�Y����h�z������n�27����ӇeOx��`*o���w����i��+ebrB�	!�4Q���s�L40�ؽ����\�uz۱mx�7ʿugq�f�}����dᵨ;�m�tVr��~P]�~��jy�|ٞ�])z�L�*|�ƃ�@��>F�6K��WZsOg���^d@�Y�&��~�K��(x?6F\�;�W�D���z�s���I��#��o�c?��$���>�9�Ҁl���u_=O�"�m��a��$�<+lP�B$zY�����s�!�H����>���cʃ������^�$��'��j�z.DSg�Q�7�=)G�J@�m0�I�"緶]B>�F������z
F`\��C�zp�V@���O�nU�7���s�I��?����׸�ط�\o�F�Dy'��(�r��/��̋d���Y��I�,=ٱI�~�zn=0����2�}a9XL�+o�&����۽0�"M�nV��21|�`cD
P^�����(U�Dl����n@f�kC�
^�����l�y4����9��\Rԓ�]��-�/��[�o�鉍}79�[mcp����/��S�V)�Q�Ѓc�!L̙/ 䠁��+b7�u��.Ç�bTV|N��Dg\mʶ;�X������x��o�z��B&L���Q=a��p�q�'ܪ�~�����?է�������7M`��y�C��S4�&����;n��!w&Z�g�G.rW%=U�,���?�aPh�o��|�*Yly|��/�u����2$g]=_aP�Rf�����0� D[���j�J,�E���5#���S�@���94�q�Xl@�֘��ݿ9\�>��ʫ�8h<C7N�/-��<r�Y�4븋t���mP;�0@-s��2�]%l|���o2�Y���W_ݟ;��T=re�~2�;m�K����i|�q�I`>�w��v�Q�	��D�~� ��Q�B�4J�c<l��9��x�Ҭ ���+��f����<��gu��������ͥ��Lz��
Z "��r�.z8��)�Va�ơ3���ZƄ����}0s�	��vz�/��w��� �1�ZT��l0�7(7*!v ']Iy�Yb!�{�H�<�v�����栅�X�8+����ō��n�V�O
�ZA�(9hDr�iL��^O��m��X�hP�ذ�z�i��&��q�����Y�<����fS��J+��ұ��-���2�=�S���GN9�<�D��tR�[�b���B_��f�eWu5<eD8LQ5��ş`��W�.)���!��:G��?ۊ��`��Ƚ�G��L�8J_��4֡<��1e� N�<<x��r"��\Ʃ��[�����yN���A�ݓy�p`tg�L�qm��
�#���B�������6��NuD�[�<�\ ��4�u�h�>t
;��Z ����
�v�i�~Q\~S}��pq�S�_~��<F��%�^���Ľ��;5'��nF�tz�yym@��&���s��
�GX,p{�l ��o��׬�$�{��Z�{e�_�M~�8��O�V�f�����~6�/�پX�b�)�}tb�N����,�t[���&�W��D�=�*cB�7�xW�+_e��w��5EФ�Qb�dV�3~���y�3}{�1Q6P��>q�؆��h�{~?���z�#��9�${��F������~�J^Ԩ1�p
��Y#p�i`Y��ك���@���u��c����ڎ:Z������b��w�����1~w�����4��.���2�u�*��|D�~�oP�����|��[QN:�����ڣw�A����eT�n9?�Va}].
M��W$��f������3F�m��a���V56�����p�s�)w���=�E�X �ǚb{H�F����8��yK�y��}A8��J��ޯ|���3y������ �\dt��ڳ�.j��%C@]b��7X#!{�O��sz��^UY$+�y~ʁ{���ơi�g�q�t�8�^���Ǆ��p�>�B�jMƘ�IUM��8�L���{�hr#���U�|th{�v��B߁!��f؅l� Rx-��i��F�#��
�8�-��Y��+��)Td�0�>�lb��������R�|;��e�A�Ы��{��N�����X�n�D'��cr�Kپ�����ȕ6/=���0�V�p9�	��#��1�r:�Dh>h�|��᳗(���G�P��%� :ӯK��ʟ��*�>퍷	��n���:h �pJ\�x�ش?� ��^s�(O�5Rb���8�"/�%)��� @�p5B\DHj��}mB���^����+:[��w?t)��k�ҧ��x���~��i؎jԒr������z&.��F�V'�.���P1�����!�ax���r�r�q�!�9, ��Z���� [s��oYW�o�b�2���I��'��}m;���(������i�J�T=!	>)v��|����Ф{D#j�?������r�V@Wi�,i&g�Ü #�g_bW��F.� b�2N�{t�\�[�z��)��`I��Ĕ
�+�g�`��5�k2r�3�L�4�A�]�F�xx�B�z���DD<��mV��ݶfmp��O�����جgo��Mǋލw����Eڧd3����uk�w��w�x��G����z)��O�fJ!��v.�[��
c+�9���7
BM�_�n��^�!�vOK(�4���q�'�� m�:͖6F0����&���}ϸMm��0Nq1e�3�9س���5��?oSn�
�f�×­-�	��t���{h*�T�S,&i/��IJԭ_�����!������9�Q�������B��Ԯ?�6*G]��O��q��V$� D1�����h��!�c�̀a��P��E��?�M� o�[eV5�S����d`�B��A�����&ŖB�ؚeu��2�yw���-|t� ��#��Tɹ�Ǣ���P3VJg���wX�4��b[�w�3���R�q�CÊ�X�c:^��(ex��"o!+6e*p��W��[��lҥqM�ȀƑ�����"K�I���s(T�=�v��D��Y��*2��T|i�����}]R8=��qաؗ7�@��c:�J>�{�e.�X�Ain��2 �~H�aA���dH��xd^��>����Br�� wG�qՄ��V�,ݨ�%o�E��>^H[~ΛB�}��/]m��_X#�Y���p�[�;�����ȉ����kEW37|�Du�;R���e�a�45���wvtx���(8_��<�<V�DQ�]��l
��B�T6tbj8��e�6�@�"kӦ[���TYIub�?c��5-v�`$)�p�1�%�g���*�3nN���z{��$C	��*�q�d��N-�@�@��M�4"nP��2��[l	�ܙ�#m��㍇��e�
.�Ο����޼�7�$G�9�O��e���x��e��" �����bVӅ��f��=�	�&$��Cpe+��>ϺXPz�!Y'.�>hHs ����E9�=m&zD�+`�E���kQl�Nt-#��٨���¤�1�+��WAP����2�(sY�M�9v�Hڣ�)�� Z��	�L���6�9�м�qp���J��w�]$�"�w�-Л�ï�R�AWC*��Vg�È~ P�� i$�1�����
>T���y~����&E�HR�t DA���T�jn$��Ty���0p��즀��U�dܳ0 /P998���hOX7&��i�E�elo�^���jHO��Y1���@O��M,������N%�*%߫� V�:�lɭ���e�1�w��?���W|YI%�� ckF��L���׾A�I�\�(�\oT��N��Ѡ~"K�0Q��D���W�׆�~yr$�9���mQH����f�+��r�,Xc�Z~2j3���K��ͤIk�&N�
zX������ޗF��P��]?ن⹠��u�`cėH�����:��J�s�ͰX�Ie�!9���o,��7�#ȵAPt9��'�����=��$IrOn����������w��|�D�����\?���I%uR�D�:3�;<����p��sg���e�1���d�p�ܓD9�e�����Jx�v�aܡ ����bVN�:φ������]�$�w��J��9���u��\nՆD ��s�د��G^\D!� _�S������A�i��(��tD�`��]CȆ(Ț��?� �2H��Y5��9��b�?7Y�2�n�0*s���N����a�-R[�R�A��\�p"1,���Z�0 �4�9���O���&����:�%淏E54��}%A�J
��߄�9����&�f^�OX�%J�n3�`�t�?ω||��7�M˽�h~*��"�qD>B��-�?,���C4�+}�:(��Ge����han.Mu�S������εÉ��� ���-�CbeS4V�m��q�q�OR�NM�8qa�Y$�p�^��@e��X���
��V��y�*�r	��'��5���+�z�Z�*hY����*_ٞ�ɉ�@Ƚ?�l�Q�6zK�����zy��R����2�4���b��>t��>R�N�^ۆv_�_h:�2.vQ�Y�0Ӹ�W4=^�tǿ�>/6���Gj5Gsq:q��k���3��t��@nX��#�1�y<���!��U]��*�� �>J9Ȏ95��#��%MmI���%o[���!N��&-�RL�\r� q�|��^��p�%�ᕈ~��zϒ�
A3w�/\����-�Q_���m��Oу�l`�5O�[�Y9�.�?-0���
�F��H�g�h��6`���������a=�g�8�shAtL\�jq����;��A����� �D}��q_A��lo���Q�`�$@R�ɤy����-Hl�t�.��>{y��"�Io�/ja�$g�wjµ��C�����(i��ڡ��D�dȗ�*n���D�Ikȃ�dv�Vj�"�ܧ��vo�\7I5eo���E�H�H"%�&a��?)3r]�j�T�㽧��P�:$�Wy��ʾ"�6�F<p/'*h��wj8=E.��������1�朽����O��k��p���:j�?߆6o��I(��u���2OֳAX.:���QWC"��%��d:��&��<��/�����&�pԚ��n^�;�y������2'm��-�x���N^~ }\9��;��E?|Pr�D6����#��G��/'#��m酖8ɋ\�t�3賤���m9�`	<[�H�7�պ*R^(�h���t�I�q�����oNqG�e�7Z�4l���%x��A��N�Ϟ�7��mK6�1+��h�$&[�t$��腢� �T�j
��í�oH���d��!x����p�r�MĞeɄ�����c\杗d�2q��H�F��A*}L�*1~�X��`�����f9Y?��F\v�R�K:O|$g��DI[^?�vEmM<{�gb/� ��4�R��/ 
�K�!�t�U/o���/�� ����ĲZWg�i�M'��֙կ���N�ǈ�^�]��ȑ��[�N��9�ib��F��G�WH��7!zd7Ѐd�9,NO���i��*Ko;�b'D�	�W�]*n8��Uo��p�Oo�ω��4*!������
�,�Kj`Z義V@ ~/��� LBFk�7f2�F�a�#p�kOE#�:�5���|u8�ͬ4]������䘄'FO�'�W�{�X-�u@+�<LrH%;�A�T��\n��K������Cs!F.�JQ�U�������X�L�=���qLË��QN5RU����[�)�O*~�Ǵ9z���Tx$Ÿ5���h0�B�j!+�me���y;�jэ��BDR��D��������s�ʍ=��A����b�3R��l��,Z�Z@N���7��s���"Q*O4 �� �=����Ոy���6v7;�B�im9e�!�Z�����-��[��'���c0߂-�aA���{t|֚���wv�n�|膨�c` ��C�P��g��Ϡ���i�9s�A�Y�i�%�S���s�c5�fo ��Ů�m�xlK�}�=x�G����?��ڨ����E���t���q��ަ��-݈[ܪ��ZB����IW�YK��J,�&G"j,���=��{xILcqo�C���:�t+?��K�(��Q�i�5�Uc]���x�Y*�t�	�7z(
��KO#H���<d�ۄ���|�;���H`�
7�:���6xW��k
���B� ��>�c��ܷ=��V���8B�ns�{.'YSh|�Ȕ��;�Z!F �ҿZ }Wz���2y��V�C��G�~�R��"E� �ֿ��9���0������g��<�_�;��/6I�s�� �&��10��)�-~d@�>�����K�����|(4�-!��E�<|{9.�{�P���C�j`��pu�,�n>R�j��t���ߵB?�j�3��i�7|+儈}]�s����W�s�}q����mn�J���RLLnC��c�m�0��5@6���~��KjT&V9��e�._�LB^S�p oj�kT�j��Cr}���'�ikST��8�AgH�
��k���;���	������H� ����x�c��,��塊m����n��ϝ��oy�¤��#�C{�	�Y�#jR�]b�iJ^S�%�WN����3C!��C���T�H��M6	Z~���%4~����Չ�a?�.6��m��Bo�5|@�iT.f��[%eP�g�&pk����sf�+� x 1���������mT�N1L6�L���8u+D��Ú�z�i��yG�n�5�2�p�sUU�����%���zX�ؾ6A�
�Ȥ�\�ۈr�`f�k�m>�h��-��D�@v84)�
�,Y�d��ȗ��-���Q��O׊t+���b��$�Jq�xw�pc�^v����)�;'qr�NPS^�3���l�Q��KN �aQ
�o�cﯖ���Ҏ�˒"
��:%^�bS�*��xH�x��P� m���Tf���9s�(�>�5K���x5�vrA�s��
��pɇ{�T�n�A���-h������P��Y��BAo;��-�pk�.7-m�k��I�3���)�ܖ�K���G�I%��lN��ް�ZkQ��R$�}U������R�R΍w��I1��e�ʮN.@�S�m�E ���J��MeoHb�o��i�˙�w��ki�Ag0mXcj�7�W�So����I�L*�/�<���6L�D�_��+o۠~gn��6J�(S�+��Ws|]�NM�`LB(6��q��U��>&��-L���-2!gU�c�N�^�>Ź�g'��㇑f1uN)i��jF�����l�ڡ(��թi;:�IN�^Ż�����^���}�����M ]�E^����j�y")�}���"ƵB�rjY��6r@�ϑa�|ل�'�D�3%�AԘ�����x�P�jZ���Y�EfL)S�����ܗj���Ds+o��!�.C���;� �Z��ox*�N��ᱝuj�0?��39w1B�w����S�F䥬`z��> X�R �NIO���V;ԥo(���4�G�Bծ�F+��P��3�����C����#��h��?}v��>�k�[6i��4��ޯJ,�U�:�A:�9(E���d��H�aoe!Ί(*h�c&A��M��l�`d	��J�5��I�(+�^'Q��^5�7�o�1��<~Fׂ��/��I�-t����Lc��7
f]��
;wL�|$���40��u��a��*������=������Fz�wz'���|�c�Y�8�C�вU]\e�U7��˫d��"&@dZ׳�9�*��R/�P���"�Ձ2���KNs��m��ZY��P�/�jȫl�M���^�����LtJ��٤�p�������uTB�~6mAy�z��ek�j����v�,e�zQO�=a_6��Z��LV5�;]��z����:d4�nv�B��=�w\-w�9���ʢ�R�W��6]h��1Q�vܕ�Z�2}�a�oL�֌.<
�EF�A���}@�O���z]k�#��Zmh)a�o�=C�z�7+c�4qk����8�5Tܯ�G�<�x��	�얤���f�j��%�����`�������D�c����Ĥ+��i.VR$�W��,�{�-����h٢$N�܌M�8����ofƕBW��0\��|�����Rzg�n �6�ݩ���BCS�қy�z@o"㥠bwǲ�U�=�Yj;6��
���ʏ L�)�X7�Y���Y����^��& yHF)��"�2�8bԟ��q�9x-m�qm([+�oK9���1U���F���g+���n*��&��������S��9�}Sgt<���q4l�u��NVW���$Q�nW2^��UH�in�D��s�E��:��i?Fz��+��r����Ç�%��>�������!�C53�;�(oT7�i�j#�Y:�;�����5����:�Ȣ���H�o�fS�p�nm�Hp	�P\��,�!F/Q]���0O����;�����'�h��]J��I�|���6-���s7����=^������)��2Tchm��W�矹0���.~{����q�n�-��Օ:�c�wL������-�'�O���4��i����0b�}Cڳ�Iܕ���<[���a,n{�w����i>�4QS*�4��-��p(� �Zּ�^��;��^�`rAs&T2�p�A�nH3U��ل���}��30� ����ߔ���g�z�T�ڥ�� Wثv%7ЪKk�%�����%��G��j*�}X��b�� ����*a*�J	���&����
5�zޮ]_�e/��M�s֍����cd0@��e\"Eލe��C�yԕ�dcXu�a0�g��qE3����3��!��'چ�ރ-��� �̳����m'_�@�-����+2%�70O���/��ʬ�{遌H?�vX�4s�g,��c��{�'U����x��uyRap.#\��?�]���nN�*V`eL UK�.�0��M2tW�J	Z57v��x���i�*1�?)�ݴ����tO^@P����g��tt�X^��4(p/�|�OC>��S���}�+��T���c��}�!��玻�Ⱥ����m�y7��`+G�Ý����E�بʶV����I�:#/�<��=_��䈧DgN%���ԯ�7���|ABwWyc�n�^�n�Q%r3�邺D�V�V��i�M��	���o͞���F�A����ј/�)偽K�����bv���_�Uc������{8n��Z�4��$�]��q$�1,���ou[�g��Oy����6����p",of3�{-���Q$�͐��yU�V��� ტh�\�Ӥ�g�Pa>�~h�ëߓy�)�Ň
#�,uh��pH:��y��$$��:P�O�eLDm�g{���wyq�f�z�HPo��)u�"�e�j��
r�flm`�	OT�.��H�eM���Qށ�g�������5\ޅ	�oD�Y�aq�d�/�湴��A��+f �`�]��Pv�7X���h0�T�2�y�5�����} n���o٣rH��Bh�[��]�M�#Vё(���Ad�Ћ����˹�0}�C]ai���l~�ѓ���r&њ�2��9~r��u�v���<o�
򎵡!�y�KT��E�7ۺ�(��j�y���{A���8�u�(�/�'�8�v3��.z>�V� #N��vN>�����R�8)\}�6�ubY7�q��U���9aT|К�ʷ*+�ri� !���wL�!������٘��#u��BW�!1���b����1>=�T��a�z������y�A�� �4�A���*��F��+9 �	'��U�и��HK� y`�GQ�҂	� &w��#����Hr�O��:Dk��bN-C@��8�to����S��Ͽ~;!vQe��J��/B�����-u~G���)Cc�	�("��at?�<.����m#)��f�)J��٬�tmI�=�|~TlU�+��n[x�����*�]˘2��6d_�����ѵ��?&��9��U~H%�_�	����*����W!}g���9�9�j́�V :���(��9�7:�1�qdn���6�ak�dc�o��"�	���և��^��]Nbe}�����jt���Z�Fh���z��ru��dqc�	^I)e����6�X�=x�Nq��Ɲ�	#����-\��?xMS��_�J�8P� �:25"�.��
*��e}�%ֆoRO��G/+����R�~sl�3E��"�	�0�*�z2���l��������/]���6{T�.�w��v�t��0��b�(2@4� k�N�>��p�s~����M�=�5�h/��[}}��?4�g��>�	J������4Ex?\�m�fm�,�n��=Oo���;�j�!� JDq"��ª��?'N��>�#��H���Cv��4Pf9��z\��l��MF,�0��`��Q�'#�3m�c�d/@%c���9��CdB��V�3;|�͈N�<զX���**��[`t�<<�W�Bؘi����[��d(Z*2H��&�q���r�w���s8/|OA+W����?k��#؛��"��7�%�Ρ��P����� 7�Ft�!F��f'�iL��:|�U�\X���ȓ�`��K�3��Z�����v���<5<!��>�/�"�|(pe������F��~�r���D�����I�
����
k|���)�U��mq�:2���]�Y�n��W"'�������-zk�(�M�{H`M�A�4�тk
��:��9� MXϘ�!���,\|�d\�)����XFiZ�"���3���ٝH*�z���_/D��'�4/dM�8W�Goka`��}���`Qo`No�t�����X�X�y�H��>g5z�-JN�!���6��Y��t.y�G!�[ߵ)��_���t ��P�J:ܻ��&��@J�T���䫐G~*�j!ݘH���u9��s��f��=&����ؚnృ�#|���^4��+��'��wӞ��?��U��%*BP?�!�Ye"a�^i�?QH!ށ�awn�c��Tw�P���/�|� ]ue�rwя+ȓNF�aǐ6�aF��o�mWh��V�) C��R�"ѫ�tjnwq7�$n�O[����I7���Hp<p��$TZ�S�*͐��o+/�[�ƌK� QU��C=/�#�o��f����B�ރ���j�$�8�*W���Fy���O��ǽ����dD%�4@>a�*�n��H��pR6+�n��
 ��TӋM�d����a�Nw<A.�t8��Ps�
�%����3��.y�T��M}���ϩ@<�����G,�2q�I���	.�Ns�����g��S�~|�M}~.���ǟM��Yu%�7�4.錹+a���""mkTSu�^!��9�����ď���-��5�?���o�"�5��Jf2����P�&��Ƨ��|����H��|��s�{ͫ+3��n·���ւs-��|_�L�D�?�I�@��/=g��V�"�m��n��9�'�u�Bl{\��V�S�E�lv�6pm����`h`J)��	�ȧ�&P]Z��ۘ;��i��P�)�r�.p=�熆� %�ݡ���I��ͼO��	����u�x����@���	Ȋ���pS���a�/q�=�Q����`C�x�Y͸�Km9���Y�i���r��\:,�c`�ؕI�uϱ�%!g(�4hұ�8w�_�2�y�o�罞�ѿ}�����f�{��RN8|uN��P�/�&zC�\�8�j����n��h�����Dk���B4�Qg墜G͛=�3�9�Y=�&Ci1�����T/�V�����و�G�V�z� �siun�|�)Rֈ����Y.ǒ�r��v4��u�š�Y��<EA�E7�'�����B�Y^!�V�nG7w��J�������s��U�mԋŚf���IN�����-�o��X�#K(䢣�6����f�@�j_����=g�C'őy��^bxJD�)�v�	�����Uo�_Q�s:g����դùL�b���/_�ZɚM��z�Uʇ�:�{�ei߿�F}?�[�ǅpys��%q��sˋ2z[�v{�퇄5��oDֿ/��R���d4�9�����^n��^�ȭ^��!�V-����l�T��]�>
������d�cS�<�l��%����7`����+( �1(��5@����?i�9](�V��<mk�{O��b�>AO�{�wd�w��� H9��Q�Ǥ%�W��/����pʠT�?�,��� �|~U�G-�u��I7H��yL�	�0N{��I.��cs]�.��T��O�X�{��;�9� T����"�p_Ү���&~����\�|
ǒ�T֌�i|�����'�޾a���{�|���+4	9�AO���W��߇h��7;-�B��8���w�5<��6�J}JV� #��uJ���)�[�&����H��EZ�0�5UV�%&��O�ł��]M�͓*
��ws;N��A댬fI���q�$ ڥ<��N"=Yk�1����>���(�a��@0���D�D"�\x�e�-�_D
&>�F�/+�B2o�������� �6|%--s}�s�����a��j�mgT�p�֗ju�o�uy9�o���ya�����������3�'���;��si�\�L`W�f�������}^I�4ًvK�䅐E��kR���f�;���eLQ��:u��T�Eֶ1H�B�����	:�-��s*��hO��� �
�_\^9p
`�S�( t(��z�g�F=;g�R_l�-�̇5�p�:%��I���t��[�p��o������K����ҎBIG�+����E�Y�n���\KE�����|K:,�C�4z}�%] �`�([Iǒ%,�`�fI�q`f�O�5���Uբu�{��zn;�!_,�Sz��֗��Q�{�V*��2S�fP���@W���ؐ1m�R�V�0$�R��TW���`I��t��]B�`��~Sm��1�4t��C�� $�3.T�l�oJ۷���j0a��HBt����u`�u�(�h1������2���=��l-���R��c��}�| �8'�PBEcRT��U�ά���%��':@�
����{�qF�� ��Q��vEZmӗ��lHk�~���l����#8j
}L#��5W��#|����}��bx���#�v�z�t{_B ��7���.�����q<c�r�T�'�hF<�E���ٴ�Lp#@�hɚ�����x�79�_(����͊gE��9�i�j���B��>�F�D�H	����4���n-֗�#!^��ⓧrM���SH��t�����-���e���a�b���R}��;}<��\���TvD;0�����F{�Q�H�`�p��\����g������bh�
�����h?�λ���`t�
l�i���(1��
o�3�`^�3P����3@���3̽ہW�x|�wh�ۥ.�����\��(���)���8z��)����ٚ�v��yp���J;��3��ӽv��R����0r��wF�q#��[*j@ڶ	R+���`��2�r��Fuft	��g#:/�b��H����*(7"�+�jP�8�<�5nD��n��+%�z�tD5���\�O�}3R�G��<�K��e($0K�ȼ|wY�W�e��?�X�ڨa�O�礐�Q0��*��4U���}�^�8PC:��	( 42iv�X��W�
��`�觙��b��bI��iyPD��^M�N�+��JT���.(���|&�m�a���,*�x[�>���czFW���ݎ�A�=�3�9�G����j[��n�/L_clM=���ｺm�N��C[�kH���Q���Қ�T�9u4L����L�p�d�aN����텯�w(�NF�j5)v�J����AK�����w������/�az�2�TCC!���u����4$� �>���V�������6C�D�F�w{��exc.�PJ^�7/[�{�p$G��aJ4�ld��m�B������L�m�lf5�|�J↵�2?�m�Pit#nk4�'�Q��%O>:&��bt�yy"�׆�"ď�.�N����Y𞘰/+}�!�����%A�8�؇[�����,���u�z�I��G�>����O\���kM�P��~B�e��3k+i$��̡8���G�K�Y�O�4�Dt���\��.�ޤ]�gj���4_�\TG��s��%7�����T�`p6Z�k�=_�`^ �=����N}D3Q�?�l���	q*�F��t��])-��\��=[�#�XA+.9�"T��O�Kä[��+��z'E�v�ѥr�0��3�)�'[��|i�&�)k��`#�'���}������ϩ�o_��&Au 8X�H��Z���g�యzW� ����S�A�.�م�S�񎸞[2(�u�}�R���׾��� ����A.�m�����'�*.g�����4	*X	'omn5�;@<��3�h���J�j�>��r= �P��s+x�Z7��L"EJ���s�$*�%\��؏S�k��(�ܢ��βx�3A%G�+�����r*�ޮPǱͭ{���A��"Q ���D�{�C���WD��-k��U����D��o�D<�;��T��d�6��(�-(W�W��}!= �n*�Z�^h�{��9�#��^>q0�Bt�8弄�`�I��1��||�)a2���2�+�N�ٓ���`��j�_=
����,+���␶��t�u�).�~���k\Zn1b�Ң�\wU��?��$ �"���aRY���`�#�L�؈�q*U�Ǒ|DA͙7�Iv��� I��1F ���%Q���Ή$VH�/�lO�E�E��:a�������-�>t�/�x�[?�ޥr��cF�(�R�#Z*�)"��v���	�  ��	�V�r��Œ�*G���.\�[�[ú��#�$lW�<��uA�E҇
cogk�"�z#,Z	iR��."���e���m�����7x�0��wC�N���'C`t����$5����6<#1��G�(?E�dwqC֘F)���N\�#(mX�g�bj�Ā@�O�H��J;�wuH��'.·��R���@��g�&�'�#����0#[�`�g�5���K�����2���ˊ�����~�P� $��&8� �9�G��_��=$��_C��8�]�R=��_W��2��`@���:%��>G��(���v��+��I�E=~��>�t���W<��Ha?�W:�X��8��'"9�T�����x�bQ�h�EVt�����ׅh-Lބn�7OF��|��c\��j�!G�~������:ꨆ1��([�e�%�r(]�	�4X7����Ê��`e�� �
�~T�3�ҿ�[SzV���>_�\ ҘK�[��. ��U�}1^��d��0Ep��dzL��S2�PÉLy��?~tV2|�Ҏ1I����-�#٧`����b,#��Ѓ�>�F�dPmK�[.O�	Q!Ӟ	�?#�g��L�����O�N0�� c�N���wwլB8���Q�%�=@A Z9�ɐB��Ҥo�ڀ��ݪ��*cO1+���ckQ�eS:�E�i��Y7&L��ʏ�}���Q��}p�+�L��"$k��\���w�I�\Gm��Z���	���W�zvV3O!U~�A�*<f����)�P� E�e�����P3P3w\+z��%�0^�b����{�����3U��=���P�`@֫l��X��hs�^�P�B/�P��?��4�W�]�xh� �Ƶ�rծ��J~����l[��\���I��D�b$,kl������9E^z����֖<�b�=<��'[��3f��GӧL3^����L2��(HaFep'�^b�	� ƙ���7Z��{q�@P�-9M���^%
<hB.���\�c�H&��4�	us�܁�\t"bI��� �S���t�YIA��R�Ga1�)���O�\/��>;2�c�M#"x�ˆ����%�s*&9�uz]*p��M���4D�2FRBg6�q�nJ�Yu�	���b.��km�Ѫ{�~����9z1S�0��Tͽs>�� Չ�:�%��9(3	k��X� �6�?D�8�'}�!�49�3Ɓz�D4d2��p���#YQ1�;���N�Ծ���XVX��8�����C�>}�����}jx
�W�:Z����7*�D�٦����*���Cr.7Kh*}���\M��Xvw�rt��@���<<U�Rݦ�t�(ۏ�V�Fvm}���2��Q��ӥ�:gj �e�����Y�k A'��I��+L�4N�=^�vn��Us�!��PXso�>ˏ¿@4i0�i��綷Ĳ	OL�wȔ'�Y��bV�mNTԭ��4���#z]��q������tM������������ID,Ϲ�9�	:օ�����/S��UU/�cW�`:��x���9���9]�����D�p�ۅ�V������mV�t�?7��4n1�d����0��	�����_P%J>��sl��N+�ɬ�#������Y��܀�i[����%�D���3\�֟�;B0��*:���������r�LA�V½(��'��y������ϢV��_\N�+�Ml�" -����}X �BMy��{7���4��K����������εEo�0�S����Zv7�0v��]ua5'�4�y�Ψ?l[�]	�t�� n��_b������� ��
��M=A) �q&Ht)�� 뙡��
�]�!E� F�����`,����!zD�����<��9 �i�������3佦1!=�~����"�ĻA�ܐ1�-C��b���L�J��1 \
�/�	�_��&��)m\�[]�D�1��p�M�}��ɻy,��&���s�J�$>�X�TB�����$b�8p��T@x���o���8c���>�N�%��|T~6�as���7��0�__T��ݴ��� F}i��-�"7I��Q�q���	��N[�J�FY|$�J����O�����⻁���Oor>�cl�4��YJ����V�b�h8��XKd�O%(;fZ_�1ݒ�������e�;� �N]3��K��T:);�k!G�	�3�^���Y�7�u���2��@ٱ��/�RQ��_�.р����;ѕ�FL�E���Ğj�M>�|_Iqw�� (=_� �y�������>Z��!:!��6,�X㐛���r���'�mQ�®�k ��^�&-:�����bhV�`oU&�Ygډ��O�#�KJpr�V�Y�'�l�����c!�+�!��̗�c�k)ٓ�*ŭ8�Vx�~5��Z��u�cp�/O�}��+�I d�Ъ��3�����a��O��^*���T��������Y�`��f�IǶ�ކ���.W�zz ��@�I~8L~]Sg�(8l�!@c������Mマ0;��!�Q�[�MM��-J�̈́��*F��1�;&ؑ�χ�|�Re�ܟ�)��*��P^[����|$�&�[D9C �8� R��݇Y�5!ȟ7��u���S���]�Wp�܄��TF=ʰ�4JƦ+�Fa؇׽�@T��AŁ�8�D��n(`�~��H�/�^��G!6;0��=Գ�������ji*�ӣ%>�����`��hn��]8y�*I"�T��EL#�]� ���B��3��6u��ɥ�*Г;9�r�={H=$>���4�N�]��V� &ϲ"�%ߜp������Z��Jؕ	s�ۤ�k�N=���LUV>{�� ����{;½;��j�A�Y��8����um�޾ �vT3�A𓚄�WB�j�I�Ӛ��t���}F��2O[����!���)��*E_��ǫo,v(K�	�af8�3�`A��wGZ���uy����ܚ�Mc6oG�I1ut�4f�;m$Q-��V�hx���y�";��׸o{{���� ���� [wX;&�b��f=R'͈O�A�\��I�f(Ov ���v�VX/i%u��C�*��y��TcZ��2��_B�W�z^㝛��.Y�� �J�17�[��=�Qlx�g:���C̩<������Y!��>>P�?������Wn�d$����.ա�=�=Gm$>�x�3c�z.�:���]9p�~�z{��E��^L{{dW���2���KM�f'`�k�- ��^"��:�8pb��n�".�G��\=���Lq��hh�~ˋ������Zyi�7��C��.��_��Џ�Z��z yBؾ �6]	� �VLl��P�;Bބ�� yY?K���˕:U�+��,�U��b
�z�o�E�s�6��lh�uRt�ǥ�ˍ��F�j��f���$۳��k��ݽ�cM�V/�g���-N�Rw]��9��ߝ^T;��s���VAu��C�-�Lv�AB���4��a�*>�P��{������3�H���w3�։��'��2�(T�{�$�5�XO��s����s����Fޤ�`&�])���)cgj޴Es�u�`Bӡ4�
�[����p��pK�|���\�"�q9�e`��{��P��R��}�0@�|	'm� m���)Q���Z$��R�r6�K�$؄23�U�û`�B[d~����ӿk܏x��#��I��.��o2]=��E��>W�ؚ��0�a��F���{�h�'ؕ�����?jn˷Z����k��ѩz����	�������n�裺n�^��p�Fg�ϤQ���)�B�1�*�x�L�V�Z�N���S�ܩ�':nm  �~�r�$�+rKu3ՍM�әj���i��؜�<	��%O��)�K?{��U�tpуmS�ic���7- �Ƨh��7��!Q�5��(�;z�o`³;�&"�.�NY-��ʂ^�>"9K��О�gKR�<`ǚ����3+4��G��	�~�v�|"��)���וb���MI�j�[0���NG(�L��\@2�'���&ȗ�v8���z&rAٗ@���PY��9��ۂY�QE�O���8�`���?5PR�#��,��]\�xia�'j�g�D�ԃ5�>�0I�zť��惨(��d�I{E��CC����OܡS0�e�5;��O*w>�����[l(��僌��˴-�ٗq�ɽ]��GA�E0�s�	�FNGb�[�#�?��dp��mŪ&���?ch���을��z�;����|/jN("�&���S -ժ� �5���G'��n��G�cRF�2���-� �@/�@�F+>$���9+�������5�$N	㙷NDVy��	��5G�1y����yy�?6��,{��*��\=��Q��WH���L�dn��S��f�IՉ�$��co`$��{�Ġ�G��&^��V������*.��8���P�@I���%@c�MB\�w����&���b\�M�a !Ԇ�C�����1�ZWϨ"SX`��R�J���:}��|�
��{�㲅���ҝK@t��P�r�Hk�N�^9����3	��@�5�K�[*��v���5���y&I b޻t����;+�L���2��K�J��]z�L'h��V�-)Ɩe���E^\]n����4�Tl�T�'��,�CКf�:��w*T*�W���;���?��(�m"�TU:� �u����Fj�Pvx��x�Δ�i���(����=5���k5��]����ڊ�r�w<���x9ץ���ЦD��opQ�S����X��	5S!/��� 3��$TQ�F=����������E��9��mV9�c��|/k�Uۊn�7�B�rɳhk��ˎ�:I��1�P�!r(�M�f��r��̜0S5�l����iR��C&��Ksl
�S�/wyҘI�����LD6t�d)#���tB��n>A�-5a�Õ����������_+��)~���7s�-�'C����b(�FI)�� ���ëJ�E�S��ލ�u��%6�l��)F�9�U��ОyF��(�\;Kz'�NC*}}�w���q�<��O����}YӃ�@�a��D�Q�T_0D����<	W�.'��{(�t���F&�L�Tε���Sl�� �y���ԝ
[��y�������(Mvy�}�'���_te$��tI>P6*�`
$0&V�WlA�v��I� ަ�+�9{��SG�}4��"�h��=<v@`�᲻E���:�=�Q��C S3��InV�^6�-�<>�j��%i�n���[�ڿF0�"ͅ��-�I�4�}����@iR)(K|��[�W�E�$ԗ쾀��l�y��_Y�E?xz�H����pjU�@�x����R �W.x��M��!�������ئ�L?�c�W�hK(��#���loi�����C�"�΁V��p��Ù��G�<�O�~*E��陕*��tO2�5�FKg�c#;�6���tc�h3x�_�3��۠�	��)|-9A7��9-�wz|�<�j~%�����ƨV���Ӟ��Z��<�6hx��&���:я��7��jx��Fk[)�tu9�jK�38�s�lz>�h�y���N]	� '1`k��RIF�/�������΍��PO���T=���R4����aW�Wy:S�
��[BFt�"]5v���>� 9���q��[��JR�,sФ(w�V7�Ö7�V'�"V�3�x��P�cQ~$��=�$/��������>~}|� {:Z�K����Qf�8,�vI� DG3d��1oŝR,S(c���!������<�1''F�E��=X�J���_�)Pѹʀ��a7�ʼ���ζ�f��l� W=OV��ELT�d�UߧL����PЇ�?}��)t�
��qD�1F�T�Qc�;�NڭX����q�$��A>��m f���k�s�����%�.�F�J�!.�jO�H���@?J�����&(��<k95a�1	�,�R��e-��Ӯ���p�f�?CCU	w��z�>X�� R��Q�CA)����ž��
f	��!M�\���� ���BF�i���03i�/�����|�9�38���mM�Z�,_��'I��,�$��)gL4v��~�Rf/���G㦕��;�~���6
���G�
ԗ(��Ic�xЏ�⌠�\���H�%=Pi�n�\uk�s-�L��޽�7(�'63]}NK�c3�x������=�(���������7���G^�x,/���w��nk��].�XI��u亸m�d��;��܈,�z��7i�|�œ��*fu�m�R��	��do�_Hpm0o#����&�HBv?�?��~�O\��PɅ�O��U����z����xT=��bj�������������KX�3�t��7��㱟"F<W���M~sI�����%S��P�*���@�Y��ad_��X��[�Z~��n��O����PW����0]pZ΍ՏV�5 �,	bC����I���֘"f6}��!�#��!�)�jgχ�<��BQx3	J�Jx189!�O>c�I��o�~n����z������-�L7����7�����WӠm-P�8�1�$�Jç:ɼ���-9�U N�p���n�Ja��׋fkN��u���U��Y�H|�!�G�B����t�����NK�9�jӕyH�d8"?�	{6m�9�H_�d���=C������;��1���7}KJ�2OSMT��D�r���ܰ�z*�&���7���jg�Sa�#R�e�+�ix���c���[� 	Z���Ů"�U*NF�\�=3|R�Q�����c�Л�a��d:����>�+9uRF�k�~�_��N $E�+�q='�\��y�Oh�|T�.]0��:Pۍ|Mv��K�$Ո���X� �����t�:.�?E*-9�so���jg�2g�{gU�*X��X�w�J�n?���O�&*�0�J7���]��'gY��Y�j�����I[���'�i�����>^yv��/�N#{6@���7�Z��P��;X�6Q����[��823
�p����N�H(�qc~��w�6�Q~���i�8�T��Xɍ�Qh]�}b�+����^v�j{/�C���:2�uD�$�:o�Vz�����L����g�;B-���:�ʐ�4"�K�Ho´�O8���@�4ڣ0�d��je��k��yI8�ow�ǭO���W)kn�_59��HI��m9���� �b&#C�]9����Ug[N���̒h��<�Ӱ�=�d�>j 73~��)8����ʢ�c����lImT���5�3|��YJ�M3�����v�3�T�.��L��(Zx�T1���`&��󯑪v��.��,����Sp8������}��VFp>�O�Xbmչ�U��屄h�(D/�}�^���3����_�I�r�<*{W� 7���M�9Q��p���J��[���>m��_�7a�T��vC�?�a�P'�t���hQ7!�֥��ě��׊M$.�S-ԟ�Z$ռ�:�YD�Cj^>:^�.�/�c� (��N�G
y��T�L ��溣��q&g�-r"��4Э�B��U�N�8!:r��I�xf_l��3�M��o��t�2��x�4����B�\O�;JƷ�%�5���O+�y<�`-[U��֌a�CU�cujU�U�z�Xd��:�u�e���u���Zdj��pYL�9�^U�#�f�Ć���wF	[u�Ε�/�Wf���cQ��go�4��8����h�=`�Q�
(�c!̓.�C���gM��~:,C���W�O���4�$Dq h�6���z��Nj�Xb�����}�ʰy��[%'I��v2�#��4-��MW;������_J<G%Ӳ��H�eU��:�q�J�E;d��ӤX�^\`}
>r?��T�Ӈ;��6da&!��T��ڣ��l�|�0��Apбd�r�!�M�^^�6��$L�Q�a&�Ü�/�7M��3��N�6,!C�]���CT�Cp:ͱ�N�@��,�X)��׬��d4�) �н'��\,�Uؾ��ފ��֓`��2-G"<8q߂Ò�2P �ĸNޗ�qu6ŋj���?�@'U�y��2�(8~~v�$Z�l`�s���L&����0 �g����rQV�U�o���Mΐ&���m�ק� �
�~>�q�p���BN���[C�U�ӎ)�]���8=�vh��*��
�� 2Z;(��T�����vg<�,4�vc���1H��Z!��њU���57H���t��'@D��QEG��{�B�k��e����75�Y�$�X`�дC����L�R@>�]ʯp�N���U[���˓����{��{��{��4���,��k[A�fK tO�{�~>9N/�xP��4�!��I�MzZ�Kg���#T]clʈJ��T0Qȉ`����0W������K斳�WXk��͕1�Ĳ�ϲ	p���;�4Ӑp��'�q�$��`��	漄��W}�j�B���C�aH}O����@��(=�*�#y��.�x��s�92��!�+��ǅ�e2���9��K�	7�vC�&f��R9��A���!��t��p8cFɖ>��}�:a,�@�s����5���Z��U�*��V��+����M�7���#���lv)�.t�� |�Sq��j��KrWoՠn$�0�kc��/��qe�#��7�W�U�����ʀq��+R'����:�H=��:lw�r�0��<aU	�<j�p��h^%c�
�%���=3u�/yćNfY��#sr�2F��l �) ����+�kE�ۘ�ߴ�����:\k�q��5߱ňA5Ka0j?L[I�ZKo<��o�ޏ�^ŨQ����L��e���U�/����k��b9@��4���g�"q �3�Z��J��w)�I���G9��Y������B��Șʹ�AV�}�FB0�<��<�.���>N�+Ŕ�I �nE��s�8�¶z�Pj�q3�����	�-�cAX;���?���ƅ �&,��В��{��wQy�f��y"d��y=�4���[��Ϣ��#iƦ��j�¨v������ry��iz�#7�%.�ԤҶ�;0n�)u���8~����gk�h!a��K4��m�������17�a'�ͣs�(�����k�v�t��Uv�`B�*ѣY0s�7:�,Uy�%O4L�#R�],��<��Wm��l�4e��i��ZФ������z �!��X(4���D�?D»�ܣ�C"
��?��1mh�v_�}����̚6ӌ�*h��*ٮ7�~��u
C����|��i�FI=?RJ��C"�/a�5L&�*������4m��1?���%��'������4����M�d�M�$����_Y�@&���q��-���!e�d��b����wmY���Q" q�bd�GfK����\,��	����}���S�rΫ~���	H���V����v�v�7����}�� <(yzkԅ�x?|2���o�N����j�ީ��I����M��	l�^�;�2�՛C��C��^>D�,V��\YA&F�=�ӑ5�,��cf#N��k�<W��bZ���$4�{��#ԅ=�T�V-���"[D.��~���#f�"K�����"�}A��	y���փf�3|�d���J`Xw-�ÌҺ�f�I���1��������^���q(ew����$w��<b�80q�B�q� ^�7k����+�Sv}c�����Ĩ�F'̈́Q�O->��m^��",Qku`�{�h��1GG�ǀ&8k�j�7w�.���ʤvq-�%`�`/E��MJ"�Z��>ȶ%��,v�c=q��a'�"��3����w�nnb��?7\����3ӿ�<7x�[h/mNf�1���e��g�T���&�!��I��`�#��6P���C
/Ea��T��D�����ҟ̻e�1�3X��n}�m�SK��#���j���b��\��aå������E�z'B�k���|���&T���L����_����qg%�N}`�n>��xh����z<]Ԥ� ��1�y�~Mkb������l���?�����5�7R�y�$%�����(��R�y,Y���N��ٚ���6�'\�w�0➨�h��Ϛ��x�9m��w
=)p#�An�:�Iߖr��q:zqy�p�{��n��6��;�E�gt�T�$�B�,:Zg�G!x�-jF�->�}e=�L'�r1m��vp��H��y��D0m��V��'�	xF����LINkg�aj����8a��C�|2ɿU��/��k�qV�f�y�aŸ*��,1�Tk�@
�|εby�[Xo����(��\�"�
�@��9tPO���5H9��}!���9f���B �R��C$,�!������@\?67�{uӥ2)4�e��?%�&��������5I�Qۧ���[�{XᲹ��eܛU���B�%����Y0�æ�ZRɒd�dރ�|���߭è֞=��ޕ=�1�1b�M:=/3*�D�Ĥ��1x�h΂��NU��4N�r�誖��2�w =��t��FlG�ޤ�_Յ������zz��]��T֪���*��r���nױ�L*B-�D���m4[��fT��hhA��[�
�I�F�\�EZ�Jw��>^�b��e�Ш�͉�c�K6�����B
]6b�ҁ?.���X�g���83�����Om��&YN7U_���C�C�w#������Uzκ���m��aǵ�w��R�: �3��P�+-�gMd
$!�}��YfKj�U��R�nd[ɜR懹�*�s/�q�?��v�lv�Ԅ1l1�䤯�Ï�n���}q8��y���S������ۖo�`��|��>"~���]���.��.1�}������[}ޟ:U��%������2L3���X^�k9����Xv��Ț�����V;�}n	�E����n 9�6�sb[�ߌ��q��R���H����	x�;|l��v5�S�P���� v(�������D��Φ,f��4���z��XD��ғAE I�<�˻u	㑍�`����f��ҫ�"
>�u�ʹ���o����*7��y�r�����`l�"f�-��0��|d�h	��/�!�Ff���?�	ּ��jB����\��W�uC�vT(v��´~�ₙ:���ɦQ!4>I���	���.�]�����;lGU�Ѷ6jK�V���G��[�,�lZ��K��M8���7a8�1hn���-~��.�Xx ���Q�$VUT��׷a��r�v%�����f��3���6�5��ܜ���Q�T�vk~���[è��k����`P���h}��|j�Hlp���Ye41�"��[�+㮷b`|��H�D��)�� ��LV�݆�f+F�W	8�T8��a+��?�c�9�ޯ������0�|^���H彊�#;�(էC�M���֭R�M���\��;K���8����Ֆ@t\Rr�lR�>���6�T�c/����TkJ�7���L8s5���O���Jn�6n�����M���7�-�>��k��q��{�.~H�:�͎��7=����
��!�7�E�L�p(��m��g�KH�Coz���LrP�^:٦������\�P:ڻ��E�nd�0~�k�23��<Ѻ]�wq�1�rC�����s�QS[&?@� e��Z�r������.�_i���|�U<�L�7�����9�x�ٰ$�d���WSh�����0b��w��.\9x���z9����8)S�Y�?% :�Gt�C&�w���Yピ6JR�@:�`
t9���$��p��2��3��k�&��ò3�ϫ�@�^ �C�]j�=N��>?�!yzv�Dw�r��&aJ��
�3�/�X2/8�aA�>� �(U=���J`=h��[�`�9H��xcG �(&�Vh�Ѕ��JE\��y.z�LNsE�5��R�W�dr��<�jlP����m�+�=a�I�(�k�_|��5�P�C�9H�>�N�Bw�C8��Ym������!+B������7?���U�D�T'�coI����s����vB��B`�i(��ox�"���m�Y\�����N* ȋ�Sm�Ł@V���m���VcH��)lo��u��TN*�H�qC�
i
"fG+��;��*H�#;@`�莿 ���-�X�qOkJٯ�sĥ6U���q��r�DfB�S{z ���, K�rӝ	K	�qK
��S�볚 ���h����'�{1�UT�.�s����ďBz��G>j^�����K�5�������(3�Oɦ?�'ֈ�VKzq�@4�N5���S.ԷM����4���{�)�-��0 *�*�j��39��p�m`�S7v�)yu[�\����+��6����@"�����O���bC#Ik��o�)v�I�QRC�&r��A�h�Tj�ߤ���~5���=}��$�g��|Ǭ�[.`�9��M����j����5����Ǔ�i=l�Ur�"��H��kP8���}�"����D v���8f�~=��U_��!�%�T "ǰ��3�$�h�T4g���;.-m�ǃT�s"#��?^
n1n���4��ڎ�e�"Zbs�b�Td(�?P�4���ה������a�g��e��,Fo
�󵁱:ZHO�9#��%5jV��8ާ\9}	��ߏOq���۲,DRM��[���� �?�1a�pZ��]���C��`�]��m�W/;T�
5��ɡ	��^�~�|&b�YU$�Vx���9���ΰ�\���%Lv��9�V�V�)
4�7��q�o�Ljev������/��`O�����m+�I�!��&6�|R8�/���
��h����wEW2�$�|PX�8V��k!�
Qx�nԉ���;hFT���Cc�Y�S,
�-�$�[�������P[knC���A�af5�|��,��@P[�����Ka�-s)4��>�A�T:��㧖Y�� B�/��d�Z{�3腲��CS`FOoq�@�j�����.c;e-�Id����?�*���bg�4
}��E�^�*�e�ܐ����x�xnKb2�����X�h�0z��A��w�"�ֿ�Gt% ���r��� �@��$����P���dm�h��Es���!�y�o-x��~3E�������c%L�I�D2�	�	�߉��6
��)޻>o��J8�z�cl��,��Q���1�iHT�qKWy	g<4�@���I�x�D^Ŕ�^�(5:C)]��_�^�[�{}T�}����X�f�y޶5H��-mL5he0k8Ǡ��P�O��Z�^�4�>�B-p�i#6Ha�]�=X�1�w�R��,rn~�0�(HY���/�:	a[7U�;u:43��\��)��et˹4=XNu����yQ�!��Q�h$���kgҷ��:Ht�=�3)Oj��o_���Q^u&c�ȗ�dN��,ȋ3�5y��3|[�G�/u�����>��Ɔhևڳ�C8;m�6;r��@�帓�E���׵XS��kܻq��=_/R�/��9-8�p)�Ŏ���'�o�B�Ӈ���6409�J6����k?��I�a����P�R6&�y�� ��1�y+�y��dryS���J�ؠ�޳\k��H���9��he� ennY��n��N��f�y��c�ڱ'��a�tޜ-����������۴0����%�{2?:�`��.�&Q?RN嫳��	�-c��Du�;�uz�Y����P{8n�@��ckm����	���zwҗg��ժ��{�pSH	^upso���8��C4Ci��;�`{��!H6�-� xzoX�f`U�eT��D��҉]��a��:�JR������/N�q���W���O>@�.��^v���ž�1�
�9t/�}�+��䏙FJ���M�l�U3�}%���3�|歾tX�qÖ��&�i�b�Z �~w#�>��")���Y6�uv#���U
ג.�0=��	�J�:U���l��y!���w�9��d��$9e#�,�Hu,�2�h�]�u���FnmMu��V	��Iv����6
T"���D;���&`��C��g���c�Xr]L#�'�Ȝ{>,A;���P�K��z�� S�Y]����4���8�Ĭ��������&���ܥ��T�ĝDa�����O�V�:6�ĵ̠ڨ���Vӝ��Je�v�!fS�%b>�Vu|�k2���ҽ-��D`<��\f�t��7f�}@w��k�I^�����T���$�I:�f<7�%}�T���k=�M�p��u�������K��˷�S6��h�����4Q����k%���|��0�#_WD���?>����0�>��'�?�=��fp ��_O�zV0����@R�^ิ~vh�;?#Fi����D����k�������b�ƕc�w����r��8�SѪ�JExu�UXW�95$�q�;��8
.�S�5̫vI��i�zr�l��}Vn^Iu�D-��^�r 9P7�6l������`��AM�7����U�ä�ֽ2�%z^E�wH��[iv�� n]&�]Y�zTL�yw���[Z47/�&�|���,��a7�y9cc^�OB����O-'��T,�*-tВg��G��6q�v����E��q�{��l}P�o��@�E}1C�E,e!�d�i�᮶o�4�;�A��䤺�𒰗
�Y��U�����;��]q;N���N��0C�^�d�	��ֆ��x�d�-��=׿<em���?C#|+�,��Gxm̼V"^Sn�'t��~ˑw���P�̲4F7����_��6���r$���1R���:�[2���e����cM�����0�;���N����j2��G<�K�Q��=�C�<�&'B������IkmS
8`b���Lu�Hv�IcsG��GrY����׼=�W�dɵϙ��
-��
\��0�B��4CM?��"a����3P�K۬57e�U����' ����V�N���SnL�%5�2�B����e�Hn�:��x������l�rݎ�
>V e!�D��/�,&�l{5�r��r�G�"}8YL0D���|�N[��sf6�G��>�k�����j��W ˑh������c� �>�ЊR�"	=��'�3%��K
?��7�y��>⁝X`j���&��x���d�WL��M󰩜T��lC�^�_���(@L�f���E���N����5�$��k��j�{��{M��8��Ӿ�d��c�+��԰��["�/��7.T��W��l��A��K �yFJ�7�}����\,�ۈ����M�}y��sR\���A�w3ͣ��nB�w��I���^/CT���F#&�]I�_�G�ae��r����_1l	Q�o$	��$��G=H�4��z{֙�-r���K�dc��,�ܷ}Ǔ�]:�b�w+�`>S�h1OxK��:��"�V���_���}��\H��h�ߒ���n�Vt'��^�9f��j���:w`BG
0��=��������m��[��6�>c�e�k�^_w�]>3O�C��9}�`e�*��-YG^��P�&����Qr�B��`0�O5��Ȃ�a>�Ё��W��6�r:�C&3����M��-@�"	#)��b�!�Q�Ed}λ�^9�K��S�v�H� _���0��s
�ʹM���3)��n��P��;�W�#��_<h�B�(��������l�*3'�'0��Tyc3��ۄ��o�w�����
!�ϳz���>s�p�w�[X��H�@ۂ�X2��!����~�����Z��R�,*�R<S���Y�W�{��:pX���b���Ew�atР(�E��&��P7���W,�u�U�_"�4|���F�d��"�l�S�F��,g�9��\oHJXt��0G�3q�^F.N9�ZQ��ߐ"��p2�+���uh��9�.� ��~ ~��t#3x�n<G������C~��x�I��#%:~ݒ9����l�J 4x���.��Z�E��t�o=�!���>~8�$��ށ�x����J�D�%���J��&ﲼ�嬡A|�P��W6��.�7?K��IL�����z��	�,�<Ǌ���JcC�gɓU��O��{���h%��Z'&����a���#�YQ�=k�uF��It���9>0S���E�d�g/}�!��P���z׭r�'U�*jZ���"H���2������t�w�'0~ ����?�H��I��牗C�l!a������F�_ z���'d�d�����|zJ[{�qv������.D��3R�1�y�L�2�sp�ŰQጹmq�J��G����+O�6>��秥/�9��.�4�Jx��`ӫ'c:?�W�N����=y���YU�@�jS�/U��;��< ��Y�����-ٟq�.f�G�!X����[�����>��7��!��ۥ]���Q$�#i-~�� Υ���*�F䧒�I��^g�����g��?H����l�I�����-������Ԑ�tsW�_��>-�!��r����e�ް�~A5 #��3C����W/�YY�����(h��4(�T$ʾ��c�(�s>!���߈��l)ݑ�0]c+�Z k����S9�XI
��M�,��y��NU1o�NH��Jԯ�{IH26���"<d�k�iJ��/4�	@	*�9DJ�D#������:�F�ܺ����i�կ����=���،���
M��Z�~s��<�v��+˵�)d���;9CH��/�Y:R��]߯�D�������k��Z�z]��b���,��@ �q��������>�.\_YR}�*�)d�&�tB��@:�:�����_q�'U5OnM�߄qЗ�4�R�ʂ�(FS���@���i�����;�J&��������	�������0b`�-Yɼ�q���Ӓ����b��C��,f	�((��*�'�?Ȯ�7��$a���*w�;����{�#ͽ%g�Ǌ7��°~<}���邃��+%J�dL��t��V�ȸMhvRV�4�,�)q	����s���t��'�F�A�y-�C�!�U�b���4��A�M�)��/;�v?E�<�}�b���]�%����Y]se<�lt�(y?  �<�2�Τ�C�w�d��O���<�Du����F9$����EźrtS�fؕ�Զ%����|Ӻ�:���sC�i��7�̠���Ro��$����+�>,"�l�%,[f0������J/��⋚h7�k�}��:��oҸZ��:���z�Pt�#xN諶:s��u>�<G��92d2�T�iV�U��1ۮ�׹�\lS�3���3��[\z�Vkʡ�]3�N�=�O��@��=oF� bk ��O�J`c:K�
��>����}�ǉ
�R�̾�̞A+�0Gƿ��NrDQ�3%79Bo�:�W s�Z���'�pL$�u�?G0
�R���_4��R����X��Fh��C/��i-�I��a�_:kd�,�/T�� ���L$k��uP֍p7��9����-���1(5˼{�����ˮ/Č��
)��)�$مs����g��R���o#?����1^�.ֈ��y}�lv`['�tO:X�I�#ks�r�����	+f�3cE���e|����Ⰱ��{�-u�C����|S���Y[+IR�E%v�gn[9=��(cL/�'Zq��x���Nb��c�,`�q�h^ſe�M�f��xl�U�GGv?k�C��fDv��w7��E?�#���@���%��2A7wtGځ5�����n��l^]
�#�=��IM��}H@ ��J�(5.���~��&�`ȓ��v����2��(F�qR`���a��� �`Y����`�2!����&M��uV�����u�ھ�����d4��"�x��֤S���nH�X;�6{%�Pa�,xE�|����W���ࡘ�my�T7i�F�*�&֊�#A�ջ��K�Cq�D�{m���k����{�.�"�^��}hEbp���C5����������rc۷f��
m�m��:2�	\�4if�4��Wa�$����۱��Q��5���GCq&	5�x�����Ѽ�*�S>�q��i	�Xs����p�x�6w����5Wυ�m������H��C�Y� �2���E����=V�@� �/��Fܦ�t�XS>S�am��i��X���X�%��뗐�:a�MW�"��2X��-��Jz��ݡ�RډFe��:���i�q�$:h=(`�%��yfn�~�N*Bd�4D�UA��p�� ��S
���)J3F�ۏu*�4�p&��A]�E)ڛ���K��Īy7���iͱ��X*�w�6+V~�K�����Y>Ea���T:[Z�?Q� D�u��G���D��o>An��=�(v`/��b0��m����o_o��'f)�
��sc�^�;a�h���>3��	�A��)ۖ,]hI`N	x�f�Ko��hJ���[��TS����[��q�R�í�N#i!��������(��l���Y������D!���W�&b��Զ�P�I|xx5��P��s�w����uJ�ڷ��z�A��pթs��驋*� �;:CADM��M�M��9��)sIz���gxLc9�����מ�X��V��P0��S�6E�yT�!�q;���9�L��n�3��1�:��D�!�U���{3� 7ִ)���癖���hF�w��Y��M�����9�	|�Al�/+�94Rv��5뎘��tr>W9DK�K^$W�1�I�Iw[�`8�6���X�3����Q���4�ب �&��H�9�eND���%>�_�����AY�P(�lB����x҂vz�]��I��T�ñ���8X}.����t�#+܊�c	�N���wU�i�u�W��X��l(ah�lj��6Z���q�߹����=)�����+@���mp��G����1��vo׬�"e;a9�T= �<wf�xe��ǐ&t�C� K&Z[t�lY53Q<>��F�Ϡ����0<��>�2��Bs2p"~_*�(�;&��,���u�� -du��=|R`Oq�j;���J�t�3��Zn�q^b�a���h��^d���j/K��U^𜢼K�a��p�g�%$���l�Ƕ]��S���G��9�R����\���Iw)��bڸJ �A��U6��k�8����z�i�^i�9���� �4�v�iMzP���Y�[�[�@�m]�-�f�C��>���<E)�AZ�[�'G���
Ja&���mnC1�^"<hR�p�����؋��+j�s�;��z)��ZT��Ϩ�i+�>�jN�FE��Y�-r�ky� J�e�?��q��xh�a8�Mu��ʝnP[l�&�в%��C5QF�
��_@ˉ8�v(�S}�'q*�Ow��Fǐ�$?[,�2�n��1���3C�9���>��I$�'��F��N&P�����ٜ����be�g���XҰ.Y��I�_Dr!`�yI���L�/�I�?��'�E�5ܛ��k�,�Aʢ�ǡ�/�II������{Ϻ�f�����~�6�����d�ñ>�8硦����+�[K�s������_S6���x�:�¯�z�Mֿx�"�9������E�WD~n=�s���\��h�%b���1K�p#�Q1�h=��H[�hL�N\˨���� ����Q ���Ǹ(tQxn��t�T��}���}��S�����O��L��f�t��d�1H?�)%�H�0z�J��.�<m^�,Gf�H��ꯓS'�̮��� �ǐ@ș���@׳/�=��Y�>F���a��"9K"Z^��r��ƫ�_��U�utעb>��&���+��L`2��_��_(��DM���a:i��sY���eD�Y�"-Ch`���b�i@��z���$j ���R��Tx��W�i�B�	����V�$sZj<-�|>�A��l�i�f:�==
��"*MO7?L�&���Xl�����AQNP��'	���c ��������ʨA���&n{9��{(�F\q�\�e��v.�������pa�ʗ�xb$�����)���l'�5���=N�����Wo��̰8�=�LFcU��TB�F%�=�?<�"��TMJ�3)����[k@���!���kiWA$��8�'3�PX��M!r}]Y�Sn���)� ����?�xM��$�jQn��t��LR�*K��{��*����vi�A�]2�|Ot�m��9v�5aK�z@� hd�8���-~�(Ũ���U`�|!aQ���*�z���5�������璖)]��Ho�S�4��9��bE��+�I�;M��r�7�C��9	5	^�!Y\��R�^!�%�L����'����T���Z1�y�{\��R�?o��d�x23
|@���.�-�J��D�Jerv����SW�L�E5��(�T\a�% �i�����B��g9l��ǿ���v�P8:"��^�".�����Q8��kmLM��R��QO]y��>��
��5|梦�$�V$�Ԥ~�&%	%��!a�F@jNs��	��7nҿ �x�B](�Q�\���}!�3�0����F��R:��(�}��Ly9�G�>�ۨ�{�op!S�n�Cx�V�ŎcM�$gZ�����?�ӰYz@�ζ]L�W*t,q�ȕ����e�[�&�L7�X
J�.�<'^�R~ q���{��+@���o���_4�j�U�29��i�����@�������܋��·^Sr)��٥&��tc+?�&�p=N��������S���y9��x�)V+bv���I_d���9Q15;�i)�n�b+*��.���Iz������gċz��#.6!|��	C�7L���( v:*	~d圕��"���}�R�13��x�_�)��b	b.X��7+�L�V8�y�
_s�oX��(�ݧ�8�zA$o(HN׀u�+D��jɓ�1�V��ڦ�bd��n�h����R�}$��ZF�YЯ��C �M��"?/��@Q<��,�NaP�B��F� ۄ(���ps�X���h�|f���_����_�޺�ֈ���X���d�^-�mB����Xm�Ο�Q��ϴ��,����&0���k>+���\"��K���#L��������*���*�i����^A}��D��GT�T:�4ev�zQb3�p����CCw��Z(���9�P	[�0�r�ݧ������p�O�tz𠂏����Lv�x���?b���N%�.PD�[y��7h��!�ː;�wH?��%��@'�M,�8��?�/���+C֗-˶o���/ʆ��|*���%����]7��kc���ܜ��5�Ό�H���v�Y�[o����mm;��Bے��4���@%����)�Nl�~���HXi��d4&�T��Jb&$f5��ǵzє�$(��e��o󴛦���W�ك��d4�\�M��Һ8^-���$���S��!s���$�O�$��O����(�v���D�z[G�`��@� ȩ�(�@�=n����|�����H8�..�z�z�p���tDP�E�7X�ԡ:�����[x9~j\���tt�Woc��!;9B��B����P�~>pZCE��V�&!� ��<��N�����c�J)h���+�O�$�[M��d��f�ޙlH䴊Y����vu?�8"��]9��Q��g��ci��O��b������>6W���C�w��UV��_�ɰ�3��ۜ��˲/�T�ѽ��H�'K/S���~3Gn@�8�	�z.u��W�g"?�gM\�T+�K�[u˖��;�K�%����;�2r�36����(��~3���-���o����ۺz�
4Fa8�v�ٞ9.RU�Kֹ��RPO�:pD[��taI��q�Ľ�����R��<i'&)��H���Bq<����5�F�߀���ˆ����T`ŗ��LH%"5��i���.��L	�/�PdP;��5s3t�� ��G�����߻��";�dz���r0�q��H!����ߏt��3|���O兀�=�_�~���������C:�<LQ�J�����굃*�FHI��e��6��d�C�]�Rk4��w��f�y��~qm��\!��>3j߶E�H[8;˳�{}��B
T�C8_X.�b�R��'�>-08␶1��Z
����8J�mX�F=�ę�$�=:Q�&�������w���
��X������ḍC�n5����MD����4�(�i�]\B�G�T	 �|��4ЭP��o/�R��x�]*��������yuZ�ї��kc8W��v�^��E;��y�Hfv>웍�U7�;M�OP�0xS��¢è[Qa�QI3(U�B�V��\O����ƛTaC�F� ���/����!V#J.!� ��}�H䵛8��Ne��C��\�}�����-�5'R7z 
�<�L?�tBp�-�+�1������c���C<I��*pWYG�� �k�^����*uQ��������|I{Gn
�H��2u�3�-���Ҷ���ڛ��wP�[� a�w:��y<S9f�/�NG�v(P�� 7�RZ�A �MQ-ݱd��I���_BV��b>�҂q�f[�z�Iv.�0�8��?�A�Rm�����!<p�)�w�2�
!G��La�4��]`:�K����P{@��7xЇL��tK8=a^O#��"��k�{\��m����B�~��bs�z�)�:�ɸv��f7�Op����h����>G-Y6p?P�a�05m7��L�9�Nw�����$��y5��(�B�G)�#����J}	ŏ<_P�^�+$��ɿ�.x\	ז��zOjD�@�
~Sq�Ϟ�k�?k��7CX|E�>Y�V��[�ŉ��i�"���!�E#�j�)�m:�`���o󯋬Py>�w�f�'������І�;�v�_7h�a��W ]���Q�!ڔ�����<���׊]�)�#���&�hK��b�\���-������o�q`��J	�Ū���{�d���S�.���ͨvǄ�+F�'�.9��3*���D+n��B�aibp��ֵ��< .��~�*[x.�Ġ�:��o��i�j[�����ْ��sEd�3�V��S� M$%A��4�H����Y{�ڢ����=0h�}�^�`	P�w0�,&j��z�y�g��
�x;
(^E3J:A��T���}�:���$�%�F���
�/�dP�\�ǧdvi�g��
T<���ZЅ�ێ��&�J���#�@����`t��G�;�OMGo��0j�g��9�1=�-�j�_�
)h�w�x]�W�M��Z��)_!;*���/1�Y�]휪�X�'a24+wYW�]Փ�'Y�Z�)}���ĸ#X
~#�|�]�:�i!�E~��Q��H���IZ8FJ���1��(u�c��v�ݙ��Hsf�#�
���ݛ�	�lM?��&5t�><����jC�!���&��J�-#�)��*��1|�V8�`_��\��S$�|�uJC�ݽ����CLO1�rJP(`�8sC�y����{�M�Et��GI+�m�`�hk)�y��$����\������+hE�PtV�,[Xy�a|��W��@k^[V9(�l�=!�uV�Yc��HLS�O���P=��9���K�j�x/���oӌ-Σ��� ��_���;��(�z(ų`�u	��Zez�(�X~?!��ĉ�[��8�Uos$/�'V�N�:�y[�>�.?���
=��Q@(�����[OtL�yo�@�!�C����l����(	��I��)�,�UG�+�Ԁ���v%�)[�3R<��2,`7�/�ȣ��Lq��&[������V�%�ȇKK�f�?������MtY��ds�U:�)�nlw.�9�|s�M�9$��c��3\V����2�Ș&ot�r2S4|�:��Z�נ_5���@�a�5Of�xur��.x]�B�lᩌ�F����m�wG`.>�BuK˖��]@�~:
V�sY}�|UX_����F�����ZtUL����s������vZ�X�t]����>���^U0�s�u%y6��qa[𖎝��(y�[n���Ȁ���8�7v^�J9a� ç�0t���]��Uz��]H/�>�h
Ea۪R=9���r`WN/�n;��|�rҙ`��	w�b�I~�Nr�V���5D�Ҝi���g]�ܣ���!�JXi͹c#���i��[ނ���_"B���G�f��|kcK��1
���V��U��`2�f@�7(u"�	=V�<��
t"�#� ����|�Y�9�N��nuE��/�|sx�'o��Ԯ��Ϸ�����6����V�g���I1���m�}/���D�l����-�"ޛ��2�
��h���C���p��rHq}�0.������>L@%[��O�7p���ˊ/�W���i�w�Xkeu��=��1�`Lݝ�ڱ���%8�KV G['��'w���-r��h�8�6�L�^�<��7!+���"#�|�t��i�I4:�xK����c�\�S���������S3&N��U���fX�/�g,s+SZ4vs�s�U,c���$����V�|��	�3�*��kO3��)��3[���F5~Y�O!��R�C�9t0���r�S䯜�=2NP��y�pOͲt�R%y�|�*�NI�o��mҞ�UC���P聼�a�7�F9meid���W}��M7&�������2�<�J���/j���\.��:Ӂԋ��C�v�� �C���l�#p�JٴQ��\��z{����|Ut���n����?���d���li(�N�/���F�ё1�`�ܑ������ߢr��l�8� �D����_K��aﲬf��x�<��W��mJr��I���W����oW�$���6�L��/-�ġAt�3�DJy�6�"��+s)�)@�$�w��� ���˼DV}�؂`9>�oH��|S�}�S��cW����}|�!����\��L��(+Y����Z�=h� ���X�x����A8�|�C��*��"3ή'5d��^���~�z���^`,-�	�@�7O���hux��ʤ�ؖ�N����0�C���9�F�%�^?�y"�^|�s��Q��cՄ�u*�$�*7�)G&$���w_O�ĺZ�L�����y��-�G��擝��\B4ZX��S�>�:���n��5��x�����qt�6X�ͯ��
QxY���6���"�9fod�n?W�s�B99�����\�����Fs�F��N�9F�I��Ԋ�����pP���;��73X�P@�nR1Iԛj���n��C�LmHI"�f���?��c��#
ƣb�(
�B�J��{S��:�� ��>��j���9nY��r�PDt�df�����k���<�^�_�)�HS���ͺ�'^��V��|X��Ȅ��u���i�d�� �pT]��WW���^ЗS�}��J�0tӦ4�[2�Zo3�A��;�<�ͯb�����\��ʣ�f:�XTx�|-��R>Y�L��M�hgbҧh�!6��1�NWE%�K�h��E��7���)�'&��èpS3_��
�~��'F
 �R��69~��N{<����0R�{9r�G�Z'4�bC��/�
��i~ �W-Rv��p��ꬍ�>\���Н\{�L��m�Q-��R({W�	K������e��H�9@��*3/�"�<����D�wm:�'�� �߇6�,up�q��$��a�J�/"���lM휐O?��� A9k���ys���VgW��D��l�6`��W��\a��VQtV��_s�� �8�׎1_yOs�;��S@�/�����%TpS4ggUɇΡ��ϗQ�/�3�@��4�8?*?)o��su43��=� :\̝֬'��.�3P�-��G��}�H�%���Yq���U�]a�D�x�Qg���g��\7P�/e�-�1��W�\��S#}��.�g��+�	>E;*v#$����l/-��Yƞ�F?�t0�{�צ>���5��st��;�z�"���W9|̫�f80r�
�Px�z9�	�Ʀ�ݧ⊠�/���(�ʱ�J`�C�}X�^c��	�=���<^���eF2��Bkg��ņɔ��r \�ۋ���F4)$'&9�
����Д!9R���GQ����g�t�hE:gj
2#u��4�����ocM���R�!�b�|U����������	��6��?�w��mh�^�y��M!�p�V��]>
;B����A	���w^j!k,g�9�HF�S�P����+�C���c;ڔhM��[Q��4��	�[X��J�>3OA�G�T�A����dR�qh����52���f��D��Գ(�&���|�-��	�ݝ���2�[���h�h"H�ɺ#q��Z��k�V�neIK{��8e,=�&�̔[sXB���R}��f����Q!�J�my��;�S�mJ��s��x���̹mI �0�ry(�6��3d�Mmv�#��?vs�&��V��1��J����_�$�F�[�I����,n���p{�3����^���S3G3��a^�gСm��|7KDk�a�Q�����@ׂ$ΖN=�5�v_�G�<�IY����O���.Ԋ���cr��
�F��A�]9DR.vgƸ�wF��� Gm�/B\%m[
:�,�Yi�\�����`� ��$�3�FV9g�L��1������ǁ� �a�.�z�2}5��&-���m���
��ծ�>�Qm��7K�l���%�Wګ���D������k�����f�d����Ob���~�'�� �G�Fp^� �a��i%|*
��u
ܸ��$7�����B5�-�^�c<j�K��V�6y��W��~��n�F�d�2ZTz��M-]�PI/�~�q�m�j|I<�%%�����F�%ד�/4����y�9��if2�\�<;����&�la����5bMzTkU|�>(�����mh�lKѰ���RIã���,��*h�bj^}�
Ћ�v�.��f�C�J��I)=I��|��VGq������^��tp51�����`�[���y:H���e��E_"R޲�Nd&/�Q�^i�����g:~ڛ��{�X�w�U���T���S�r��q��8
������Wۭ��.��xO׮�����9�|��S�ۅ8@E��v�o�����U��-rsS�lK�ԯ[5'[F�>�����j�Q�K��$u�y�9�u��ɍ��V������j�d���i���>�����6O+����9�,�xS�d�)�l{��� �w�b�����{�ʁ�)b�k:8m�)8
��	[�I�H'��1�yf)�LA��"]�	�0��q!���1X��]"�ih_��7'�cKz�����1#��Q�N���Gk���C�}�$m���U�"lv{v=��x��3���0��T�� ;-�l:�{�(�ݝ4��z��LQLF�W"�'���{�_g}��k?���|7�S��a�=1���Io�=�Jɀ���η_-A7�π�@��e	��~���B�x�3��x�+t�jj%n:��+(Q��h\�p����Ǻ����g���4�a�G��������{;��������YbN�κ��~���e;e�{������Ϝ�ϙ�U��0�P�j�#��%��fn$����>{$���8���� ��:�ݘ���A�E>�:����,��"���OSS��*pF�l��Ok�ij�k�j�#�9���V�����(!�r��Đl�;�&��u�#��4�\Q:�,D^�o_�BHf�'?��nk��B{����^-�6�̍�@���U_���:�vg�}�����n#M�$�i�豘h�Þ1B��
~0�� gQ� n
��$��Q; s�S�Nr�<��9#~���,mF���}k��jmb��6�7kl@��ǻ�`
 ���彅�:lV�-Y
P�F�DfX��a�m�%��xgِRL��s�l�ݍ�T)'���w�0��6N6d3���B�4BJ� 
����-�p�Zt%��3V��xǖ������jsN�|�K���L��dAol�,���q��џ8B����x�C��^��`�h��$k��=Mo�Ip�,'�SH�a�<y�����v7�|RP�
<�i���L��҅,Տ�@�y(�[gr��4���mm�@��]�?���Ӏ�!pl"�$ɂ��@�W�� <�a�9�L�ѦB�n^&长C�a
\��n|rhE�y�J�m׋�B7x�%_;TU�8��M)guUYM�tJq"Ս;������'����;���3�8�5�Y�U��|���	_��e��d����^�ۤ����5$�����#��Z�����3���]SM�7�5�u����H���q	�mw��՗!��ٽ4�=P���b���mX ��o�{RM��h6v�EDkQ��9u�o����C�%`;� b�)� ��'�chDU��ٶ�g5����0�Iwy�����f�o$�Q�N�hK/m�ѦӪ~� ��������>Q6�{b="Xg��rN(r��Uu���`Q��q��ԙ(�B'BЩ2Sy�A��DS��փ8W�Л�x�`����h/"|�*:N��iK���ݸ��M�x&�R�sܕC�L��0�X�Vąh��##�'=�����xxOXoD@����/�3A�~ƃ �k=�����:�ɎA��ʅ�h�f���ƅF\���i)���_��m9)b Ξf<C:eiQ�|g ��l���%���,��Ͽ��sF�kl0��荒3p����O�a*}[���=�e�[c�aj}M x�
����7c���� vVs~D��.�?U��/��
����K�o��f�r�+@��+O�RJ�����?�]�9.),���k��+F#���G5��#�Sa-Xon�0x�>U�� >�|�;�,�Ę!�u�3n�%�[?z�f-�k�ݬ屻��C�G$�vS�F�Uj��bWҧͷ���:�7=�4X[%��&�)�����v��7�w3��a��Q'���y������f]�CC���!8��6�Ʊ�टz)ſS�^v�U��f1T�T'=�a�<����{@Y�T�=�p�M(R7#0�{��t2�U�n`��}B��j���qLpx�'��E�J{Y�k_�����)�v�������A���%���$(od1H�";!QJ�ޓ�a�`lT�פr%��b8�h��w	����[��}�N�����=�(�Ů*�|Hf^xK���2�>��C=�'��o��W���̆:����a�a�c�nwm��~�u��?d�:^2V�4���̂o(����(�aU�*�1����d�����j7(���	c��7� ����g����lGdw�����o��B��.NZ錐al��P�\����y�M=E`j���ܵ�{��W��������p�b����#����ga��ax��IpfA��:μ��!����Ib]R��E�܃����սD�x�c�S��O�����{��<gV����/�����]�a��X����XB�����h��v���M#��
H�����x�4��
���U0��WK=����I�]�k��B��n�4|��'J��L�Ƞ��/�R���`�E�����`�E�LX�.�2Ш�0?6�[-���D�i����EޙO��b���]�*�E����Y��{7�8$���bq
Z��l�Df �w�Q2	Ot�j%��l���W'�^���E�DQ�q3��eF�"y܀.ŞKu�����/K��H���q��ɔC,�d�w$��Oi�t��?�c2 ��ytS�tk{�cM����a��B�n�&:sq˒�z����?jTYb�3�/0�I�W�+�ԅ%;UHÜ$�Ž�����m��	jsA�YU:�nO�.�eF�5T+�`���y,�(+�l��*�خRq�W�}!�-��)8�Jf��ҷ���)�/� ��&� �VX��`۵���ݤ��a�R����ʉ�6A��W��߳�t8��~�c�h���}�1Fp޷�d]��&�ֻ�ɘ^����Sg�bj-(*^U��6
!"�T���]��о��$B�^��V��Վ��I���-��\4d�ކ� \.ܵ+=�J�C�DP�Gba��l�����c�pp�� hH��u�9M�ь�qC��"������{z���8=C9����,L��Ѭz4�ey&�L�>���$L��&��p�_���l� )���y�1v��i�f&�$�/�H�I�Y�,'�P.����N�0%&i+����"$�����&��7u��4g�\j�Y��]+��<}�O*0�(Om�J�}�;CyW׺�H�<�z}�([�s$r�%�4�b:��i�͡�a��$��� �uH�k-��+'c,�H�!0�A�QSH��n�J��g�ޥ�u+~��&x��Z��~��:vlُ�ehW��!���O3'���C�b5��<uo�vV<�ܚ!⧿�$W$.,V�U��rr����C�W�������8�I�U�9uN5Y���\�]T����l��n�7���ܫ�_Z�̿���XW����X��u �Q��;�����0CcF��:�u]�i���7G�n�<1G�j�d'�����g���bz�b��ς|.�6R�C�tK��'ɬ?ɓc��ȶ��`ܵ
�
f�:�.n�Ȕ�����5D���(V'��>�c6lh�˓W�� ��
��΢cԶC._Z!��d>��>
�"�t8{0��b�kXMKV���A����\���].�p��E$ �E�D��:��_�_l���ui����
��W�<m�=��=|�9��
@j�42��sh�����{ry��*��Q�;��M)]6���G���y�P�>��Gܫ���XƚP@=dM�B#p�Xn�W�n�2��O���e�'� ��4�+�n���5���-K�_�|7���W�u��C����E�Q� �u�"���Z8��#���z8.�)U��4����g`1��i���<��_V���'�͚g�tPq?-�����)5�t�j�S�Ώ� e�D2/�a��Ǆ�Kֹ*�P�yCJ��_�[�V�u;a�N,�?�}2/�FrL��^L��G�����a�
��u�Ц�n�i9-w��m�M���t�Tv�}����8,��ЯA�)gu+�_k�z�(��w�n��(}��}�c�����3�	�o~����Q@��Զ&���5?��z���[���"`sy&QzL(�(���^�ڹ��*�}~\R�͉���ʢ��ę�x٪OO��0]9g����I����[Tn�1e��)Q����~�,O^�7Q\b�f���'�6�o��N��$��j3�D5�%���%!�r�\�t�p `��]ȕ#�膓m[�ez��\��x�wn�oe�#�5(�EW- �q-�f;գ\��~��Q�TY�JB]�m#�M���<Z[\|��A�t�����*f�#�����YHI��%������Ȝ�2�	n�AT�8�>B��d�!��&�M���q�_����'،C�<6L!v@p�����\f_8v�*Y�r���	g��+�w�ʤ~�����j�<9�~��1m�:1����G��d�6��3�W$��"2�+�����{Ąm�WM.s�,���Hl$F�8�[An�C˦DY�2_3�*�KY0n�q��S6g�{C��w"���h�
����3��@�C�1�.�F=�^��v�O^r���1��c�+�����}<�E�z�y2���a޾R��iG��/���_��_����o%��ǼNY:XQ�4 h?3��|+�傼5��Tg��K�2�n�!$�7WИ,�n����ZA��0��� (>r_�,�� ��VB�=��):�u�����~�FŖ�]IqK��X��
������M[��E�$ct�<�qs7,���=7f�	���ڂ���?�-5�+�NK�lp-��l�Y�M�i?�j��Sǯ��@�%�=v�6� �JqH4�uM3�5j�r���$׊Qޓ�w�Z��a~g�/�{�ސ
Z�����S�k=Y�9+��v[<~���f�i�-=^�>����5����o��D]�1C`�� ߒ�8٧v/lu��@?o�8�ۍBumJ��ԁ�Fj�2����W_��A�3��Ņ�j)���!Mq����@�c8���.�*V�ir��Du���OU��{֑vY{nz�I��-�4ڌk���ʭ�M��F9�q;=95]���bc���"0@�E��I��93��9q��q��=�r�|~�������M~S�`w��ZТ�l݇[� �V�,4�sÞ̈́��1�l�p@fT���FyC.����CR* _�$6�3����Z���P�ψL��<s��G��q�ҝC�Z�,qj�ç�F��W7h%�R�M��a�u��g��qb�GP>����q{��>*�������MF����0�o݀��9Ľ�_��|/ew�]n�^�P�lp}ƪ���D����?�����.�+饩ĵ���߃[�@̅�D���9�|��4����_B%���}����*�,�+`��DjӺ�Ж^���|/���������k�q��PS0p�o荾~�3���T��ᦲ�T�1;�M�|/Va��r&��a�,�"�l���~�nz���X��~��ǂh�X-G��yX��%���i(����?��X�YJ�@�F<ƿL���j^�כ���l���v�CN4���?�w����,�A{ �����lc�i�� U%��3��z��G��u��_����L�hp���DC���՜�s��i��:���{>��K���^ w�ٶ�8�A���[������RǼ�y�f=��%=#v�{ذ���;;�\ڼ�2n>��@�NN�&�)�2�V;5�v�=j��#P��n�u��4q�5����4��FȁU	:��0�I���l�K�+*��ص��M�'>$
E�>��<7 �#�Ip�z) T]������X䁠u����`���,���Pa	#V�"
��1����+��zD��T���r����l�4�{	P�(�vQ�����ű���w%_R�~6#�Dg��O��Zvʰ���Åz��<'8Bc�מYI�G;�eMa-r����\�e�)7�xG3�D��/���x����'^���u�,���C�P��rǻ��e8�xo"Q�Z�
@����zѾ�X�y�'~���*���E��:�e�F�x��_�M�xsN ?� wf�k�
r �RF����؟�t ���&n��p.a�}u��p���(��*���\E���Lp
���&55�!Iw������R�@�*��Mم̥�y`�0�R�|H����oB��2�ص�����x���|Ji{��(x���}t.�b�6vX�Z#b�1��$��=C(�t��a�2G֤��J�M2��	m9@�VJ�����`�M+'"p�=9ǆ�3��U�x���^��'��Z�{d����Sd\I�����;"`|��h���1�C,����Pd��c˯��e��< �ɘŧ7����r���C=�M!yՠ���7v�~��4N	o,(�7��X��ņ
�~�̵Qjɾ��@UD�5����qv����(X�l�dw�V'N��E������Lm�'F�&O�pڌ6�+&{W:=��k�����B�IeTڥ�]lc�1,��_XҼ5�(�XC�b;��?��E.-����ǟ��F��C�t	Boӛ��MY���|�;��0��i�CBKe�����X	
�A��J��L���5������M+jkطf8*�O3[ǒ���G� �)�P0�����j����n�KsQ������nP��ﰝD�i������c�,�A�q�A�F,���af��,D��_N���=��2���/̑�jt����Tr�ɇc���!pʠ(#�W����2��p(�a\/t��������a| 5FA���oh���Gω�6��+%���<�2\��Y� u��)��AR�n������m�ݶ_�����N{��;��Y0E<�r��oRb�57�&��pWV�R�6j�/�L�(ƻ)��7�
�eZM�G� ��pk�CD���ш�"��X�%�X�*�����O����.ļV����|6���rҲ��\�N�2�s����c�2���Lp��QML^`):]À�؏毜����C��z绾VlL���x�e��Ͱ; �\Zg��'Y/pjT$��%Q��Z�A�O�/;�?5o1
{'�'@���¬y�c�۔Ϫr
�zM�JR����V���`�7��N�
2i�%AtYO%�Ќ� Q�q�ޟj�d!�s	�q����� %��/JH�ջ<�(�H�2�<g�����U��x�M�d����<��M.�z� ��6�d�7n������߰u�⏌�OG�L벓L��G���kfE���F�$�A 6�|��m�h�uj�/��[B׊?�)�,���b�iH�O_��r>W��3]�u�|ګ��	��X�m	�����0��_B�w)�}SX�sN��_�++�"��,�Zz����l�4��E*C��
;��[�G�Wo����Y_�]K�z��^I�X�ֽq��e�ǯ�l[�~�Ē��U�y���]]!At�V��}�Q�����ʟ�0P�
�ܯ ��Ӷ�����j���;� 2֦��PrW��>�@�nz��퉭��%�T�5Aej�nqn4f�an��jI�sx�m���W�4!���=���zH��ރ`P��{R�$�9sNk�G��q��g����?�@)��D:g��!2�W�|�/���[�^�h���벴��O���f5�f�������z|�zAJ�=3љ^���{9�Bzm�3�%˜�c��"��X[��Qַ���EE.�lu�H&:3,��ҡ�)j9����C8@�ͅ�~}���S7�_�����/E��{t���F(��[��wt쫮	|����Ȗ�S�gAȉ�����*�u\d��JIdT^��s!��`�92�3	_S�$��-əf7�N�@b��#F�[8-h���	��γ����@��x�&�V�C�������ٰ"|U��r�iF�T��
�
.i�$i��'��P�5%9�΅�>6�x���U�Ȭ 2��c���A�ʟ�A�X�<g��h�ٳJ�|²�s���:��#/�_�R@�_�[�$ܒ��#NtR�ph?�k���O�ܗ�����|mU=+�0��d���v��S)1�~���a�|�6�27>�d�����es�b5��+�����[ a��mg��^�(d�Cf��W�D��Nػ���M᠐���nZ�W����>�֣W�O ٓ7�j���J2Z�����kS����)i���Ұ�d�,L�S�[�v#�Ʉ�3��K��E�i=�}��@[<g	h!�����
�N��˯�&e��mܗDB�t���Y5s+�;͋��R_2��4��M����}\��c�O����C��N@�9�j+v�5Z|9�ы�(9�3T���"Bqrm���y�l�~�JHY�́�~]އ���� Q�p��G��|^�*��l���G��&��jL� ��N����k1o��[�����P���S{v�{uvb��q�:�ŠZ����,�'uC�!U��`�cٙv��i������wʗ��F�_�VL"�RՊ��V��C$XoE���s��\���;gRaS~P���VC7�ǵ���\�i�����muc�\�����ۨ��K�Is\4�D"���5��V@]Sp@2�o
0d*��LV��}�R\L[�,�P�Ë��O�|�:�H�-!C��K}
��@.��نԙ�Z�mR,S�����>����&���o��+� ��C���FR�u�:��
�R�,
c�э��[ձ=$cw�\��8uυ�Mk�!���<�2W�?����� L��o��	�Q��h}�Qex���+��+��r~B�_��~,<�ؓO!��5&0���ߣ��
��a3���9�g�**�_� j릇�'�[���y��bV�6/�C���)��.�:ǐ��]�Y� ����?�ǫ_��&�śnB��&�Q��4���*���ƬM6�K�B^�L_#��	�H��9��x*��ЯOӯ����*�	���`/-�`p��4��ΤQ�bm�9��� Th�����( 1�M9���.fE��a�G���=��cc�IC�"Y���-�<=�@�.�����)�^{�-�A����;�ʹx�0,��qn�U���3ߞ�P��1�0]�z�ѭ���3��)䛜��G����^��ڪ��*='i�2}�|�q�as�	����n�Y	��X�<���w�S�1"�?�����s��	"����9ٷ�"�]}N�����ϔ�{�E�����U-��1TBM(��m�?]�e�E�sW��w�6qi�6���p�y��6Uu*t$�&L��( �����~d��Ͼ�Jvg��쿽�FC���q�]C*'�,�E��ۺ��Wv�r㿎�����4�sDJ��G|��}0�f�s��$y5:A���=a����I~&�/����H�<zS�Uk�&p�EM��LL�������+,�q��r�[�z���������:��%���ƅ@.��ir��P��*d|���@�B:R���}��̓m�gH�o|Vh� �&q���G(y<�7R�'�IS$S�?6X44JO}F��[�c�+��J�4��ʺ�%4)	y���	pq֏3�}W2�a(=�U�?\�*�ܙ��4�W�Q"��F��<��f�$�ӘI:���q���.ɭ����W�18Ǌ?X�؍Dh�v�s���?J�����wC�K0�ѿt[
��K�`@���/��3�P�Y߫�#�|�v��:͠��r��HkA�Ϭ� ���an�Ԝ*}��1C���!u0��;k'�g?��:�l�/����'��w��4q�R}�&�ve.���t����s����Q�s4��'Exe�ZT�pO:�Vo�g,�����5rނ �]k�7����Q��[\�KHn�	�#��3��z�/7ʕI���kX��#ӹE.Ot`�G�f����[kH�
�9���HK֜�S_QT�OD\����W-C%��<��؜U3u�Hs�1���ࡥ����%�{�x���lF��YK�#�����[�=e�=\�9?�y,Me�5���Y9��s���Yw]��d(�nʳw#��hb[_�F5�6
k�_�r�y�S�;���%�~S�}k~Ǖ,��iN������V��]7�AϾRTDb��w�(�oe�Q)%�����Z�@�6g"�h���к���I ����<k{�
�3�_���g�Pho&]U���{�].���5���$�\ ��o`����t<���*4&�0��1����e�Ï;��b����oa����*1����0!f
i��p�F���~s^����s^�j�D�=��;�J�a�t�2D�ͦ��������X�<�R�F��s�uѼ8���1�zb�Y�q�F,@�����K�k�e����w{��'a'�~æ�4ඞ���JK�R��#�0���@��N1��|�:������v;n9���dq`�/!�;��� F|f�eL��&~P���.�{�>��wWc�E<&h�&ҠR,c�A�l�f����e�cL7У����u����żD4��m�켃��g�	&_������O�PN���n7h9�qC�M�-4�� w�gj_��4�F�v�﷣<��Z4�
�m�+I@�<>�F*B�.�p��K�R2+�=w��/ZQ�&�Ws���>J�g��`��LV�`r�_FG�au��J'Q����~��dAY���s��+8Y�:���]&���,;x�w�b]߇�ǒ��9���DqӈC�Eg'�u�$6�3J�"�"��a��W^[픋�$P�qG'uQ�kn�*�M#��$�ٛ
�G׃�g��o^����.I?~^pX���P�
���˾�����s�U�v<ҍ� �/�B� c�W�G��;���`�6�6ƿ(rT���N5ƽ|[�m�ƺ�	y���^���CkƋs�M���/R_Y
^�z'�\w���aG�f��]?<]�{`��iN&b��f���3щ��oY]Cu��WrGW�������$'A�΢�gp�4�Y@Q��*�I��J�K��K|�U�S�t�;�r~�\�M����y�6�	���_�{b���o �?'���	��՟	� �6�j��gUEUĆVtDm��XBCe�U��YMNѶ���i�$�%�^������k,=r�R��N�5��C��d|�AT^�/���ݾc+pa��<=��6��J-M��EB����X���N=�"�g�"����4Yu���]9��)�x�J5Z�
����e�Q�ُP<xl����Hs�Rk@���Dn�����ڝ����n~FM�y�.G��0��I�\.�aX�*Ɨ�oy3=������%Z����<=�jl6<�lJF[f�`��E��S��2��12��OO�蠕��j��Z�9��T@�����iI�#G�i�����Q;g濻�$Az���?�_UQ� -"�MS��iN�l�G�e���m'�d)�� �s5p~�6 ��[�7����#)�V�J�uY��k�����l�����'����T�i���x�g�Jy��❇�;��?�pp<gk�3�{:B��9'�t��uF�X9f0���u��A_��O;���У�\ޮ�Ǡ�p��j&S`&X��/θ�&��/j�!<����]N�Se,J���"=xiQ���o�U�J+��u�׍h�[�j,��f���7f>$�Y��i���hhl��S��v�󨿋V�(����Ɔ�LZ��8&�ގ�y(0<�D�>J<���ȹ�p��-a� s�	kĒ|��i3�8�w�J���7��g��}q+�Y�m$'�J�|R��1�Ԩ�/m���@Ѭ���u&$�Xg��D�L5 k�R�Y]]v?S�+���G��k\l���屽K=��G��ĴtM�l���o��/��~P�Z�����%�>�ߥ�
�5���y�>��u>�0@��}챐�{������d�5ses �����{�K���I)��P56�
B� P!֛yg����lDC[

<�+^���tmi�"�f�����zц�PZ$
�@�r	k��¥v~�A�,�D�R�b��l3���2����E킯9�;��*�rRj��Җ!c�UȂ������i>G]�T!��C�,��}M.#�ś
/������Ŧ�b[ª��d��1d�By��|�`]�#�x������)F
�������򾘘2m���C�툡�g�H<����ll��/K�!��7����~�����'�pn�)$�wcH�p�?����L���2 ����b�����UwQ���W��r�!2�epdzN<�F��_�̳�NY&������+�.���4��GW8�T�%��rCO��zos��y��w;ӗh7꺢K�?�/~]��t��fQc~~��q��0p����>	�A
�߆b�O���r��l:�X.����U�/�?������ȏ�g�������|����x}~?����Y����nUEu��Q���0�rKc���}5�U�@$�ƛo��.4EUPz2c�_��.Mץ�}+_T��k�A�f������[*b��*�-�gi{�dȈ��i�|�/��l6&q	�ר��8B���/�a- sץ�i"�d���y�ҕ��c�"��'I.Aj�À'
��J�Wu����ƿ
�^�l��̬fW(�M5?v�\6wLBA��t���hg�3�@VL�+N���0s3_�\d4 =h�dg��Kի��^@�t�`Zƀd�}+O��$�m���*�|���#���.kha�	Ҕx1��"^}�%�����8w�g��i=V�����8���;G��E��̌��/�= �|)|'*b��`t�,FQ���I&$5Λ���Kz������&�3+2����m������:I�)�����܇�[ۇj�VƤZm��ɗ�B�"5{RWeWu�8�|4FsvZs�G��7�}2Zd�d��ȡ�s��a���ݟ�5K�Ϻc�'n�D��Mgo@�o�m��`yw���=��	�ÀQtΜ�������:�@����4�2,X�C����f��?S7o���-f�$�1�dIX��_ɵ���9��\�_�r2֤8\)�%tB��xNxFP����i��LP�L���S w_w��G���J�,�D���Oх�H�/�l`rF���V��Em�M����ܟ[�kt�Yg�+�.�Jn_���ś�$���RC;�x�X�?*x�N�S���U�L���(�9"Y��!@h�o���ᨨ�9��y	Wt'�M��ىP/۲3X���0�I�>�I�ocv0fs�]H�����1N�}�*%������(���#�Җ�!�TV|z��wk_���G��8�Ϯ�o���`�U���C�=}�)W��&��W/�6]�&j�@�;c����ޯ!,T�� /K8��+�e��?iK2"�YA���AW6_�@k����s,��}�}��e{��Z���9�,s�VI���H'�s������Q(ķ�EF��#�p��Y㓺���
��#����0 �V�$V�%�	���.�2&���|+5ch!����w�Ji��C��b����4���3le'q4y���봉^ۼɉw�����W��tS�o���S�"�6��b"�Η�ѸYN�5)Rϥ1e�44������ތ�zr茼Z���y[u�>y��7�����:5�E �fv��V=���'־v)�9���4�G�x,����$�f��<��F�$�:��@�Yi��+J���M�ߢ���P�����wڌR%|���Yz��x���u���W9%~��yg9{��7<�u<��t�~7�� <�ｘ�b��G
�q��\FZ^L`�Gȣ�^z��̡�����"
�R`� 2����]�/;�xR�+>���$�}(��g��A��5�-Z�����Gr���Ц�����lŝ�sXր�TyP��R���e�'w�k�7�,�|�!�� �FXc��V%)D~����#2Kȳ�=|����#�@��]�
ZW�a��tU��S��z쯯�2�0G�����>�4��7n]�(�����z�։Y�Ƃ�ͧ��z�}��� =�������1�>�����I��\�cR�~T�	�Զ߭��W��jG�vs{��U����K��t���k�z���RPyr�
���N�cf�n��D���:�c���%����;˨f�~�5 �X&`����֩	�u݄S���h���o�����2(A�R�G�
%�_��T��Qڏу�p>�_��-��ֺ,`�$���b
z}-���FU#���:��4>?
�[Gk{T{vr���Lr�v�(e0)m�v��S�+�FC�$-q���K��\x��w��^6�e�67-�u\54m�x��jnAXȊ�_����=�Fn������=�LL ���u#�s���.��Gc�hb��I�+^"vp�����eTU��=B컇U�%��	e}�)A 9#�~|I����E�R�o3�S�ڳTz�����$��Sìx�խ�7;
��n"�Gwv��aʜ[ڟî��&�� Ц��Y-��2PU�J�i�Ó2��V���Q�m�nEN�Sn&�9�fhC���d�U�A�&_O�vm�I>6��О�?/�O�w;�I���2ؚy~���(۪��6t T�g-�^P��^���G
�.�۵��<�/�a�^r c�����"H��fR8�����6X�"n�{��p\u��C�*�L.���{-5�8���ڶeњC��)<g��8�Y#�K�.�^�����Y�Pt�m� �MA�'����f���B�Ր�U?-��	��q��'�a7�[��-C�D�o�=U2��'4�{�=���k�L��l�P�E����%��J��bû��̢��S'�2GU���Ϧ����	AG�{O]݋M"Sb�cVR>�o��G5�(Qx F|����-���a3EY�go�������1��K K����9�67�Fː�jIk�����~fnخi�^p뷟��X.���Ga5-j<X(h<�M��jM13���b<"4�`��ra��k����X�D�-�����k�ڲi��
�pEn��2c:��ܡg��ٲo�G����p?��<ω������;.�����B�)V�[��
�b�(bs�+ݖ��P�����<�'|���������j�A� �y\߿&�����C��A�O��@�ECNw��gQ�d9��K{W���|Ҁ��{��,���IQS�ʻ�s.3�g�Ө���R&1���Hi�?�"��RP�'-�*�a��`F��rÄ!�{]7`@�ZN�1���c���B0�:��(i]�����X����GI��p�]	��ܭ��,������]��L���啚c�Y��y��I0��Ƌ�W��|#�=4���c�H�-�B������X�^L룦���!����MorF�.~�b�dUј�F�ԻE
$::Q��U�2`�E�>`&Yܚ�x`��%�v�4�\�R۴-�p���хҨrg��<�A��܂�`�� F��3��5���L�j��E�����:�F	}{���R����_�X�������Q��+x;�y�P�>,؊z�����Xј\,���'(0�u-����R-���d�X(��^�p;��D�e*|Ʈa|�u���[�V������ }�R���<1�p�Ω3>]=)wM+zOa>�Wp�Yb���f��3��z_扸�T��k��:��>G�1�(��ӿV�\���&�#6A�Ў�0��(#��Cv�A�;X���5g-�A49ܭ�/k�<OAt���#���������[�[�pX��'��
H���=�Jx�ϕo�٩D)Ȭ�g�:�P.�9Ȃ`�>I}�yN��V�B����3��;��� Y
Fd���&J�������'�����7C�ME��AOyf$r�e�
Ī+��M���N��[N&ְS-4W�ts#_ �h^JQ��j6���｛]�I�\�C<^H�βISQ(:�F�Ү�5&:�K�����3��']�1$��'Z�H$)�	yM=I�@�Jӌa���+�I�哲�V7��e_�'�|U6��5mw�tqD�S��9�
o&��eo�y*똵=y�#�^B��e�˖!���7��G��,?F{���S�.[�D���8���2�����Z%Ƿ�3J����0��)�ͭ��ƮB��,�=%Y��:�����w�+~w�d�
��밝EGIT�f,�`"9����iM���L�1 H�!�T5,�t	��ȩ����.�q�w0R-��qs��?���lm0�lk�L�'��q�nt4�@��,+%/�#܌.8f�k��9~\Bmn���rRBԓ�)BY��xEjCA���%s���g
kVC��3JK��3oS����EӍ|A^l��b������(uVbW�q0K�ZB�ϧ�L��&`u��mb^0Ğ�DQ�h�P>�R��IS��d,���p1��4��h�-ֆ��r��[��8<�jk�ƳcT3y�А,�
J�r?�08�p��8/�s�<��,� <A�_1ќ��U[D���F��P������׳�Z����h���᪩0F���i#Dmx3�D�x�|J4qF:��ފ�vC;&'nY�o����l�1�&��[,w�=��"�7
�
$�^�:|�W�<Ou˸_�)(�͖k���d]��\�+'�����Z>�?�d�M��]��j9ਣ��.��Y�����Um��㊱}�>q%��,�!����u��>�}�ije���r}ЌV�Smf��m\�:�?I*���x�)����?���i�@'��W����wvb�@]�ſzj9z'���J�HT���$ 0%�9ޱpR����3����A��Y�̏�Ǖg��!,�L���
q�~�F~q<g��D%G�{OQ"y���%	~�(l�����@����Ľ����3V�������d-HIgIkb7�'S�V"��\6�a�{�
�wA/��H��ީ�������W���>�(3�)�b����qL���	�%��OZ��?[$.������?C�Q;2�h�W��'���"����P_H�
��՞a��#�-����~ݠ�k����mr(��%$y��g���X�3�l�h1�p1�Wؽ�P�j�]�3�%�h�38˫�y��2J��������6^�^��C����p�BH�&m��8�E��P�l%�s�gr�Y��_���h�S^�vާ��Eyp��H_v��I_Q��
�0I\�&?3���\���m���&=㕰�	��mruՃ��!0l=�c�I�E/=U�\��/Ð$�N��S=�h[��Dn�g��
�װue�)3�<�� ��actCT`��<��O.͙:��@EY{v4�W�e��L�Ӣ�}d��/�x�b�&�a���e�
���|]س K����鍝F � y0�&~$��6�ϼ�G�ݦ�W?(��+:u^�b?oyT�e��nS;$�]	NQ+����+�2�����*�<fP���
|Sֲ'T3�#z�����=�/�h�<����f���0Q��Z5�lM�pbm�Q|b�
�Eb������S��6���uK 0J�&�� �׍C���ʋ��_�_���w�\O �y���~�0֒�݂���9g�hT�௯=`\@t'qv�~�oH*%������928GGF�5H��Jġ?�>���f��ɽ<]�be��I�!]��J ~3x-K_P8�' ��_�J۰P�f��E��c��x~w��3\���أ:�(��J�苁j���z/B���V�� '5q���sԭ�6TJ��źd��L �("p��j�^���%Е
�GpAù��=��}�RPxq�8�a�Za�`�X�s�<j�!�.l�:�~�J�˒�e\��P=jFGՕ�\��_PlU7�;�
Xe�!G���=�����Gr�S̼�MH5�'��
\z)�3�¿h�F�yke1�;�ڞyo��R�ԝ�������w�u5�j��hE���k���Dť���u���������Φ���Q*�$%ӲaPR��uq Z���vn�q���4S�zO�<g~4Q=XU����~A����AW5�x��p�q�~$�o�N�-&�&���5�y��t�1�n�L�����b�r�dh���O�" �|Lv�g9�.�'����� �HN��z��� xA���+aQ`�7��q�^W�		9�g]��v�m{��;��m��3��#x�?�p K��}�AT�|���f�Ex�����tT?����d�0;/k{�\Ǥe����{!��J`B�Z	'6G蛋�w���3e�e�֖|���[k@83�q�hv,1��RjXN��+�!�Z�2�	W 4�J��4v[��^�[
�}�X5�f�5\s�Ne����Dx�l�=ο�k�A�R׎��a�5��Cu�0|��f�����bę#������-Xt��B �<X��v)�H<�y�\(6K�/7�a��+ ۆ�IJ�:�B��ZL��7A�a�v��-�bb��G֩By?�q�Y�8�?�k��/o:r���jAb�	����8��Ah����W�&0@�ѯ�/�P�K2Ǵ�h�Wb�M��`͜�+_W��S�[b���^�0?i��sCh3>�S�^��vM�FH5��?���HF"'��'�����K�d����m�5U��gf� q��[ �?K =I�Q�ƣ�.S4�k\͢+oR��T>j��v�u1INyeVҹ"2���<ϋ�?�\wyoP��@4}M&T�_%m7�1Re3%�ѥZ��� )��'u-�.�� L@\�� qy2d)�p����j�8�AF�Q��h_���ޔ��q��q�S�����L*���A l~y+��q�P���=���u����Sw.Kl�ڽ:�ќ3d[���5�'X䪢��X@{yLTW�Ւ���ZBɂ�l�{�s&�8fI1&���k����E�c�HRdǬ���V�#�_ݢ��k���hJD=ﾤ[e}��,BpAF��T]����;���u�6E9��q���g�lq���G*r�խ�7N7S�a����fB��O1�`�xWmg�̎D�'���TA���V�*���
cΟ��_�/=���X?\��=7�c��D��/5�*L���Y��!)9X8�>9����v��J��&�X��X �r�����|�?�F�8��c)�Z�ޅ��N�����e�v�\Sү��TE�Ŋom>IE���Xȶ򾦶���1? _o~��hXS��FUf�vY���+�60h���v�l�Ke�H�(���֪"ң�G�����
~�����Q ���CK3�5��2�S��}u=�X(civȼ�qz��n��>����V1]��Hn�2��ǏGn�Y����#Xŋg�6�ςP$׹�{k�C�<�ZS3f?�
��4�D�*Р��'�x��,���-6�rD�X37?tޏ�Aa]�!���{�����
�>~���nh�����w4 ������c+��X��.��[��keQhF����s|�O�H�ܓc��K��`H�����?=�/"RhI���'�	�jſ���������~A�F�&�V�Iڭ�/��\М+�t�UzO����\��*(ﾲ�L��n��Ap=e՞+�8��.4�TKQ�`<�B��#-AQP��B'��-�O���(������C�×{b��d��͵� ��6���.�|�'�k�����]��/� ���~�i�a�h��.��<F��"���[�E8�h�A�]ejCA�M;" =D�e�ˇX��k+9�Hq��G�Gڌr@����~�wA��G,��Z7*�r����*'�S�`�	�,n�8�^O3���hj۽_;�{Vf�7f(�b��L��"�-�d@x?h����/����6H1Ps�X%���K)z���8(��_��U�D0�٠R)b��K,��drQ\�(�?
���>���^a()�C[�p	UQ�q�����@�U�PF-�YG�ΈRz�S�,ƥ%~���V��=�l�bq�~���"̬9��;K�ڵ$��>^:[��l��4J{P`�6!�:^g�v�P~:駾�Ѥ�|����-P�T}O�"`����D�kb6�c�� �v�	G�D�2�X�ض'2�$�Ý�©o����ܳ쪏�P(�
�66̥W�kFK 
4��_�-�N��U��Ħ��.:�<c�Uvwk�6/��2r�i���*��N�h��\L�����'���MT�?Y_U�\خ��z��D��{�q��1,��^\�jh8�60�G5�����E�x�-�d���5B�"
�@$+e]Һ��Å�� ���I!k���I��,�#�p��v�Q��`�fin�(t�dh��ݡ5����]5�"�$5�`�t��+��[%��Z�� ������|S�e�\l�{�^�������ao����7z-y�ge=��Zm��\-���t�5��Q�	�����y��9G�[��,�<���J����){VD�TgeR���Z�2�&2l��3�e�����k~v�5�E�̭���x�� FM=�0Mv�o�3ӅM�@@'�&�]�3���m}sf�#��#\�Y6yH�����!�s�l���@Pd�_��.�iA% Y+�Z��M�m����:���{\}�%�����,T�?	"i"`�>,�Qڊ�u$[G��Z"^@��o�_CB֩@4�g�����s��L�Z�8X��Lr�mlT���y2�gm������sHS�O�z>�9+��ڳ|0?�s����;�L�-��<֔j�W�2��h������d�`�B����pp7�^���>
�nYO��r�J},���?��]�G�����y�����T�L�*'}0�/�TO�xBdN|�|�K���b���V7�ߍjP�)��g��0��7 輫"��ơ�c��eOI�儹:nj��Iי|)'�|Һe���l,�MM��[��\,(�����"WV�#y��gW7x\�
HV��y�"k7�����8?Á@��%2����CD�����x�㙏#=�(��K8��h�-�j��l��	��y���З�\Ԗ~l����џ��Q]9㰨85�3M�u.��"�"媉�?�:���Wʄ,��wWv*۫`g�1#�1���@O�Y��6_iw��I�����hM\3��whʁ,��m��F��(����Ơ�=�ye;kC�5=l�-�h����'�,�ů[�|����k*s�P>x���ɕ��k⬞OKܐ/Q��7&�@$} �eW��ǍG���|W��{@��f�p��>���Rb�b��KK��M��,�lw�]$�ܯk�MzzD��3�0)F"��'��f��m�|�Θ�$Zb���kE��h��D^r6W�H�Щ�I�ҔT +]f�p���Rgq4>����Ʒ1a��X���J��F��a���6e����iV�=��i��q��%��X�)�}��'1�fC�Ѫ��:�&�+�Ld2����4.��N�����e`�L(B>6�̀!M�^���GA#��y���9^2Q����N���Y<v�foQ{O*�׸����u(���޺k_+�̆~:[h�d+A ����S���sh�;d�6����l�o����.ݿRf����!\� .��Iy�&V�"� �a��7; ͳ(W�(�
SN_����֩cOd�Q�	0�("?\�Y����Qi�]	�W
6د�P�&��!
�e���_��oi����,`���]�ʟ���ØI�L�~;��Y-��R2�i�v��_B�=O�a ����U�Vr�`M�8$���.�k�*/����
\ٯ�H���֖ѐ2��~��GK0��7)��h�
F<WՎ2���t�����a%�H��|���vt�(-6^���TF���[��L�dno�U�N �`�I� ��Pe�߂�iĉZ���8��-�ys��f�<�������d��`^���9�B{Xh�*��yG�A������}������ߗZ&k�����g�R0���J��b���K;	/C�R�N�� �W"�uU\�l(�_P��ė���6[t���n��	�e���m�3o����f�������f�V�"��l�4~����%֝ �Mfk�rd�Nl����`��]�/��8��LO6ӯ`�i^��Q$)���:'�IpI���"	�=�2�2�c�;ь��w^Ĵ�10iu��X���� m�u+/�J�����]����v��؏#9��)�?�n�d��ܻ�V�`�2t�/�?� a� 0�����R����>�̸׍;�9���� +���#�i��Bo���7���������6�;�\��c���g�)��ԎO�oK�RB�j�X����.��o�'�qRm^�^M_����z���u0h�Z��7�7���ZJf�*��(!N3=-��Jxٷ��1�`/{:R|!�#7�mD�Ю�WtˏR|FR3�rhW�&X�e�}!�8�e�Û��뫓���3��T��$\Ɉc�@m6w�x��e/D�0�/�%�#�T/H5_�f*���I*�N��1�3Uqo��Y���{�`Z�I��T��BT�^���9	.��8+�D~Ȗ�;��0�
������P0M�o���M�4�wK$���5 눗{PA0XFW��I��ġ�[*�e����{��*��щ��\�����x���V��Lk1�����.��Ѽ3�M-�Q�`���E�(ZM���C�N�Kf�����\4��#j=����@R�*l���q��4�qA��A�kJ!��(�����D�雕����P�b��8��v�S��U���0�ҿ��|��g�r���/���4����!W���0c�7��p�����K�cB������Ƀ���ʢ����ٚW���a��ant�x�Wҿ�b�C\j!7���w%)-W� ��P.�XB���n^�����nvԪn�79��w)`i��5dO�P!oC�c}
�EŔ]���v�z$5s/^���	8Q�^��P��x=��`�铳V��΀ �`��)���[ A�^!.�{w�K�B�m���9�p�ڷ�BGK��R(�f��G;��L�2E�CD�G�_���������0�bulEGj˓�ꁮ<A�d���&4Vy�c�\,���/8prk]j��3Ԗ��ٵz�<pU�+��v�]~�fTߘ�A�n��FՎ�u8S-���k�g�Oi�B��N�n��##M}E�g��h��]��(mm�~��X�L~5�D�^���\4D�0	������[�<(�)}�0tξo;���%�W�Q�����i"�oЈ`%���� J�4��ƌ�5�mp;�0�Ñq�"삦9U�P�7]�a����s<V�촹�*j�]�?^$��.��&�~��]��u���V���6�헚�hQ���D��j݊{����M_�܊�<)e4\@Ti�jj}��aP�8:~�gkuK[fX�CR�P���K��x*pZ��+�e�lgW�:d���?�\�� �;�_%Q�0���9��o�ٗ�e��\��M|B�����U���<���v.��P	�(f	�@���X�v�ѡg!�iV[�DN��|�/�.��&C�D�,l;�#]��}l���'^��^7Aq��7ӱ�Q�Z�|k_{�{	�(؟�'d"�Kf�-�M%V �G�5�0U�t2��W�hG]��)�Z��&EJ��u��1���%��G=(b;g��3��iE�˄����"�Qӱvrɑ��9P���-�,?a�/pW{j;��?$|v1�RKE��>1.�߰�CNIq�	(�nKmf�!����͘+|F�{�uT`ͣ����� �H���jȤ�kh)6�&N�Ll�q�ɹ<R���m��hM��w���A��:o��y����EV�Y�{��f/�+��S�A���� �I���s�Ik@���/Vl�gؚ����߃관���;0M�2H<�����pw�qMUYS\p�4����aJ��jaӋ��N _�Y�@�i2.�@��ap<��+ZԆ�H����gRT�P�f�#B���IjI�]�Y�J�3m�������1�X�J�l��,ť'q�M�cE�������aG�f�|K�i���5Ѷ|bȒ�8�1�B���c��!��ȷ%-�P�/������}<��8��0��vx	���lO��ʔ�\���j�XxO����y!���� ��5-d{D���l�t� �FhY��ozP����� ���J�����9j�$�Tr����V�KA$��&�#b�TO���&�w�2�D!V�q��	^�i�	EwD�0yよ�!���n���&,�5��I{yU�l��l�5����"Kj�8 �U/ 
G1���#�WƱ��:,}:��7pr>����~�/NX%��o �OS�#hϸA�w)s+��P�75��I��˙o�kx�Y/�a�#�2��e	��Vy�fW7�Qi���T��o�ҥ�m����~�_/@�1C��u�h�{��e���d���W�_��)-��7g�a����$���~��1&	�)��4�:��Anܐt2:���u�|G~/Q97�����W{��	w�>�@��j>��a���9{��H&`A�;�=)��T�y�t�Fׂ}�U�!�����c���<��)���.ksY	�#v��)�~|�`7����V�LxQ/jY�M��yQ�*iÎ��j��9d�
�����f���dF;ZLS[�ñfۭ���� 㧢L"�ҹ����:��wh�8Qt99��{�����H���@*7gk���5wm�4*%فA8�bA�թ�~�T
�D�	5�oIX;��<ޜ�3�h��I+y�8I��h���?���n�Q�ػMv��$���dS�S�luJ�L��:%
�l
��(�g
��&��V��;�se\�W�1�������38�]��O�깷h � G��E�[�l"��L�U�Ƈr*��M%rrL�pi�~������q;d�m�"�v�&�maA��p�Bx��ީ���1��������S&1� �����S����������h2����c�P
���$7��8����E��h�hc�V	ˎ���w2����r��=�&B����ֹ�� �Ŷ[R�蛸�w��f
*X��7h�>�{Y����Cr�D����!?�Zx�7��ѣKPѐG�&�#B7xz%/]6D2i�H����H����-�N��?��Y�=x9P8T��7���#�|�!&(��7�n���L�K�`}h��Sqt�>ɫN��?B�����'�+�˸��e�[�#ԝC^���4�
�nl�;O�oi�B�mz.}����$�;��l�Y��%��.s`�V\Of�l�bi�\2��,��7G��a x� *��	q�3K�Ҁn/:��$�ҵTt����b9[�-���v�o�t�0&��Z;E���ޣV�
���������U��1��$�T���s�I��I2���u���V� �A�_o�V��k���gsX��ͱS��iJ�T�[��G���KM�?���m�ÒE.K�������Ѧ��kB�7Jy��B~ C�Q������N�V���楳�8��`�f����R��E����ܽ�L_g9�uxy�-8E�p��^4�"�D�?�I�/���r�T{��1�C�Օ1Si��)^���H��ҙ-���E��i�~�;�J�R`9�$
~�V�J)D[����qIF@7�U���@���w�ޱ��"�+3"������vfn�yH=����*6SA+���Y��jGbb��|+���횎l��|eu��K.�)�e�%)��}e���}e��Ϧ��Ǜ]���j3�5��������c��lf�l���Ĝ�K�A�D��`�©�q�)��&a��Ι���a�FcA�j�0fb��g�Nc��QG'~?0ĽE�v܆��#IN���G�2	�
�xX}��)�_Jj�5��9cG�@�AD������l+�?.�T��~Nn�G���|��ILHa�\D=�
/��3߭�1�/#�o��9e��}/�u���FRE���q�;9��U�[���8A�ף����N�}���|5�^T�Y.���Z�~�`�6zdC��൭PLC��D�;��,P�uSr��g�^f��8NZ$�E��-e���}I"�}v�U�I҄]�[
���!v���k�S��P�D�R(�@�ZA���J�c��|�ye�	�V��c$`8�2]�&������#Ѱ��'	�[���2w�d��ܶ���q�V�P�1���|B����8��Y��B9F�J\*{�V��J��xR�G�W�ߑBC4��0�"ü�����&X('��DRw[`Hv�*��S�"&r��/
pw����m=@�ڌ��YЁ����8����Jv�2)f4����c� Y(ȅ��֪W���������^.����N#�@V�6 ��C��\tc���l�ũ����' ��#L��8���ND�=b��Ȓ\qPJd[��Jx���K��g��p/�1;��_�n���*�?�aK�t Κ�rX��>���Q�0͓�zاt=ʁ���_�ꇲh�����`\{�~2��m&�}�5��3{J�b �@������A.1�R��i�d�zS�-�S�L&�=y�LJ�����q�JK��j�e�3$d���|N�!`�0�m���/��
ٯ��)7�p�1��@�H�/�}�����wю���3�yڡ�9,�I��%
�@���L���F!*��1�O�o�!��Ǜz�ϡ׋k�k��%�ob�'TJX�J����r�92������ץ%;r�`��2<�#^#7�όj�EA����őhY/
��}��d���]�43�O���i��?��)n��"��x$��N�<Hk��̭�ݿp6�P��V̌��[0���1��ӿ�w,����kl�.�"�FO{4#*��=����
3�b����n��3)v��%J���V��/����y�:ہJ�l�M皩<����ǖc�czQ��e�8R-ZǞ�}B��E����|���u�K���Y�W\����0�ĭ���pA1���dZ�e�V
{*�ˍ\^=��v��`��Q��F6�lN{�����E���?�y`6C�w	�畨��z%v�`���a�Ղ���-���S��D�ʷ�e,=z�5�����?AM_�ZmHiҒ��,�I'��titԳ;%�^n�/�F�b>xm���y˯XBT�]ڀѣ�nv"��?��;a��Qp�� ��txg�Nb>mehAQ�"J�x���;X� ��BL��R�J��a��g�w��u�k�4b�c�Cǣ�'�)�Wf#\��Qm�r��P_a,��4�>>�eW-dr���[N)u��X�@J&A�������� C)W��X���\����������|95?�Fy��0�ȒFws��������Lx��u����X�h�	��4���h��Uk�ܒ���DC�N+���%g�I0��?��/��Y��R�������Y�d��s#�� ���BG��&Wo�n�gk�V
(C���(�*�q� ��PruM4��µ?��>o91z�Yo�����~�Y<��^�nXBFC<Im�M�j���y�©���|g:�l�����3S��@�/���k��UC;������7۵�s�Zy~c�����*Z���;��~���l��L.�GO%e��(/8 ��s�CV��0�n��Fn3Lب`{�����0��ȝ���wn�0m��D@+Ղ�s+'02���G��'[���7���/b̼��ĉqPok@��� t��أ����u�e���e�7�e~y����	*��m˹T_�~�5I)~�6�9��>AH�`{����i���N"��i^�
G�����ܚ7����zX�e�刎jȳ��^�ye�#E���/�-ɘ�7)��ϣ��^֟�"�,>_ͺ}�JT�w;�m�l䈹jw�C�"���q�*o��/����5y;QvK�lr�����0V^��X^���ɶ 6��ٮAoD�H�Fr����x2R�p����#���W�	�G���l؀�p"0�o/�y�|��ІE�t!����C��S|��T���W��ᤩ�ǖw�is@���洓T��e���Kg�j��"�K�Q�`��Ʌ!aH���%1�5�s@�GY�f�v�E1�,b�v�%�t�Q��r� 7Zu�q�`��e��ζ��W�#��0J���$6IoT`2�;K�8���Rj�u+JX{�H��.�B���^Å�'��}`r�}��뛍���k�W6���R�_eF\cW���r�Yv�� �2}��(�b�vCf0�y��`ΠAxs�=���*h�"�5Oh��0��N��a��X@�~�N��K��ϫm	�^XP�hp}^N)|?���^�˴@�#;���`�fS�`F[T��8B�
S/=া�ʌ��>�fa*�̔���i𰲴W�����x�H��ǣ~?��t6?�9�c������q_ʁX�I�=Ѵ҅����\��`�H����qm
�7���d��[az-������g#!���Eͪ�WM�ś�_�0�`�]�F#e�ת��%^���a)0gIz�ge��&��sBK��Uk��|čI3	�qo�F#��[�)�U�J���@�Gvs,�QBI�I��K�����Ab Fï���/��L��	��
zH���j��Ws�E��t�5� �����O
vAA��ofE����8�f4��( ?��9�c���GÛ��[I�d��oR�C�e9��oMq��a�P�-�\y�N�xJ)��Mh@���bȌQ_����-�g�\(8�4�Wl��X�K
�����C�u-1����7S�����S+�쉭j=�c�UW���9&]=]���C��Y�{�y0��Z?!�d�&����("&��
�^1�?R��0�1����M/.决�^?��]jS�>~�|�Kt�q�sS׏5��s��b�zV��^�Y�4޾��blMg]�2�9q7�����g��q���OG��z�[�d�c3�96,�H97������o�9pOI�w�}_� ш�)�Lj|YM\��osΓ�g�����y�S��&�H��D����ٖ��,�8�$/�z���-��	!�d�Z�	��+@iK�:�\�P�6ٻLH
��^�nOl�0Z�z@���%�k����`���H8�sn���� {D�z�|Eo�۪q)J�`�BJ�2���p
9qߝ� �
����wQ�Q���z��>��'�W}f�6�YN=/��<_R��e��6�*ur#q�f��(��c���&���d��11@�F��=s���[7�u�E��ҿ��$����Fuɢ��#B@��Ġo�C+A��Iu�f��@��:ظ�?�Ѿ���=��u�Wp�7!�<�Je��r֑a��<@��+j��t׊�c�Z�>��Y[�w:%��Z�t�9h)3$˄X���W�
��򅒄)/���7]�`����F4�fx�=�a� �,�-a��e^�,ꮢ&~Ȝ�q�_=xk���T��d��xJ&�(�U�v{�%�PsuTσ�>�P�&�YuF��r��o��3���H~�Ҳj�y�s&�ϟ�.���;�Y�-��%@U��Xtt���9~Otn�ǣ~��d��$�Ui
����3�����we.$�Pc���ӟ�@R��U�6�Չ��	����r$���y�"pd9����q_PLrJx�9��~;��neٍے�t�UM�{�w�a���i���}�ri�%N��� }�vj�VCO$��� �I��ŭ�C��l�9�8�[��o�U��NkG4��]�g�mM`Hw��h9�`��� ������zo��+�8]��|��p�3з(��)kIv�xf��E��ւnʒ"��A�T�8G���'�H��3D�]�%	��΃Y�<�]�/I�*;(�N��ƺ#�L)ra�&k������=���~xoA0	��
5S	y)��Rh�j4vf�3R�_�bH�{��K�G�Ʋ��,�&�4c��]�d���p��U��@ }?7	f�d'O���D�}�2�1���p��k'��n�I�`{)���D���>{&}*��"�066�+�y@�����Ѝ�NC?<���b7M>j�*gv=��B�N��ֆ�_��5A3�n��Q}b�VKѶ#��h73u��ֽ�1��)ݨ ��2f%�p�<q]I#��B\��R���=����Wei5:	1�/�9!H(*����B|�u����;�/9;����^��y�]�"A����b�^;Svg ���dC�Ѕ'�R��a��H0h�,##8}�"Z'������V���,�<�	*5R��œ�� ��1[K�}�B�Eex�ap(Z�l@��������c#�NGo�R��Սו�oD�.�0���D��X��1�9�s��w*(��E��Ɨj~�?�+\�0�T�@���S�n�:��=�<uW&Z�^�h���TY��菿&�,�8���n��v�f����챺�k�A���7�)�,�����TJ;x񦸐�t'�Ȓ�W� 5v��JB�|.
�� �1���W�`���3�7��̈́��j�I�9�;)���fY`��h�jhkܴ ���pB�JǍ ��j�Ї�q�G�1���� ����"����Y0�d�Ϊȵњ��B�ޫ��Bkr,Q�7�f�E�yN�8l5�u�ˮg�ˇ-6��o?o�����簽�#���ǆ�R��ԏ��=�j���P��&̂&(�W�2�B�[P:f�&�eo�a]�%^�iP���爈+:X��ۥ2���:=8�l�v�5��� ���ΛߢE�Ћ��.��P;g�L��V�|5^!C�U�)��@�;������,ͦ	0YEi�ou�_	��9��*	N��_�p�@b���Z�,���	������=	8�������T:'����:����3Q��g��i���O+�n_Ih�\F��l#�]�� "�\����V��U�}U=�Ĵ,���j�fͻ����r��d��Ї&
�_�O�~uO���+�-��Z�Ɋ��� ��O���;�}�h�yo��}�0)��M_��Mu�u!3۶���2�V�ˢ�[K��Yp�)��!u${�Uв{��s�N d�V7��ٳ#3����#	09Sڗ�(;�ݢZ��-�C�%t%�p$�a����Y ����Z3��K{�e����:l�����c�8��}bPU�t��y��SGG�S�5�'ulfv֝jܷ���n�k��p�S�o�������W�ZT��V�녫��8a��tK�pۯkK�`�F�uI�P��G,�9����f��g�o����QR��$�o��č���-�4`ε
Y�08�_�P�eI��RD�|�5q������;s�_�'�)���?̕�����g?���G��R
r�Q�A�44@u�o�!��<NA+����^t2�G!G��+�E��:L�i�$�ʠ�����X�n�	����3���&�1�@*z��ڧ�L\��r"�b�೶�bs����5��+X+ 7F�kI!m�X{3���O��+�K��(�:�Ѝ���<R��y�E����'�"m�C��9!f����͋\:�c�u� ��Y:{��[ԋ�^��|��ﻟ#3��.�`��,Ϧw8J	< J�����P�@�t�|,k��=(Oq3郯��<fG�������|��5�0,�H�IXJ	�Y>oB�W�j�(v