��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,G��U�	�oJZ�@�z�����>�� �F9!�/_g�T@_hm/a3^��(#z�dZ�E�����v�h��|���-�>����w,.��N����9Z�S�p�ւr�p^������[�G�C-�Dʩ/�Pm��[o���w��ׅ�-
G�)%�9.�eP��0�Bou��#�{�@�3������
�1|;ku���'�7�O���e��˗�{�$2�\���θCn�ob	A�����i��+AH	(&����;�gL�P�N�,ʙ���A�S��h�0.ީ#��=���t3�e�7����WmN��rJ��ZՆ՚=R�@��'S�s�*�[@�C���[zW����:b4�M;,�Rr=<�z���䄯`>��}���i�ƝY�_�����b�w���nӈ.��DVHx?��\�d�g�i_�3����,%t@�����^�H��	N��7a�f��<�rw�*����ֻ�Tg|э��"�ׁ$&J���P�dp���f�:%��|�b�2pi����I�ȏ�֓�0:V���4*L]���
��(�͍��1�O����~
�<ңy��p������i���/jô28�.z�Y�?}��cAL�6x��O�.�,���Y��k���T��� Z��>���yIK�����ҕ�aw��@c����L��z#M�9�ECbR�G��L�<�S8�ɿ\c |`�61�=PV�4��P1*���������6��7cC��՝�q֐Yy_�<�/G��L6&��m���{�����?�q�+��z��?�N��Y(���&�q��l��4���sӼ���Y���D�=��`�x..�H��d�,f����%�����ض�Q�n�'=?��r�R�PXl�q�|"���@`��<�O]�����]ՒyH'����B�����Bl7�k\�¢���I�]�~�q��̼��mAy�V�D4�q���_�)Z���π/$�`O+���p|��!H?�>;��}��b}�GU]�7�~�=��G�IМ��Q�s�!�%H,�|� �6��������Q�-P"�����q|��
�z���&����� �cUlY�%#F�#�i�mɬ�q��,K[[�eW��Q�����H�:!�/!���%l�oI�������1��۫g�HG�����g�e9�����V�}��n[�c�n�� <�!j�s�e�#jW���KTz���L���	ۙ�41j�#��VjK8�ܔ��^\՚�ׂ̯�0YI�#z��5hj4i�K�ʟ�N���Iszy�Ϡ]L��lw����v�ف��
w�
ky�sݙɊW��&=-})��<�y��~@/��wNZL�5���S8��f�$8W�n��C���1�.�owE�����l������^������9<����r���-f��۔����@�Y=��E{3���-l��n��!zl�����{_� �h�0ʃ�
7�>6I޲�����jRϔ��a+�Z�	�D��T�,�FUD�,��I�N&1�ϪZ�'ͺ��K
�o�s q�("��-��<���m]�a�S�ɩ{U��|�+
�<r���u�P-� ��g�&�i��ա$4 �t���X��[���R�EȆܙ��l1�eDgEp���{���b0;��-۞���^7R��4<h��ӿg:ή�/��^�����ਦ���/-������Z�k9X-�~��;k��'7���vf:��
��H�)�<�V��!�?�@|�d�F�p�T��5'QI���]yZ�'$v�C!��-�7�}'�:�㷾���M�"/��µ���b�ar����\��
 D�$�KE��v�5�D��������[{��rͨx	�JChRw.�޸��a��A���`o�;[L6.�0�=���r5$3��ǌ�ct���f� �$*��tb�h$��</�Sia��?�,S%��Mi��-��A��m��6dK�0�{�����P[����o"��Y�M��}���G�}v�/�M-"�3�V������s�ʃ��+Yq�m�+>��Bm/>ކ-N��;l�����!�1y'y�W��ۡ�Zr� Y�^�������&���Y���<��*���JZ�0��}�wϹ7W0e`[�MJ[�����%'^��G3j�=g~MăؚV_?T����;6r��Qq��i�g��*��W�n�r�*�qJrPDR��X%U�orV��2~��������L��MCF�6$&s176�Ɯ78����f�׭���h��n� P��Bt�e�c&�;Jk�/O$n�>:]�ʢ�r��۵�d�Z�K�_�[܈YUc���}`��4S�92��bꑾ�X�I��/0`v��p�d��Z�bp������Gާ�Y�CC�q���!/[�7_ .P���s�?�q��%��H�9���zz;�D�ԅ���i�?xڤ�ζ��B��w~����lJ��Ԧ�B@���ƒ�@*�V�A���ю aCMfh�"�o���79�N�}/�^�C��c�w�Ԑà�.��g�/~�9�����ւ(	�#�/>�U���O_}�<t}�$��?`]D�"����ڻ�M�����H ������zw�2�~a����+Hj-p�{J;�ޙ�y�|8��9�Az�w�#$��ߵo$4�U�޾٠"���1i���"��.,��w�xX�`��샲%1ִѩC���
�s�{#�0?���S��!��ɗH��w��{dy��ʿ���2#��.�;�����D+Q�,S��T\���|p��{����!|���dV�aʖǈ!�����<ZVc��2TS0��]P�(jG1���N�&����e�����]�,p5Tq���Yi{C.��w�P<e��S��K�j��1��1�F�K��K����a�8��/�䖛e��
�S�~��U�[�VM���.lC����ylBb�3����@�*�&/ח"�E)�g�I��Ep!R�����}���@�˕Αo�g�4�ɾ_�2���Zq��U����ޭ�UK�-��Z��5p`ȝI�e�d�%�ë ��u!�K�Ց��N�V.��ݨ�:5�_t�k<X^D�0�u�tJ4��W}���e�^��\$�ѓe{���=֯1�^:7�/�08BN�2>iw����R�c-;- #2�"%`[��`�����I)�D}4�t��meQG�j��%|��fnF�u�e'd��k&���w�Ǯ����טkk ��	h.�Q��VaAa9^c�)�#��a_�xd+�*�& ɬx�X�+Z~v?��!D������B�}�m��}U�+�U�+�j�bk.\}�|b���\zxi5����� ������3W
bm`���޷�&^�0�8�U��k�N�2��
k���V�9���,S䀙�������%j�E)�������}�ֆ��t_XY�N��:x���D�0[�p����F��0���Z+r��j;�6۠h��#��#��9Ц$^�؍��m̑�M^��9�O�%.3��:aB ʅx��G9���.��uQ�3�x��ȑ�pd!���%��E��	b�`s�Jz��(B2�iq����[��+X^�gY.1����R�r�z)��I]A!N��G���X(7�1���[C��q݇���cWƆH����3���L��!�����
W��@���ʉ������E��#����օJ��0�X�N�.;�7d��[e��L���W����0�X����ţi�z��`'�.��śȠi\���9l���&���Ի�1����Gw�ߠ@@h���y9Q&v����l۩���T�b��=擆�"N��0D$yӽ��j��Q�j��u]���E 'dS̍:=>13"��G��1��������Z�9���#Y�2&��l�\]՜4`]&I��E´�Cs/H#��{�g�o���TUz^4�%�Y7� k'���e�=13�=(�i>�d
�P�|���*� [�|w�el��~5��`	#鹠�ͼd�V*V�7��f����@�0]l��ZV�?y���KW0���m�� ���8�:�2�P!9?�>Qd��j���kŞ u3ͱ���>eG,
�'eX��$�87(�>�DN�gfx�Ӟ �ۡ��R��}�yvI@��R��L�b� �Ws�d�u��c�>0��Z�n�����7z�..2���OO=)��D�������� �V&��ȗ8_z�W��.�k螃C�p�j��?�7��[��0�<���5�j��q�u�[�<��ʴ��ǔ�bGx9�$Ζ�x�ibc��J�2�W�qQ�4;�C���X�m|