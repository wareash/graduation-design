��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jåا{�\�u�?߷�dn@6�zf��r������;��r)]��*���/�����l��%돆�]�'���4�a���7k�'��W-�I]�o��wyB��W
���t_Y���M���GoS��������/*�c���^�T�j�,#r����!�P�(r� (��i5=
p�}��@�cRd�r����"O5H�ܖ��Z{x�6؜PB+ǽ���w��p�>aC�N��*��'y�ՙ�k��}�4,��M��[xe�00"�Bw#+{/$�A�L�@�.�K��OB��&2�+��$�8�9��T�y�{2;�V�����K�l��F�H�,�#��x��y�D;��O�!B��>�k1޵�#�{ �W��7{�1���d��k��!N�mL�YQى����/��E�w�/�s���j�;P-Zp�	3Մ~�y�����ɶ&Fք�%�3:�O8��4�S9�'�hL4���;0�:�k��䭉{�ǀ�/8aS��vL|pʶ��'
rU?��&��UHe���Yv`?wh]+��l9m	;!� fɥ&�KH`��l����(Ő\��4s�5Fؾ�C
���e<+���~X�T��XW��4��Pm}֐�vl��u�Q���e]n�b��.�MF�B$���%z���+��y�����2~���ZM��㨲X�l��`S��'<�>eL�).`��8��U2��4q�Q�a���Z��ͯ����J���=d�c�O8���S]fm�D��"���	B��h6Sr���'��¿�kBd��Ί�Ri�\n���X���c�JRC���D@;]�F;��s>�B����gg5�TR�NAU���ڻ�3�C4�#�@����� ��U`����������<J���F"� ���
MBWִ����gha�X��=B�W�j�W9�����7O>��z*�Rύ��(���F����@
��$�����F�P���@�ɠ�j �(RE�1���FmXƁ�k^�1\q����w�-Kf@{	�4y�w�����[�1�2Y�����N=��z/2�c��C=���ɜ�z�Z�x���Ag�rl�X�ϡ1�k2�-zJ/f����a��ip��d��Om\�.����Rt��9�_�,T�ce���̼���5�`�^���M�6������?�,M��%�4Ѫ��Q;�f���W�Gs�y'FX4���\wd[�Wl��%�w}+>��CF����_��D;TЦrP�*�T5`#�fv��nٙ%�U��@��q4��w=�C�\�ʇ�d.Y|�&Jvr�
�}$��w`�p���s���Y�t˙��u��|���IA�����+�e�>�(�h���ڇ�	[u����O}� ��>B �o.�Ĵ��ƚB��G��W�oz�]K;G�U6h �X:Ъ�y��0e�Ú��?j6y�A� u[�PC=��uw�
��@�Ɋ5�1)��?sA Bt��6Gwo�X�p�%� ��O
Ҵ��o�$�{|cW����D�x��ѿ�)�r^MōQ�۞�;��+��AT�4��W;���������P�$�A���G��?��h{/�E�f�R/q�:ւ۱�s�里�&�|oZ���Wx��mXI$�ک�p�q�j
�f����;j���Q	�S�y���Wh�5��w;�XE�v�ȍ�S�yi��s��'��ַc1�h�+��i�̵i(~Ķ�-��)�N�>>�x$,��JMno%z��\|�����*��� ���93�&�E��үS0��lck��{/�)��C%���,��0���|�����䄼,�A�_WW$N��5��ar{�W�Ĺ�c��_���s�N���a�bG�?�G8+hf��}�8!����/�zG��4�+%���a�i�/�x���h�-O��ߟ2��_��)[��2R�
kh4��`��O��&��,4���
9R�	�t�k�Y����ν�(Qk/���`C
���X��:	<*�nUM]eˆ���,��Qa�?�qw�ڰy/�:��0�)2Z5�@���������.�&���	���Ȅ���C��B5��!�_>@G��׌��$���.�*�Kt�{lޔءs� *jn(���O��c�����u�I����� ʹ�?��>����Y�I��M�> 7U;��v�q*aox�=M�Yb�N å�#f8�Qp��#,��f�=��\���b+!�B��ퟦ�ꈿ�'o�L�d��B��z�t[��nJ���η<�C��
��wȲ�_��W�u��`,����<(@��LAA���
�,۞
��A���"�xԻ�L�~Yh�P���еj(��d���	�$�����`��>y��`d��)�b���T��Օ��d��=�#1g�_��z�p���,��U�S�Y=2�|��)�LB�q~�叭�BV)�0�	S��v6;��>���A���5�j}ݬyb�z�
߻�1�0��E^���0�R���Ǽ;��M}.��Z1{���6��)�N~��i�*��#�:(�}_�����0�S�E*���:m،ey��GX�B���ء�{!�Z&9��{��Sh}�f���e����9��5p��77'���"�#��¦M�23��=���4P7vG൤n'�T �T�.m��*I�c#�|-[x�J|�j�����s!�ɭBFƄG�C��Q��W[D0���K׫ր�Ň�u�D�<�"d1u$pb:�8����*���f�~���B���k":�k�lԊ��U�'�m��ׂ�L�� XR��u�����B��+i(S����y�CG[R�S*VWV>�N��7~��/K��V�jFR�T��(�������	� k��(����7ܞ��:Z�RRsу������*�c �h�(s�jL?!R��-0p�J�!��iJ0^"=��t�kJ���Uk����'e�<!j������/�x��9��16"�[^I����>�$�Ϸ��7��7����t�?��Lku�*�B��@�Ō���sUn �NYc�(Au�)idA���,����.�ۇ����wő��(�{��w*<g(�r��CAnEo"�\�a�B��ƻ�e��� ��(�*���g�K/�r�]����}�T���t��(�J�42Y�L
1P�oa��Q�$�Z�����J,�s��	"�(d�.�� 6Cd"T��y����b��LK�����Y�Q?#X(O�DN�t_#9A�y�:ދN�ت����].YU`}���|p��$�?�R?{���hX��w�JȋA ���,����s���ﰳf�hQ;ls���*�7)��A���/e�"aT�!<�������i�!%�F8� |蚐 �^�c �:�Dȏ�
�����������nT@	FcћU�2�@Piv��3`�Q��Ɔ�𧥭#��1��/���
�(�H���_DK�=0��=�}�CJhhr�wU�nH�q�r*����{�bW-����[�����
ڀ��!�����kA�/��'�^5�VM2gUf�S����vd�[Sl�Π�������I�E����jB-@(9	뤊7�ً촒��Z`�{�= ْ���y���q���]!�?�Y�����z��lίZ�]bg�T^{�Ƞ-�6N��R���B�*ݯ����9�h��l�:��1O��f�����?�2U����r(�[��x1f_��*�B����fa'OEݟ?��-����,����Ad�@9�p:��b�vx}��p�	�1j#�D�H���؋�RRM�7�x��w��㣃��%�V�"��z��yP��u߯��Jg�6z�����e�bR|$|�QE���i$U>���unML��!~�S�`�ߗ�3�a̬͒=_֧��Oy�Çe�/O	@��xU�
ϽsI#P.rY�Vo���'�z�q���;��E$��s��S3��ю��['i����Έ)���0�&�>����aH ���e�l��j��gt����g��Ezo�x���<����@5&(#�\jFe0e�59#��}�4F�m�Cnd���`l��x���$��Km�tꋅmD=�N�B�������"�O�\^��Ѫ��A�ux*j�-q��^�V���4�Xmd�=��D�c&��}�O�,��jǭ��bG:������^��0������&h8x�Քצ�)���**�C�/�U������e�w�hA��._ާ�Ri x�[���H"tO�j�>3�ޑ��	�K��k6��~��Mcv��{f�cͮ�6�,���<C�^��=Ut�5S_�� ��1l[b�X�J��~[�S���۟����QEG��Kh+�=s�v�ڈ�(���N�oP"+s��\�ܢ*�7�4�N������тv4�'��P�a�o3'��?@5�z̅ȯK�9���&��N�P���Jw��%�c�sYh�>��0���yBr�e?UMK\�1��"����ij��R��w{r�ocH�	ޡX	�<�v>��b�����3�����?�C��#:H ��j���ƾgZ��@�_��K!�<�X����`�)��4R>�$�rB������K�-{)x>\aN���Q�*�=5�:�3S��/"Ֆi\��"Ǣ�U�<�J��3��A���rA��ˏ{]J���o�t�c[�)��:��q��	�ZY:�LR�%�����_`6	pb�)�)�МV�_��!�?<8��e�	]q��T�1�A��)�Og�xIk��/��+�&*��8�H{��r�#Z߼`Kg7-*��2�$I ����@��س"�J��ΞƿcGn��J񕑔K�P��_��q�h�PB{�WA�w�(,�g�u�B*�bDe���2�	���H@�bocf��-v��g��(�����ݔ�Y�a����
A��r��<@ܢV��)�9Vo��M�R�(iU�1f��E�3 X^�O�3a��V�����KE9j:y�m�Y�L��f�x�R�
q�K�қ��2j�w���ϊ��9:0V�E-�l`%f������hƱ/aM��\	\X�n�1=�~�R���yF��!�?aA`E�_Н��[��^_���tw��b���
�<G"�*����oJC��G ;cR�( �R�t� ke��U�M 3��&�ZvN��8ѤF�ܛ{�D�����[!�[���T[ ������+*u�5��aD�9�I7��Nړ^��Op�c��|6`q�e���� ?	=�a�������=�
!ɕ�H����	.Y����քuO����g��UB!��"�k�yw8u�V���'�i�u>�Z��ZI��-N�`