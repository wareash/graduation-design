��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>>�Htd�g�����B9N�ٟ8R��tw���SG:1����HW0�ʿ���J���1Dy�js:�^ lq��U���\j�R=)Ԓ�Ƙ���}.�h:J ��?+W�醬)˔bZ�K�� �6#��%�Y,��������m,�*"�b���c��2��l��힬�%=�Nd���|_"g��(��n��ցu�� 1-�j0)/{�QvPM��_}Q�&�Te��ힺ2�۱l3�a3u^3�n�U�Ic���%�<N��F��*	��lgF����]=�Q�{���C�L)L����Q�i[Ň���
����b�[��~v�9�y�Y[�J��۷:̬���cQ�s���Y�_?i��w��;�>�9�5ϵ���~ �������s|��Y�+V�$��ԕw� �w�1?j���m�ʨ�9���3i3דy����x����ڹ��|ΞUÀ��,��fS-}ah�"(�?z����|{U�T�ԇ��߳��`#��x&�7�AG�j��N'�[�j
�����<E� ���P�h>���������c�>R�B��;+�Y�W˱,��U<·0�����W 6c�Ã$2��P���y?���o>�"�bJ� s�!P8��M�Z�U=����`�<�]��
#~>|��}��'��v��kD�k�,D�jQ�Tj��Y���8θ��5�+�)�^-�R�I�bT9���k9\Lٕ�R���{#ͭJ_K %V8`�al���!�A�w�ޣ�]Rx~L2�}�v���ۀ�'A_�b�JS�����d*�Ě�����c<�?�}x4�Y�ɩ�=oI*xn����mB�5�$��Cd����� v�'�3����|A��^u@-S��
��3��K�$X��-���䧍�,���o{�V�=Z�Y��R����B����]TW�|,_��՜�S��4O�˵Iܼ��`�ؒ�w��&���iE2G�z�� �B�1��{-+8y���F[]��+;&DL�оf�`o�}*!@`
 ~�Y�F�֕�q^��%<���rc�zyN���2r�ѲɠL��W�:�zx~�Y���h��U!�
K8 �7`(�3A��Ѧ#�]��}�14�:���S�lk�+l�}5ϝI$O��Y�8�϶���5.<���珋�V	����1��4�.�>F#�c�'x����R�|1�̋z�@���:!�Pࡾ������y�����"��^#�\?��8K+��R3��Qmm���H���YP6��1m���>�e�tLV:� >,�vj��E� �ˮ:yy^��{,�L�y(̶~R�P��w6�b_GEAj�O{���Ѵ2��64�|R�Y�Bg��iM�-����|S�kJ�O�.����)kF'KC�'�F�[���8�����c�J`�lxz;��!M-��;0o�B��R�E9<�Ͱ�P����ݻ��mc��їC�\�K8��^�	���r� ��V��I�y��w��*��x/pch}� ^'���L�M�j����aU�!��@�R��(@1�~؉n�*3�J���Jn�0�ŁqXK�Iv�+h�̪�`ώ_d.�U�Y�I���L��K�٪�j$��W������i�,n&ET�];Nc��`2葝�J����P��w;ٍIoSnL���C,��У`R[�Z���nA���Г��LE/.��\�ҕn^���t�$ӛU2K�U��<��l}�^ݑ����Hqя
������.�F)�.@Q~��G�|X��%�1���r)R�P}S�E5��W����gW��~�-I5�d�mM���:�\���"B��v��0K���V�`4�T;���8scC�!�C����o�5�����<�R��o�ZxͽY��Dr�� Y@�M����g`ݔ�H���[�bd�>8b��>��;Ҷ��a ��c�Bv.7$��n��R�p���DG�Rm�2	zO�7&3���	���Z�-m�x�N6��.��}�;�v9���=������>����,��#�j<U�; yTQ0�'{�=7@~�������t��_��5�I�K� ��f8Ьs�(Ɉ#�k@��n��n��������GT��OҜ��nS�H�ez�I�f"�ei�ʜ��<X�]W���_>+�K�އ�dEvQ�Ó?�e��/�+��q����/ngp��E�p B�{���u M�k�wYG��%�p�*+M����	3d+{:�Ą��+0�ŉ�H���x�:L��� ����������4��f�"�F"z*X�v�)�>�k��X���	__Aٔ�E�4G�	��#�7���Z��� �������$�1���!y�践(V��B0G��8�&ja��Y<F(�@u�LK��'��x����3�/g�������-���3>릔�*�+����p��C�]h@Ù���:�1˲&D��ʣA��
������y�)�Vs��,�Ď����>0Θ�{i,��!�^$���ZK?ۆꆭ%&��ܞ��Z��&�*�X͠j�)�$�+E��+�.7������Oe�v��1�Y��#<��+�Z�E�b�4cӤ���3���>2~g���^�0l�)�� s�V��O}2������e�4������7UⷩC� ԩo�N�	�Ӏ�)����A��PI!���=�"���ǉ�VP��ں�|)�~͕P{n���^�G�*��yE��S�]R暮#��Ї�u�����Ɓ���w�Y0η�),;��6D����f�,�b��ĭ7�q�lnC����d��:�T�A:��� �%�x�W���M�ԐFˈr��"�:��+a.���W���}ga��V�A s��#�v�kA���h-Yl���wt���P�&��8�Y�#�:,O��Ej+w���ayt���'H��v��TD��Jgc��~ᥗA`�Ӝ�_o�}��1F�R�h>m�#dQv�k���/1�b
��"Z7 �l�:����� #�W�JE��V�uN���:2xu�q�����@>�d����Q�ZX܆�����&i�c�xô=�ޔ�����f����
�B�N��ᔭ0'	��bv�>�=��r,�׽�D[��{���>(%pɬ�����wy��l�(��i��
��QhOE�l��%�+��Kϼ���'p������V'��&�	�fw�EC�W�E�y�
��w�������ע7/-��������m�pK������ܒZ R��iU��*��;m9L���Ā�0.ݧ�RcR`�A���.�(�J�>��H����X�9cPRFr>�'��2�-S��!�c&��ՋF�ƣ��_�A� c@ [�F�ڂ�Hj/�HM��a+>f4��Ƌ��~���RQ�