��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|��We����P���\-�O]4U�bWy�T��ש�ڪ�a�:�D���*m�f +'�ڤ!���~YCW8vs�bS��ϻ1R��Q�P|1_����o1zJ�?�f�����X9e�W��ݦ<����	-0u���8��R��Yʂ��ZR�я���3�K;ε-�w�&�O���8Ǭ� 7h��Wb�Σ�ʺo�.�}��(%p�eb3�3/��3DTa�J�C���0� qǭ%��0w�](��QIw��N�o���rj�Yûl)��+�\�g�5��8��W�k�W�ѓCi�[Mi#�d\G�w���@s���-�9y<�����f�?�|���7Y:�Ëw���y���UA��n�~$����A���A���[�=��/�&$U�jǿ�e�s�x^�^��,��(�:'Py��� �����N7�G�k/V2\+bTm�@C}��߅g����
���i�J�1��Y��
2�y+�D��,�6 _�n��	#�n�1���̐�om ����M��@p�`�(ן�n�}É�>
`]1�!���A�xM�>�� ��kS�����6��U<�mO�F�52��o���Vᵀi��M7�l��ta�a鷂t����"ze�X�fP�e�����N��U�ɧ��5aX�;>�D��A��c9A���2Awv��3U%̇d,���-�!�k�.�������5�;?�&��6�q�a�`�H�,X��OO��}��컂��pO3�e>���΄�����]^(�_(1r��l.By�Gd�婵�R�gL���K5����w����#6_��z�X��v_����4�V�r?����ƘuK#���y�m���
���O8�}"�8���Eo��V'j�
�&^ƍ\��@����"�i�=�7_���ٙK��q�L��f.T �JQΓ��/b=�f�c�|s��X�mAW/�v)%��~��{ʭa }���^� �C��hߗg���I��S��"li}�`��@�㕺	f���Ԑt�,*�>�m�9N����>[2W2��Alߵ�v�`������r�4�F,���T+i	fm�E��Z��^�"ZU��ۦE���PL5V:�l�Kej���!���9�G���n] I����قӂW[&Tf_y�`!����n �3w`;״���E�Ǎ��eT.Z�q�]�����!�}�������9@#���� ����2�BX6�еa�+D+�Io�� ���z"B�Bg����o=�!=��kg')*��_yq#�� �R�z0n�LJ�V�2��w9|�)D�vCΌ��m{�K� ��p>��"LT>tT����,��e-g��3ø�/�� wuma�?�� �l�7k"���&�*�G8΢?�7�Cn��C�����jm^ۇ: �k��6�ro��WxT���,7��-�+0Z�9�皃˨K���n��#�#�-E�Q,+�3I�;.�.��y|T�y�	�vED�6���@�v�J�LF��w�������4\�i��h��2���;���졕��P��6�U {�R��y喝x�����'�[�^�ŃD�O	.3�t��
)JT��P�	��3���~g�<�yFR'K���C^��X���2�rg6_��	�Dĺ����u'�$�a_�p/�'���v�x]]v1�ќ�]>��~{T(o7�̢Iۿōj5w}�۴��%�y��G�eD��1�N\5yB�y�����0�L���W%�ͬ	�3�[�����j�(_�F� ��؉}�x�{�2��H��jC�7��L[�������ugf5)� 4�T'.z�ƾu�7�e�3�Ha�IB��p8O@�X�೸�eV��R��d?�<�QC�w_��{r1Q�<�`|���g�1�����L�h����Ý�kAd����y���S�.��tR6l�E������i��.�,�:�:��B�-�|~�EV��rAb��GBR���`����Xj�mۧ
���7��p����u`���£�h�rد2p�O)?�$'m[�
cǧ�{�Q��)>;��?	�?�f��Zf�²��$`�pN����'v;�"�^N�C�Ή+x���[bvs�:�~1e�!H�ǭ��nt�.�v���L�D%*8f��\0	%�h�r���JY{X|��w3�+ҝ��|�/�	�95�Z[w�k��Ä�;GC���&�zV����#*������;X�y���TlwB��5s�ϜұJyH�ǂ_(a�{�cRͻ��*�pWP��M�X@�2��)�O��]�|R"� |)���>x�oč���
�:�2�zV�}hw)r�{{��bc1K�jL����-��۝Me�A�&�����+AG��*)�R�Q%�E�FwG��Rz���;�a&����Ԟ7KN��9:;��6-��Q������o����Ey�bi�1�`B*�[&z�� -݈��p���#�Ϻ��e,i����r�mW��V�|��S�2�+�т��cCPՌ\Ĵv>C�1��:|c�f;��j]G�E��Ɏ�k�!��Uov���e�`w��3��X~�������rħeW$� ��|%��ᚖ N���'"W���1�n4����c[��5�
)r?�5�[�0lx�9#�n)�!f�6QhI�%K �6����#|�)Ҭj�Fpߛ�Qs��� :U�Ӝ%T���sN2��7�a=�t��_�L�%�ߙ��K6�O���)�V�k�Z+/����e��ϧ��857T�(�h�ŋ+���'���3��Iھ��τT�����#N��2OO��=�:�:ZEX23\˔՗���u1E+���l
߲�b+��Z���9.oDͤ�Sj��`(��>U����C_5��q��;������򊘐��5����~�L�Sc^�3�OV�%��1]�2����QZj�V���f�Xr,��N��g���ԑ��x��]��ɣ���$��&�*�,!��5�c��z/�������6=0[d������P��sl�B;������k�tsܘ��/�]6�KL/\Au����~A�К�Tl���ǧ��f��l㚹��6`���^�~	��d�C;Tk���)�JA�^�̈����K�>�������bDG&�֌OQ�=bP,AF��w��L#j�vV��,t/p	�	
e6Ŵ�����6"@��.��L���L�*�`�$c��X��]@����uع(�]%n[�j 	M�p�^J��9A~6L�V�D��ՙ��6�s�dB}E��O�M:��%M#� ���ӂ�=!�4#�����(�s�	�p<�Av��jyb�y:=P�<���#"�S�Z���'D?����*�V%`4�M� �D�Szz���X5/��jo�v��rT���t x�=��-�p�sݦf��I�z,�G�.�t��Dn7��Ӕ�nyN��|݆g��$��w��+���Ys0������cNJQ�?�U��/}PB!"�M^��*8 ?���f�0���_�� Nl�"�02���\�'�.�qR��ܳ��[L3M�=׫�--��-�W(�9^��U��� MFUe,*�rK�SL�$q�i䴣���uwM�1��k����d���GK�$I1�,rS{r���%����OO���d��ㅬI,!�?�򷌼O$x��cNn�|ZI� ϼ#.Ğ$!�u�rݖ+��1�h��	;��k%+9�����gz�=���֓i
|_86ܝ��g������a'A��.�L}l	���IP/��K�02[�^�T#ry}ݕp�\C·����P��<21�I|��F�e�O�fu�db�'�9J����"�V��y�a��e#��y�wf��2߂'v��Aj�W?"��:	a,A�0�Or����Oڤ#~!���g�n.�F�^��P?*��A���:���^�5dƫk{ؚ.a����:�K�����1M������r	2�V�U�t]+��|��E=��-·U% ��3˸�,��cS3yEM��+�/@��9YC&�pZ����ku�y�0�44�,�d|ό���|||0�ĵ�y7b�A�T�0,���ߣa65+Ҥy�y�?�VKc{�o��m�xU>��w�E��Rk���E��n��i&I��3E?$�Z/��R0��kI[�M�l%�O^3�Ԥu�iF�k�Mk+j��"4�Go�SG���1��nh���|�W����� �����zv^>&��������CM�����< =<HN3)���n���L�dl�!Pu��ƱU%ͣN|�0��_m��pKd&���K�b��*1��*uFV��;��uw^�xa���]Y��#�; ��׻9z�#���s˚���jЪ��3U�Xt�Rњ*B��K|4[k'�hR�ez��y7^g��-���S�����y(�x+h�yc�+��"�}��"�fa,r"�.a�bc�ˏr9�%�N�]�#c;��I���}��j?	���Yq�9���{-ѲiK�CPB���'h谮��	�9h��O�ef�Ѓ)�1�p&�Eٌh�Q=���G"��^��JI�]�h���i��y���֚�_��_��-v���h��_�LdJN�$��?���.�e7mU��2ǧ���k�V���k$�kY*j$ғ�V�\"�R�T�ZƧ�,���a��g��F�z*�B�P�l�����g�\T����kU�&��$��kȏbDQ��(�]�G���:�:ܶ�ri�3�f�ÀH��
��6\�*����L�f����ʩh 乀��`����̕o3��8����!֮8��+9C�T=�?g*���+=3���aD�$Y��d�DB~�-��KEؗ�8Ulj��l��о�������X[X�*�PЌ��1Io��/E���>�~�G�wL7��InȐ��
K�b�m���=G���xy���(>�����^=��V����&�g�lߘۆ��)��dp{���7��	�vu�%�Q.��G叮�O���b���!z	ō0�м2AwS�J ��I��P���j�F1 աk߿�щ�?-e�k'�������oS�y-&bmQ�ox�H�R1˝�:U`X��Ժw��2�$oBj��j��?Q~e	q<=�>�����t\،��< ��m{���%z�rx��F�H�G��Ҫ˩^��wb@�}���~i�xG��`"F����!b��0e�WhL��*�o?�?i�8��+މ�}�b1�4�rai2��S'!��a�ʋ�o�T��큈��V���j�m��V����ӜO�<E�=헊�! F=M��菅S]�X �.����Y��uݚF�̹��F�W�U"o���Y��}$���dJ~�*���� !r��/�f�+R��t��s�6�J��`穃ǉ ��8�1ֹ���|E�[e�J�A~�
�cs>���)�#`,2�ҿ/�Ů�T8�v�T�V(����Ph���DSmF�����u��c�h�7
�b�ƅn����+k2�oVQ�,�^�O���%TS Ի����j`^=+��u��~Q%Y��Z�5�ͥ�Ge,����n�ü��I�	$B^����	E`.�{��������ȣ�W�,�c���M%&��Bv��M��wh/W���M亂A\y]s,g���Q�It�"��B�Zo#���dKri`L�!�mM��"r«%�p�Y@�8y)��������Q���,�����`m� v�Ib#�B��cs�P	+"^�uF��5�MK��*�8`���C�2���N4�<����#�=cT� ��D%�0�|�Q$͈��:�D"���zF��}�^��ֶ�D�>������c�K���jϥ���ߥ曜����OG<��d���	��[oA��}f��5��Hn���o���_Rƭs7��Q�JHH4R�9�8���,̦tf�Je��;XO�s���P�L���'Z/7s0����A�;���}Lv�)d{�Eʿ΃�ȓ�g!��+2j�����D��H/�Ul�V�Sx��=���� ���{Ze��������95{�3�5V�`�J���pL����!e�Q�Py��Q�fg���v30x�^]���-��	QxF��&�.��3�ۛ��:�񁜂5�_$D��F6}v����<���HaSܥ�>5*�\`����	x-I��v�;���]P�,|(�^G,2F����jry�vJV��F{I �~3��;�_q�t���̑qU�������2 �t�-����T�һƙ4��\"1��v�J�ߣ���%�6#p�H��f*�ғ���p�R�e���&�Zh`e�4L�o�����K��U܉�Iޘ{_�$�Qo_'؉�6���̄�*G�]���0�qF��βK���zn�3��=�؎�v�ʁ����ҙ�q�Nf�o�]>�G5Gr���fhX�=�xzM[פWjʼ�A�n~CO�J`�˕��dG�~�!ew��F�1�Zct���{���2�a��%��a�r����@@��k#yB[)M��<�~Bմ, ?I�C���F��r�������Yy�V~�L��7t����g���cīV4O�]r�ʫ� V�h֞t���BVh�Ȧ�&�	ԅe��(��]6�H��߁ƥ���jC#ܦ�8�5t�9���޺HPL���HmY� һ�!f3�˰8�F,2vWU��b���� q�=�:$l��]��vt������d~w��Q_҈a�dq�[-�e�O�ǣ���爽����1ܻS'��|��7�L̫ui��IS��O�*����]��uN��(t��<��Rj^DJ`u�
����aB��M�[�T��>�v��$ؿD��Q9e���C�*�a@d!<���y���+r&�3O�B���=���'��� �h���ڃ���aFz�
U���p������X���7˚}`%߳5+AR���%'�Y�CRoN��Ոi�����R��!�����:Od+[��u���!���?��[�t}9�>�1}��O�gX��6���)���>rO�}�����M�i9�?%%T�*�p8�gc��;��U3L*����38-Ē(5�����������ٔ�麍�.˔.�OO9KB���.�����z�<�_��G	p�
�n� �w����6�[r}�}�Q�O�z_�%�a�MX�����dl��`�ܺi3��_$߰�=8'ǐYf� �u�\�I���Xx�M[��nS?ĺdx��?T��f[�[q���)��[P�\ZD���b����=^�
�u��OרSX����������gnM$�N.b��:�'M~x*p0�˔�f񮴞Q��0��'�P�cU�/Bu(���D1�>�r�E�LVq;����^�D�-	{�����k��&��]g7{�&]y9��؏}��=�G�+=��hj�0c)m0�~�������;�lW�I���/��q���>ޅ�iW;Q����R�7�h $ޝ��`z�"��(��c���M�փ��+0c�1���Na!�ڄ=�����O�����U(?�a0���v�U*0�8�k�@EU2�'^e@��
+ι�/ ��gg\�:x�Fc͞P׹�����.b�!T�z�_��G'��jl>hKT����E�-kX��\�i�D���X��_�|�+]y��n��X���m�t���K\�F��f��~Z�8J���4����=0{�խ9����HT��MJ2b��Jdn]�s�,Ԃn!�1���ɒ%L�L�K���U�e5ExJ�hH�-M
,8�*x�9>�dm�ҋ����� r���8�=�� ��n�o]xn��k{�ʜ��ya��-�N޵1oP�$� ê������>=����p�1^+��b�w�Ҁ��t��ZF�d�R��˙~E��9��s��q�A�ǶogYY����g�7,�?pz�P����hӫU"5݀�15@��YS~��Rʣ[���S��2����(�H(36Q�h�g>��^�@ {o�	E���٥�K�V��o�X���@��o�{N�������;EW��+���k�����um�*�:�u:{��']s)�p(�WFԏ��J���KEx�� ��y7ԊLբ�}����O����<����>�t����yOF� %E�D���6`��d��@�cB}J�}_���bd��˿����>iC�+���/K�}G�]υ��:uE�G_�;ոL��3ni�Ӎ�;��`R0��#�r�dHcΞH���J�M �$���4#����Lh��ܲt�ߡ��џ����a� a�ܸ�P��I���[����hb�(�3��v�D�{�<��|�p%��hZ�Ŵ�GGu����|�R� �vOP?� !��&�ot�KȠ������@jk��P��-A僶ɫv�x�p̦�ܿ�\�Z�!�FV�ZJ�)TR�s��r����)������q��eu�=��&9dbNغV�H��kB�g>�C�=Ϡ�S6������ގ&��Lm�5���4��`'�2m�!�����ly�*��L�BU�J�	^@����_��}�t�1#f����,k �3�k2>��U�CM̓+5Ӡ{'@��e�m�����D����C�{yB��)���7t�(1�	�B�.%0iP-�6��D.�&���j�p�W��'��k�hxks;�cY�� �T�-EL�����L�i�_��l�M�q_��e�;����:H榘�-0��i#�9���۳���c������b`V�&q�u:�?��)C�V�/bڴys��HF���;*�@�?�$����æ�n������`�Ӱ��m���&:v�7�R Å�~�c��r�X6���z<lB���R*�0���`^���Q9�����zN��զ<V5�M]E2>,_ {�d����	�Q�=��;����c֤�5ē�T0��>���(���"y�iB��e�ٳ۶��D�U�|�P�Ն3I^��F_�ᮅ�tF��)m;�sL����nA��+-���׎ά�au��ۙ���iV��Ⱥ1o��c~�A��\c����=��{��!�l�Mt["1@��C����4���L��A�օf��+B�L��+$i��o�
E"�PV�u���QD�G�=�&*(9�ʨ�p���=�q��3�Nj�s���]���F��R}6�ջ�ΐEF���i�n��G)�9��)P����Ԓ^z!�f�U���u+w�g�	���&y,�؉���M��"d"�z<�u<�:�C��e?/J��6X���yi�#ϥu�,z����>h�;U�6���U.��x�<P�������z�e��q�SN�R6m�aCɲ� ��� �Ʈ��ʀ��R]Ph�����$v��W|���[���vu/!�@�C���p��Ww��@��e�����{��L�q΅|Ww���kh�����`��?��$z\��~@Σ�'���m���14�D��2|��?:�+�w�<��(#zu��lQ������9dl�PԷlgY��W�t˞C~�Z{�a+�j�-h���F�fbD�!uZ	�Y5���a��a,������sp�G�[tn�A�+f�4��d�����U���?����8r�`��	=Khq�Hj[_�r&D~�qҚ�� z�M:�$ERG�Q�.��e�.EU+�R����jV�_�(ϋhI��ݾ�YR��/���g�6���ѫ}�9F����6W*!��o+l�Lمr��v�|���SKD��֊�`��w#�#��$ĵ����p��M/пv����I���l��Ppw�4kj!�	N�g8���#^a͠�;t�C�YB$��W.��$����4 }by�5A^�'���zW~�e���0�d��}EÖ`�6�@g[�֊5��9�']���Æ�o�~���o���l�pj_Ű �j���dN~v��S`�
4�Z!��572c��N�(����,��sR���]UWU|����:+.�5�C�ߝ���?Hiħ�6_̅ߏ��Jb�rƒ�./�/M
�w�h"&�����];�����v���p��(��jL3ĥ��$
����wnY�N�Q�0hA�6��y���/�}�CAU#��Q+�Z�;��]�9l�_�;RC�P�x��*�"����ːۅ�����W��D`B��j;��e�̣�k�.����X�Bo�L=Pz��o>qj��y�Z"��k.�����>����YV�y��(A"�>��CO�g��٦Ke�J#W��l.� �����P����E�a�G�{�%����Z�|:w_���\v�|�s
'�5#�T�p�1pw���"bJ%�f��Eq�ۂ=M�uXQ�U�Q�N��:�����1�1�k�rve2����Sۙ|`RZΖi,	�D�����s�$Ʌ5�l�h�I"�x�� �(b<&��yx��8��+>��'����hߟ����ݱ�����$����k��!�7� Q�U��ɧ�.��+hâ�S�����"�g�뫷�?�a��n���ֻ��8E����Bs*5�h����u����^��{�uoV�>@�d��YM-9����N,�����1T�,�I\��0?�gܳ����+�"𩈁DP_�� ��v���8�?gFn������xo3�/��]|��yU鞔�f�2���4�)�2�
'�P�.0z�t
T�+��s�XV���2H>�I������ີ��.�	I*�.n�:�X���g�]vYbK�H�iL�S��G�=f�~E������Z�L0[}��)q_�uÎ�Ͻ����."5b�ΰ��16I3��M����ģϴ���!B�2f��3b�&�ߤL�����\#r��sj����f�.�9=���5)�p�S���I�*[��'�}�O:������xgA�9����[eq�-iHݷæ9ׂ��sMĽJ�T�O�m��3;N��GM�9� ��Vy������U&+�(8,��:TL�箅A���K/�u�jEn8�X�ʕx-�R�p[F�Z|�\�����H.�?G���1qJ� ��O��k�9	~�y�	G���p��m5 CY�����R��u���N��P��t7��b��9�1g�����g��8�%"���$O|