��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|ۧ[����&I-�M0MFɵ��za��wC"���6%З�ޭ���ɭ�&�5�D9M�@f3�� �m��1ft"�u3�j�T�������t�E_�h�e_���`z��28�����[pC=�~��b돖$W����<��a�u�W4�(*�.x��4�t8)}��JF�����J��>��G��y��Qy����C�:7^S9�aP=���m��{LּEߣ6��	�+Q��^�e���'�����g��t\�B+$���݈M��B(�:u�A1��m*eY 5�0;~��v`116��*]����n����������[LM�b�H���;�h�Ѯ�
ȁA�QXd�Q��C��r�8&�8���u�K�k�07���O���c���)t��^�$l3�e��ɲ���U�>gJkXE��H�5�R�Ƅ4�g�<HV+�����1��]lVd����?������hs�`}��#���N�s�Gc��F>w%j�l��T=
�y��K�pC�ŦO�TO%V��ԧB��G1
�u�jɲb�)S�ݷ%�:h��Yc�/A��P(�ǆ��n�Y�{�N�)����l�h�i~J`����@�W�HA��^F�q����Z����bPB�
�QGWu�y�\��T�M���z�99��n����W\��9��FA�;-��ᖣE�J������	�h����N�[	,ާ1��gaj]�]�.jh��3}�w�S�)/�=��D��y,f�+9��l_���%� �]mH�░���������c��')�����&�ן����$���uA^^�7�`�
m�~�f�Th���VD#&#4+��dAA�s�s�[,c�m�q�b�t�� �'����%ԡ{%S�Q��.�;�=c]d��Ӈ������e�>����^�x������P"��ĪKj[6KYU�]K�[�[4�BqM.�l�b� ��R*o�����D�r:3֯p�xO+c���G�|���n�Vy��*m���#���ǿ�FL�i�!ĵ�	#"\72���8���-�X�z7r����*�EO߿(C���}w��&���>�ޅ��r� νb�d���ؠ�`�G}� ��?����
&�Ʋ��5�Bx2��s�����R���9H����V�̻�z-�dp��:���'մ��ՏX-�*����pP*�5���_]�^�L�M�T�D���!\"C�`��%i�e*��NwvT���.�P#�vٻ�YtӀ��"~�#��~�7-~�Z�=�N����d61!�߭EXTOhn��)w��;�t�����L/�2q	��~�����9L�a;<I1��V��v��5�y;c���S7�tg߸���!�w��a�Ͻ��,�Q����qz�0���7�l�hH�U�"����v%(�}�Ayi�~��Ra8���3��uG��"�w+d����a�@�r�(��yBJ������f_�4�Dy�e����������.Kiڰa(.���0���`B�% B0�d��������'��U����S�{6T��l�4�ɀ�ط�{���$�;���j�V'�3�v�:E���6r�q�W���dugy�,�}�NCd� J�HgV�]�K��/��CN	���*�|��^!���o]����r!Z�ӢI�oOCŋ��?bcɳ�W~~s��{�\
�\P7�Uy��$�U����R���\�,�{D�x͸ty7H��%N�Z�/����n9�Wx���r�mQ+�3�����ج�#هF��������������������^N����q�M�	jqA*QO5���>�6/Ny���v^����(��e�?gk�Ny@�G�'r� ����_��A,�sX3=��`x��e7�y��J�_��!(g���ٟϊV�"d������m�N�h��*�2l��V]��.Zd���J�!��܀�7���EXʇ�}����]�i�l�B$�z�*��7]��gM�&�~�^���((Z���c~��7ɪ"�+3R$���(�r]h���|VkM�E�!�4��h�L^IB�9O|�7�ff�Hܬ�3-ߙ��r�&��]XgL�$b�S 	w�뱹qi��h�`��8h$>����`-��v�ً����Z�M��r-5�7�J�50>���g7j�wS`���e{-�cإ+��rb+�x#�˾.�X�>4HX[�r[�ڒ�"w��p!�կ	_pӻ~Fe��G�A;W�������1�{O�Z�6?jw�ȟ�t��M��=�^����e�6Ic��+��i��.���O�E>�	~�	���<�	�FM�O��i�~f�jr�O����-�����V��72��
	y���q!m���(Z<uM�L�bk2�2�� ��� X��8�`I#��䰾}�#?�6�k�z�^�C�#Z�	d��Z��@��.�H)�̝yj���-2�g�9o�0v��pz��ũz�ia?�i����!q��	�5���ʻ����ٷ�u��	=+	����f����
���ކ�Ek�����?=���W��[�����ظ+ڠ>��Q�f����z9w}ލ�m��?A���**H�2��ԫT�I�t�'g&Z�>�`~���`�ho�ʴw�a����-"/s�%]X/����ђ-�S�q�~��%*��[�C 4�h3d�>:���qS���cu�6��O^JT����������A��V]����l��5�`Eζ��W�b�4,��U&�4|�z������=����^�I/K��G�+�R��-�A��k�Sd�fis!��V_�����~Bb$��˴_��/I�g�Xt,�{��03��L�H�������-������<J�z��++���2H֎'唴m8���@�K�6`	0Oe*�F=���
����i���jN�KG�$�����0�v u�q�&P��rqi�g��D���U�&5�FcG�N�_�>�X,��F��#z��v��<�Ku�0ֲ�a[Sp,׷ �!_�z��l)U�Y��z����#�<-���_���g7�7v�/�ۆ�i��Ǩ,P;^�up8_�[b2�kɾ���>�2�Q0�s.�.�C?�XM�#�7���c�e����F�5�j����@nNu�G�YHZ�Wf�24�1��F��~�_�����h��O�F��������h���{5z���58
����o �`��=-�A��Cɹ(��Xc6%G�@�ZY�-���/?�c��3O�l���:W~Lz����r=`э~�[{w��3VH��m8�����j4�)QbC&���Q]W����qx6�H�٨��~C�Ds�w|)�|�<�;v6m��;`|���T%�b<��	�=W��z���H/U���Wů7�@��Jн�/�Ӫ<q !\qdӷ?��8>o��J)����Ճ�i>��������zv����?����m�C�I�/��#�*ϧ��m�F�~eg��9uL���}h�o�}n+��Η��u
����op+��-_�0�F~�Dz��u�*�M{��<'�K�e�uD�����<���PlFB7��IS�U�7λz���D�+=�����~�i�<����
}o[�{�EX�YR$BY�R��o������ <c��oG�r�T�*����Ol˿��#�
&������K�J��gN�#���Ę]�4Ѷe)���sư� ������90~�lt;����,:u�E�əx0���*;%����W�|vb�w<�YzR�,���LIE(�n2� П����A�;�j�����šO �u�l�q���UJC��G��� �|����/�M�蘖B�~�0
/?�����A��hX���֜��	�j�}��Z�(�M>��"�Q�<���`t�D0"l<���L���Oخ�4�_�]ҍ�碂]�ʁ��}��BǁI���R���p�\�������[�?�[aiV�C��>IڄHs��������$�6ǂl�/�Q��f�Ja���z�N���nH!��6��cO�4u�	�����Y�4Ή{�v݈����W��8���wrjnј�� wS��;��~ؕv�|h��zIX��F�#�Q��jBuQi�8\������Vw5w5�:�zPPjU�Ǩ���d+����L��!��6���킃'�i���ǽ������Eu� �S��ߤ Bws��������{��?:�p����(�kyn�g�fԬ?>8%U#ot�!��E�~��}g�mb�<̟�Hgސ���i����IZ��;��I�v�*�),��(L�!�Zb�˄ZI�}?�m^�莡7~�V;�sy(�j�a��S[XO�;Pi>�o��H�o奈���x<4u�3��=iad�U"��8;\K6�Q�3Y���c���Hd1���&�YLo������ǦnW�No9&DXHg�\%ݦ_��hL'7+��B$����S�ˠ�8%�r��d��B?��@��&��8�SUi2st549��L^W�=g�s�VCm��A��!�cArM� zn�C�����0�[u ��׺�v>m�|����1W��r�f��4��K�Hw�	�c�$)Ƞ���ל�a;\HaO�9`���n���1u sMBB�B���͝��$��T��H���t$x�Wk��2�8�h͡O[��Jd�aib �I�0h�p��o�����d��_e�b9l����	��[H��N��ſ���Xj���FL<��e���$��~eZ�9x���"�z��	Z��$�
)��m㋾��"�tGg�F�����(��V�v֔6'_��hg޼�5�5g`T+� �-�kR�n�T����A'��_P�Z��"j�=֍$��BUOվR"�QH��c�*fc^��Z�f��g)��J����iů�k�/W.�m$���=+K�/���xM���ٻs<AA]_�9F� �͟�oF~�c�~@-�����H:�}��]g;� P�u�/��vŮXn�$�K�p�M�O�c�HypC�	��� ���������H	�\�~cT ���J���ͷ؍�Q��#i�ߗx��n��1�LB�3�i�[H��=���p �������h��m9u7z�&�w������E�C4�ę���{���v|�*�&D�8@ʑjq�AC:ʹp��P���+ �b����T'Dq+͈��W0slXN -; �-�@#mH:{�eS�������R�zx,B��FJ?��v-vj(YN��K|+�' ��M���YHl�D k��G�^�O�?ϕ���}<WS`�7L �e�Zt|��4 p������H��N��|5Ϛ��d�B���GuY��)Z�q��+GC�잌~��p�o�p.i��]�ar��D*�zy�,�����p28�a��X�B���;�/�#Q)��]�N�|��B3����/Yp"�iAI��pD<�O�fP�03K}�(vٲ��E(���p�ʞSU'��~4�!�����t�+��4��<�o������Sk/�T[)Bl5��N=�
��uK�F��I�>��1��_�l�+E� ��ԅ��<&n����ƈ��%_�ۼ�=�3h���n
�"�i;�BGV�ui:�&p�&4�*��Jh�JA�?�7�G���j�WP�h�e�g�#�k��A�Ѧ_0��
�_m�����n����A��zB�8�U
��\?�d��l����R�3�S����ȣ.�un��EҜ�57������`�T�v�{�q]p~E��F�F�ڵ�N�b� ����Ǩ��;��0y�6�
BK@j�r��?���i��OC <��/���G,oNE/������z����A2:\� # Hp0��Kf�y���{@_���'*p�*���3F�/�����e�ET4�i�s?�A�����&o�'����f*=��H�PZ3�n���I�C"�!����c��S���#58K;����5����xX�oe4
���qA�[�aJQ���΂����#P�"�W������G�p	
5�X;O������G囲�r��C��2���;D�h����������l�"a1W� �k��*�އg��_��f��XF{^���g>��փǘ7/Lv�1�	�����g`.���O��pR�j�X���<s�֡�ʵ]\RH��A��ʷ���N¸`�A,=$�3v`�Md#�f��h���2*��+2`a<�oV������wQ��;cT�3�^�j,}��q%���ªu�q&�l� �M;W~�4�K_7O9+|�i�_ԝ�R۪ W�:p%qj�w+0o~��Pk#l沙�$��IL`�Y��+�Vy ��Gz1��Ӿ�sm>#̛B_)$a���� ��$��N����r%}L3/JL��w(6��Ԁ&'3,J��2cф�-����0(�Y��)�bw7�2�Z�᱅�G��#�[B-�FD�q|�btL��j��� -��j0:,�ʷ���Ў���c�?s��AO�U�F�v�={��{5���������(�h"�c+�r�¦-�rY� ��ͻT(�9�z��0X����Nj ����|6���z��TC5$~�U�={�9���xHӟOs<���>Ǯ�&L����bǏ�C�:���c�%�B�Mz//+_�^���g٫��^x�bo�3�m.�:�c���;ԡ1�U^`\v�I�¡�[`�|�CnT�'�E1�'qB�;z����pH�+�aI�g�-Hf�]��}.V��_�x8Y�y�V|���%��i�F�$��Ě�.Q�wJ�0�*dop�^0n=�j,j�nRKѨ<3j|�(�w��TN#�d�z���0�A����gI��ae��U����^�{���{-:�ݪ�534�7̲�S��1�g��/L�=!d����'�!]�Hw�"��hW(�c�T�X\[���}y�7����w����ѽU��A��T��DP��Z٢�h
�8�2'�q���XK���@mN�uXE�.
�M�}����B�:6�J[�'�(���\zͦ���s�i��rsN���I��NB��^��NԎ����(��L��r����]=T"��w7�����Ш$�w��[�z�}�] ��a��l��x�̀���g������L5H{l����r.O�݅@{w`kiu�zz3��Ɠ9}Kf�HԻ?E���z"l����!�,�W�F�
��ƅ�"��I=+�3��7�H�}���8QRGN��!EW����[����q�;�m3���#��0~腏�sW��lpc4�:��nA�ee �����K��<�ý)�8z`�_�\P�[@��А�.�V%�g[�wI�	����X���/�I-�`, �=����5m!{B!�\[��U�F�1�W�?�]��(�|�.�9~H3J�!��9��,,�-�U1�y4���+�H�i�@;0�&�8��ߏ�Y
-mY�m��,��ql|�_X[�����YU���K�f����R�(�s,e��Br�(��]�#�iagµ�`��s�Qik��#�g��a7_Jw��ˬ����aC�n[(0w�'7�G!K���	"��A@��T�R��}M���K5�>?7�=V󿶫b�u0�
��'��Ev]�c�E6R�+�J�.D�Q���y'�Cu0]�����������{���*mN��"mپ�p�ZjR�u��B���z����I�x��;�v�_��:�]� �3�����jVt�p�*$�H��q��)��ԃ�����x��p˰�E�@_���$w���hט����"x�(�8�X	����Ё���(��i<��n�������Xi�l����F��eNC6��R�c��y�9j�D�A({ҳ0E)�M����i��`Wb�Z斞Ji�&�y!�5��6�ׯ[��ǌ��
�pA�:�`���{�p�u�.��q�Sԛgb$k�	�~o��A�W)���]�lA5�菻��a���.v{`�����$2Ϫ�W�O�[;j*[\Z�{X?�����\��ʚ]�D,k�hZ	��Ҏ87��r-E*�x=VX:&�s��6�	�#�Cp�*�Q���?ͼ�>0���l��L j��R&�@��%�E��\ʙ�1�.�X�4�U����T��]k�vqψ��g��롵:
3[3i|5�V�$s7%�5�=���1 ���4�(�~��Ѱ����S�L,_̼oC�B77FV�^FU��J�k�q����� �\��W����iǩz��3` &� �z�6��ݷ�ề�:�#�̙�}�px���W���1ܚ�4����W�t��UG���ǃ[�^k�gv���͑�v���z��7�M� rtz�X˙@$�HG�������Oa}j��t'�����+O���Eic�B��פ� ��C�5%�	ڛd���A�p�rz�	�L�k��o-@����ã�ա��l��3zhdz~�0{:j�"��,���)2�"�/�`�gE�(*��C�
#�6�_�ݲ^��.Wd{d�5m�]!g�=�+��cH�[�m*P:i���������Y%
:'�A�yÛ`^kW-3Y�N~��Ș�L[�c�ˍ=%�Se�ֆ��&,�No�q;}���z�܏�~� ���u�4���(%8�����2��Y���r�˜`3)��>nAY*��)A)X�1"�����S�MS3��b�2���岪�V6[G�k�V[j�I�4������K��T���q��V����+��b\��W�E���	,�'��?�����xneB��bŏ`ۉr�a���}���'��+�ްY�n`� �+�Bϳ����
Z�:���Ψ*Հ%�e���3md�%H_sRZ����)9�I\x),��[hA�7��]�k��}6D�ᵋY{<�dƷ܁�Ṏ0w\C.[I�"�4,Q��6&J��ം�C����-c
���k�P'�Q���%~	e辯3���!\-3w.�\�Y^G�KNb�?U�A��ۀh������ǜ|GR$@g��๬��I�&�;�.��aZD�%�s����g}/6/�k^\�ˍ-ߌڝs���}n���-���-l�#h[{1F�9��S����N�B��8B�P5?Wu=N
D ������g�8��vK͋;��([VrT��i�b���wp*V�%�V> ���ϓ3�,5ҥ|��^,�$$jݜ�����&��q�؁cV�"�8�]F�B�<.R�|ϋ���5\�Mh�3�C����b�p�^�mP��c8H�ANK��τV+%��S��0Wx\��4$�S��L����3�׋��*��Į�������V��2��l9��l_���ŀ������-#��Z�g<�H>�� ���%���*~W�p�Q |��D���������"���ǅk�<R�
�����3��_��{6�
������|u�<�2k�Ϫد��=�p�Ina���K#vB.��>����"N����0�l��A]���4p��pEn��sX���uj�t8Zx�G,��R �F��ڠ�!x6��UKy���UA��<p-���I��n�t�Mҫ��%Wp�(��ol�'3��|8�P~3R|]u��K��0L�({���d�+����S:V��p>�O�-(0%?mU6YJoVMX�%�&���w�L�Z>7�';a�j����1�{PIq��]�
C�95��y�n�ۑ���}3�D9,��X7j����ᖠ%~*<�z�T*<�mF�|�0�����{P'��®���3��y��c��D�\�s.�xJ=��9s��«zؘ�����#�[�ޣ3�CPN}��HV���|f��\W�jα �mLx:E��r]	.d�K�U|��*+�̌��>��=��b
���Y4-N�Ac��i��t���(4�o-��	LSy�
_���d����?t$�1\�Qj;�^�� X�Mw��)�t(�Kn�lcs���8$���3$�ÉS׏T�W����)Q9�d����[P]6s�y�!Re�@ҋ5�%V���m����O�E5����������ܮ�0s���-�vJ��߳�����,�L�=�­�ER*�`�������lD
����ԭ�^?�nʶr�7$�"��!~�HO��mZ<fO���Xr�*�(�:�m��R�';��TV��<E��T��>˓<�̑�=���+�[�<$�y��˘���r�=ZnC��]�GZ�A}��L܍ϼ/�-���������o����S�~��s����2l�Y�e*���8�G5��=�Y���p�PI+Q�<P�N��3�j�;m��Q�:�v�9�����{����#��?i9��ˇ���MNN=�~wxN��`<9^�*A�^�7u}Aʥ-F������X��,L&@[���������Ѐ��ht{��N��]��Qg�Xk���|iX�8��g���|?;�?D�li%�>�6	Ni��:���@.9'���6��b�-w��ߔ�uVW�#��"B�+��`4���JW]i~Ě��_��q���@Јl7(9���(��6E�~�����5|�F�a]��������@��UX�PJ�w]v^���:��-X"ޣ�\kj]�}>��M� ���LL�I�cɽ{� ;��0�uUO%��ڢ��D�\\�&"�_	�`(�i콷��C/�1�:-?`G�+C��W�P��uq�)Hl6�^��t��������c�{rͳ�����<��P�}��x���X�/��L�����&�Oyp�r}���~<�Xk�9G�W�8;�J��"ݟT�Y�ΞH{�j�����M����Ȕ�o��5Ƈȉ���0&7`�ztm��r݉r����KG ��ſ��޳��ߨ�c�\�bȖ	nP��h�̓�4h'�v�By9�L8��s����o��bN{NN>�=�����CR� ]�2
�}5�Z)� r	��7�ŕ���G+�Sw�@�>��~�!������*2�[���c�X\�h�"�t��v�8�i��K[�L;MX������o������_�������s�J,u-1g&u�]{�; �=B���j�`Y�1ێVRx�A�Uk}��Pm�D�[:4<h���$f`�*eE�K��JO�*�XB*#���,"�t�O5�o�M*�T&ĿtE���N��T��>6�%H�fQ�h�-ɐ���L����R�8�}�Os�]R.��+5r�E�fya[����n��Ү���8��� ����d��Ws�G�\O�jT�x[��-p�;���%�ߑ|Z�m&�\�Vp8�eZ-*I��,m-@�+�+UHbǰ]�K�2"����ۊ�;K_[-��i���r<��xP�n40����~-s��#���p)��s+ ��x��B���ּ2��hɃl����g�+�J� �;�<IQ�:z-�BX��Q��T����\>,�.L�	���"w��>�I��K�{���a��7k�BMug_�w�X�kK^�����`�����/�e�+�[P65��~R��K� ���~�q�%+�m���ZSt61��{92��p�Y�������ؼGU��4�n�ٯժA�k(Ey��lZ>6	ZY��N$ L4��;��
�x�����SC��S��X��[k+���ĚT��s�-�K�`!�y��H�UA̺���[���Ա��^2И�"�P@I��&���'���w�� i��;N���$2P�$У^��B�j������z�&VM�=��Z�4�	�g��5�$��Zu����k��ɦ��k����z����бŘ$�p㾲�'4�P@w���8GOI`����7��m�7�8V��ϑo�")7���S7o4�V+	d���h7��X��.]�I���&��T��l�g��c�Tds��֞B�]�	D��$����=��aKTЯ��W�S|�_$9�A�������*}е��[6usF 9�JJ��+���9o\���n�5����=~G�`zB7�D�z5M���x���!J�А(�}[?�?&P�9"��t����ܜ_�D
-�d���nca����4V�尶;3���!W�{�:X�'��AAi�C�U��.ADXSX�y�NG���t�r&��^���?�����Id��ߨ�kF��a7:�T(�z��6�W#��v_1ʦt�[� V�5�P��b#j���	:�Oc�5�sQJ��}��ދVD��['��{�3%��U�<A`ݦ�M�p5�e7e�Eй>���Cۖ�pxW�	��"�[00������ϋ��:`N��N���i�������s Jv!�]�\�p�'Mv�31��BlR���;pzQ�Ɋ����[�_ٹ�߹�6�E�lDnz�(��7�z/�M;<���&.X�kd�c��!�/S���KI��İ`�������ƓG-3�(���
�f�g5�J߻���@�)��2���|mtZ��Fc��g
6�_
�6�����Ц*��3\7��bq�vDUg�Ҷ�ZD�yVyZ�%S�{�a5�O��(�A�G�rt+�̱C.� !O�H��ө�'�'#��т塱Q�#� ������	[{�cV��2�)�a7�l��`Pcc֒V��bL����ӿo
5=��
hFI����t!q�����c�H�����KPx)e��EO)�E��đ���ݗ01�$�!Zu)ɦ���Ǐ�*AVj�1�;,l �!<
����.At�Q���g2������p%��xq-+u�h��z�SbcG�J(mOb�]0�P�����]����^��5j@��w%*�!P�-�f�)#�m	�SdP����Pp2�(f��˻<RG$�/�O�61'{қ���׾a�"�j�)�3�-X'���o�
տ��M���[�_�)=G��Z^���Y������Cg O�5uv�#�tsޝ��&CF@/��V��Gn^eK��ç��N4��~Sh��d�*��yTu? �R��#��V�5ciǮ���CE��i��lC��D�5��fPN�ԙ��{�|�!����Ɉnyb�^�Q!P��F�����Lf^X���@�]���[��ϓ�-�Q�!�Q#��9n� \�����o�إ���H"���7T�4����yb�z*�+����W��a6Ƒ�[���H�����ғ�{{B�7H]W߲R=�����ߘ��<�PZᩬ������qx��j�%9H	���U?��Y�w���¾3i��8�����m ���^'���nη�l��/�f���Sie� o�P\sc�������E�s*k���2�tK��U�Y�k���	$��*^V�{��B�z�eVaS����W�W��Cj������S�T3���|�B:]Jg�ɶnINWc�O ,ۑ�*�K���Ҁ���;�T��֡A�	}�l"����t�^$���MA}p�T(�����Lz���khg`Fkvx�P��yx��Y�~��TT�*9Ԥ��p�	�Q�a���ڜ\�p1p��Sǹ�F����[�_��l:Ǫh�JMZ�B��q�{���P/?ɦ�����Q��H
	'j���(��Ye�7�x<��H9���m���%[\��q���qe��YwO��:�4DBë�б�R��dy��]�΅��}�fEE��|��(D����m�@j:�Q:W�>L�\��i|R/�M�5͍�ԿY������2�Ʋ5oЛ0�������d1�܅<]�3������&U�����jf���m�Fګ�V�O���3N�a�OU0�`�6���N D"�j�4M5���� �Q�"^�"�����)�!�a�W���������xf�r�����SL��m��)(,�Mt�r���T�˱�9|��B�Q>B������X'-��|a�F��0�g[�ne|!AD��]�䪼�C��
��3�Dj�p�����-|�	A��P�<ڑڦ�l�������M7�{Րӝ�\O+���x7�v�.��JH�@f���?��9^`��zko�yM�nBk����!����-/z�
��w�DU�^���j�y�-f��;��9��8��W���۬)/�[����мd��p��i`w���A�잍��^�����nɲ8c����H���"D���p�P�
c&����fh��s��ǳ?og-����~�W���R%Z�
��O��n+�,O���%z��!!�3/��� /��ʬ@BY8E!u�d�|�A���3�-n���y2d�ЪB�]�r��Q�Sc/��@���7.�-�-�0@p�����~Rs��mm�Y�b��m\L�C�V9�e�
CC����tA�K	;k�]�^�qi	&5�����D�s~�÷3CWĹF�K�Z��w�ݫ!���/1�>���˕�$�q��=��$1:k.�DL��	�l���Q�ϥ���=�F�Vv�"?�|q{ն)ff0(��r	d��C�q>:�Mc�Ƣ�����\��;�7����_�C���CA���	��T��W���l�����΍*L��{���9��,{��)7��FU�k�!t�
�0UG�55��d\V����g�4�z��7b�tW{�ꢼ9�'���D�Rz�u[���b��h�M�g/�7J�im�y��v�uq���Ah3t�,R���o�%��d�nU��D+��ښ.!M[AZ��Q`uW�O�+l�E�a1hBT������0T����Y̑"�P A=�"����<�k��Ixtˣ�Ԑ"U2��ݠ'*��R�ڞ�Ʀ5��K���2@��E����l�M��/� ���^�H���q�*�D��� (�dv!~�R��KQ_�'O�k�P�K����	��>@��ʊ�W�/���Ɛ )�׌�H�
�6�a|����� �G�k������?��t�/zȣ;�M�I������)/����E�ќ�:g����e)j�5T�=Y���n�3��+A�W>��ܞ
 o$1��W]��z�v�L�!z�yh4�Nq_K�t�%���!)K�"��_��;7U�ܚ�Ş�H��o��|)!a��b��_c�u/�։��e���*
	2	F��Y+��8������f4�s��Gmvz�
�2"��)��j`���Y�ϰ
?�ސK��hI�������e�7��n�@c�����/|-;YT�3ǩ3ӊ��?�w�ɘp�"m��]'��
��k�A��N���`�n���1�b��)�h��{A
�^���o�F^~:*�_��ї�)+�:����^��$�5q��)֯�|��pm�$����[b����1r�+���?�#�H��?,Y��Y��<���T�]Xĉ��
���k�B�%�Ϫ,���Ă�+�,�ceYн�.K����u-��N���}��^��pw�j-��0��\w�Fa#�ѥ��Q<qDh����Cj)�_�.��A���	'AG-n���U��j5��
!�Gu�mM�}��t84�C)��W\��jZk��)��&P&���so��-�"MQ���ю��;��=��%r%�J�~6����*6(mLҨ��؅9��4������|铂w���G�)�4V��jE�v�3=m�ϣ87w�!�z�tH��o���w�?�XC+aF�aem� &���i�� 5Yvb��k��K苹_�8C�\��ۉ~��q,�f��x����ڊ��p�عs��F�b���z�xgZ���H᳍��p=�A��H�Qر��lp&�n���<D�+]BRʥ��˰��̱Օ�((�W�+#�`���̱=Y���+U:�j��b�\�H9�+�ñG��0��<��Q�_��E��9�H�~�{��Fd)�	�>�h�օl, ��BVX���<�+�޹��J�Ծ\QRP���X���X�[�RK	_��j�/�r.���,�D��&��a����|:WP��W׀i����x�@������-����?���s\O�Am,�����f����l �9����rkͥ-~�h�����~�B}�+`�P̐m�B����<��l__6���1���	�za� Hi�#���{�f"�zf���L/� n�Y�zC�l�2B����:KV^�,t_����k}âSH�� �`RS�Qu�I�/B%�&hEp��~I�$D��<�o����JgOMk�d%Q#����e�f�w�����}�8�K�n�[:��D�h�d��h�;0)Y@���J�ġ+�]O3�>�`�"J��f.�n�@��cD׳H��'�|%y������������9	�˾��1�;٬��5��$vZ�Z�s��B�2+���?FED��a%`��j7���������N��I�5�o-�9�c�"�;9�(Aa�ݑ�&��'���S�w�_Ń�}[�e�2��O����}�я�ک�=Do�K�8o��d9�X<�o�L-�'��8������'�\�|�.Kr	 G!��p#tT&���8�,��R�.�jq��̟�{�.Vҡ��g���^��� �q��t�V}�[��
��7>���p�;������+�|�6�[�m���[�c����r�%-�<<a�.�f��3��L9{h&�������=�m>��̊�
y��/��C�nu�U����?��+��MX�=��%�@�zˌ!�yF|TX�HR\?M�n<y\��2�"�ä*k�S/Q��ZP=*��BmSj��*���.�4M�E��G�)`qg�����X@��wU~�����,�6-��j�Wĕ9=�ǚ��F+�B��ޛm�H-=�d��T1�G	<�Y�F=n�����#��[�:sO2&�)̛�Z��9����|74�|�üRp=D�d�(7���)��)����ĜTl�9d���fbK<��0���9�;q�r
���इɿ9�X�|K9�j���,��#hs4��̪AP7�hM�G>���l��@U�v�Pj�+�a���^��~%�i�'�06���-��Y�w�y(z��R�M��P�R���tq��.Hu�u�"�ݛ��5�L�����siŐߊ��ÝC�>�wc�淭g���PB��E�E�͌w?lr���Ҁ���:Wn�J�fV��ay��)0f��!LF��s�{AN�>t��+�#;m!2�����MR��]��2�e,m&�]`���jљo�:�j������w�U�:���nc�X��������+��#/��VA�<?�X��ֶ�p[c�I�Y+j�2���|Ω$%V��H��Uo������  `�|��9"nv�@�%��)�
~��g�%}! -*��qrl�]���׌S�*��h;�M��� "j�3X������P ;�R�օ���r�*�(��n����1Ƭ��fk,W cM&j��U!��K����� �e�ˇ�3�̎��`�H6u����=�W6������ �"R��"����.Z;M�4gtF�ɒf�LZoG�͛�q��&��K�����9�[��I�!�!�X������o&pDF6��+V/��7 R�,��*���3���L���/��\�u0���L�k��0G$�'כ��g�������s�*�(��Z������}�.j�~��=r2�(f}Ť���bLk�c��U�o�-C`�BO���l�:c��	�.cl����b�� �5��I�Z� �

�2-�?��%b�M0�h��.s
��#B���ł�
ɹwW��8'�[�7���S.��V��+��ʲ��S�.��?+푽��2����-�'*�g���^�0ob�Jc�\�]-'�}� �eݯQ�l4\u����'+�0o��N!x�B��g��8�G���(�5(���:�Z�&;k������}Z_&��դH֫̀�6s�J��bw�0�tTfC^ 0��_��ZM����E���:�s}��$��w0Q(�i�@-ΔN3�󨜶/���I�mӚ[��6��ء�jl�"�	�č�#�Z��cҬ!*iԉ�5�:˗Ӹwm����cO#O��{(;��TUਗ਼#�#��d�2����K�H��3hJ΋�犰I*2��2�J��^W��<�~�k��$yϯ#�e6Ĵ�T�����l�6s�Q��R��y�ꤜ?(2�h<%`����Ť:-k��^I���4�mmUW���#7�O,�a�e�./���Ӆ�E?�Z��-��|��}�Ôt���wV:"�u�9O$e3�����R�9�o����W_V��J�C.� xu��.���Fԩ��N��&��;�e��UV��Ŏ�+$����(E��X̮B�<��[�1�I}�e����M������Z9W�RI���4L� �I_�,#�qc�>��|{q���ً��:c�NC��$��_?��+L� ����BL�L��2)>�8o#���N?�W�*�zC�	]�F=�o���Եy����x��"���Bjz�oZg�	H�٣�I�M�|"�U��h�}QQpj�_J7���o��WY��@����R�wTacO)�u��3-�mlwZ������Y
��T�m;T���h�y���4m��g�>=�l/��/ԛ�X
��v��(|7Q@�]������� V����+������D>r�C�f��$��3IGHp�,'Ņv������^<��z*vѷ|E���'JBI�K@��t�a.����C�p�b����rJ��(ۆ�Q=EĹ8}�.*���l�Q�����xo@��A{�������XƏ�L���*��b���{��]�~�����"qٮ�!c��O��Y&����ʴ�����-s���_��u�1^�C�d~��dm��
��`�򁵈���?��Z�Ԅqt1�s�D@_�^Z���������;tq�/W�Њ��Q\�1(��\i��z�>Q��x��ɽ3��`)� �@i����>���-G�VP<���x�-a,�U�
���-f�g���w�J��4�*r��i%�K�������V��y�W/a�\�˔G9%� ɔ�R�ǖ��HOjj�i�[6h��<Yvз��i%��񱘾�k�~����0k��8e��k���o�\�("�ܦ�I�_����![7;�XK-L���f���&��
��Ҭ�\� ��~V/m
��ЉU�.�֔��Sd��Kʧ$���u��?��_�X#��p"�Y=Il���HF�&��(�Kȫ�ׄy�n">7�a\�(��(Pb���m��^ߧ��~�p�%^c�up��)ȭ$�"!����3\��
=�0�ګ�@A���'%#hb'��mR�L��m��S3�!�yc�D-�@�����y�����@&�q�S��FO�Q,�Y;�z�j�my�ɋ�6iQ��5�M8����A^�����p�|s�j�7]�|u�yR3�p�_�3���<�<oz���R�����|�i���߶�t�f�j8~X�ڦ�
��'	��J�l|�Bd1��m�3���f�K�k���@���V�ѱ�槺��X�nG����v�;V�ۿ�DI��Z����c���ѹц���6p�y0���4Z����n���/��Z��<	i0�x�oH 5m��?3�Mb�Z)ʲ<gK=j�B�:������J���"�l������'&�T�}Nn</�$K|��"�dІ<���$���0L"�]�����4�)i=��Rp��^�D��XBF	��S�H�����|�HR��7�P�/e���%���%� ���1��nk�$�nt-a2�zΉ�����ь������ʩ3�19�ό��3�n ��h�&;�k��J�ߔ��W��dr]t	��~eD&�'盯+-y;�*�\[�޵>���I����x
`*,q����q"��7�l�['��yJ�����t���ܾ�̻�Oe7-&� �҆�s����٤�j@���l�f�9�����q�:W�W%|����!�߶Ʈ��h�N�.��P�`�«yjW�<����~��=����� {l�ƅ���n���Uf���m�
����^�J>����L~[1TCApP����`�,(���sQ������75&燩#���������KE�g�m�H*`t�hq$di\�u�>���ze�iF����Tx$W�|�.@z7��M������p���S�8����y����e`ڑ,�P�6�	�^k�9�2!�۞�`p\<=,����Ązy�j����-Jq�!6�����>ݺ�_�z_A��3s���pQ<���+��֗	����i�'��?����u���ºG�m�~���b ��>��l���E-!�O�
�A�$�îj%��Hٌ'�f��`�Ũ�V~{��Jo�L^ݿ,�
^̴?���f�wXvsR��&X]�)`��?��]Q�؜����a"�Y�B��L�����T�~n�� ttn=�c����_z
օ	��պu4�� ��k@5]�@H�l
�:��ť `M!�(�\�zNS���k����;���hk�'����2\1��$k�hdWAA��1�{�|�@�N?-��Z�Uq��3��6�������!8@�x�A�Y�p�_���͌<g"|{���N�q~��]�j��z��D�;|P�t�N�H�)�o�L2�<j�A�;7/��q�(��MȂ����l���ӆˬ��q6����`*CHpHn;�lvqHʨ�~�I����u���%�>!W���[{}2���:��4��;�yR���Y���v &1�AF_t��N��`8�Rj�[B)H~l[EE���n�?�Z�wY]	�РT��>�:�[��)7�ޤ�٘�����qZ<G(/����	B���a]PZ��5S̷�}�aj����%�}��a:�P�>Bd�ʤz~w�Ժ�Vhy-lG�3I���(��Cz}�%�ܬAD��i�\���F@Cm��N� �5�G�3�|�+�,������-������P�x̚��+�n�9Uy�ekD�y����X��h�<�����G��pP�zNl7�G��
?��'$^���m5EtTT�D\�24�\���#p��$�i-i�;�d+!�_�GYW=���X���+x�c�I���)�PY���}�A��w�iV����œ�n�}Vg�c!��23�q�U(N�QB���@�G��f���UT��C��������J�E��)t�#m������y����Bv���Y�C닎'a=I+`f�W �*oI��'�������w�D�*����Ws�03�J��4ׂY�.8�Udj��*�Ϋg�kΩ�^h�\&T�&���AR���|P}.QY�F��MK���v��D��&0sE�u�X����%�m�` ��*��{B��'ЃG�t��B��>��Ȑ��'1�zy\䱼lgY;��y�\�3}��h�κ�F�=<ѧ[�/!�&�u��C��uRi�]� ٵ#Y�x�q��i�4<�H�����~��[	A?�PL�v �:�fk��5 ����\ab�!��(��������l������K~`0a>��"�mU�d#��pBI�`�|��=�Ć��c�Nx���p��,7���c��i-��f�ԏ���٤������ł�JH�����y&�T�/��9���Ј����ǣ��Μ� ر���A� �$Ii,��	;
���w�4���ʧ)�+ne;�%�؟�.Y�IP��(.���)jƏId�A�T]�@���s�����~�?� ��%C������u�n-��+�����x��b1%)9^��V�3`n��%M]ۿ��,]�� �^ΩK��S�-���B}^�-������a�����,BEh7���o��9�!�6)��;>3����X���eBV��<���f:��qۮͰw�,'�0,(�$�O}V�0��n�f��VW����D뤊A���'gˏ�����y��S���"��<D*�Ȓ�ҽ�DIi���cZ:4�o�w��&��zYG蒅C
���.dL�m�2������2����.0���yǺD���}S?sh�m=e�[x��^�?OM�%��b��Ʀ����y�u��Hw��;���+ـ��K,apUp��Q�PJ��,�b�r�dSRp�ȍ;LMU�7U�V�������˱�����Ř��q/[�6�u�_�R*g����܃%{����5b��3h���#�
��l�(�$�[��̮��A����X�v��sKk<�Zn�v-�"л�jH�;Q��ު}��<N῀�6�^Z���fq]W�0u�p���F���+�!�&
��[��k�9O���*�uį3~3P�l0֛���Z�m�×�����hp��������R;I� ����C�� ���	�~�[����-�B���ә'c4��ۺR��	��F�Y���i���Z�(|r.�W���_��=g�g�M�xP��l���F���s�T��g��vqvE[}���vH�v�.VC�=���G�0�A���=��P�8-� ��Q�׏_���o?u�ArH��0p�l3����O�.��íCP�N\;ޖm�|�Ju&�~_6j��Co5O�'g��+��6�:E^�W���Je�i�%U|��l����/��[�Z�qc��g>��b�Q)*xL�
�*�a��γ��  ����?cƷ���g�(#�{@ڼD]�3��dg&�i5G�Em5)�@����Ac�;U&+e3���p�.z̞���N=k=-7�oF���"�s\�ׇpF^��"0�7�h�XY�q;��W�)B��7u[Ǘ�O�A1��;�^K>���a��M������B�D�	a�%L�����CӢN^���Q�f���*͘"4�z�,V�#���C7%G��i�CIZ���o�v88o��)����%j���O�K�{��k�+F@�{D]N��IV�ͮZsJZ�4���a�"=���E0v�I�Y�W}�f߱���v�*�D�~㸂壳ƈG$��c���簑}Z���S�>�~�j���"��-�5�譫�g�_,�W �<�}VO6v�Q&�\�%�k�����3Bx��⑝�����߉?u��~+��fw},��}��Q�����@3l�1^��0^��d�r=����H��d����;>�_U�s$�^�Ys���k��=���gq`K�)1��+S�!)���޻�r��܇�*|���`C]^��plJX�F,��.���Th�%zV^�u�c�r'�TT��}��h����Fkh�2�^N"����<y)r�"[�(��^������0��3��1ҊS"����Bg�d�E��!w��s��1��>?��͹�Bf�02��t������Y�^��#Gxf+VH�^9��)�s�6o9�����v:{Ŧ�rs��J�����RZ��R~ъ}�~x�+��x��=�w>��>
+O�vDB�|v�p��m��?�ߋ���_'�ӫ6�:��Ԅ&0�c�%�=+V� �ف�Y�-!��4K��|1��uM|	�셷��t���hX��EcR� G�[�DF���)m���u��q��u�GaA|y ������=�^�M����5�]Ҝ�����/-���ؒBg%��2u��$�Yh� �u_	��l���Fu�C��d��A����%��!�dr˅�"�&��2F���>�i" �}Z��K���K�(�>��Fu�q�P(���4+T6��G���g���A�ϫ�lɡ2�Q�=�Yxk��uD���#�q�OnEPu��^�>�@�����`�@�a�!^����NaWT�jcy�Mу�*�𱽰���Vm��;��i�-�u��aRP�/I�&����
����|4�W^u"X��N,�Ky͍��X6���O���.�^Ҿ]Td��}��$e�=��h�����t�.�wa?�����!E����Q%?lwq���6�d�Y����\� ��٨��<�56-�H,�X����I��w_��I�C8$�}��L�>.P��G{�~GX�;H���t���%�~{t=�{V=S+� G#?�����$;Mu϶
.�
�$�O� N����u捐va�g7܆u�&C�t��m�M8'+��z`<�x��ِ3LХ�k'�Xw�Kw���q�Ɓ�>��E$�̺���m���+����.�W"h)x8�[5�*�j��j�x��{��Ġ��(D��2��S댿U�dK�6f��i�6����/���:��*�Qe^Vnڛ��!�E�V97��YEn&����zC���4 .X���_��Q*���O�Y���jA��/0�9yr뽂�:J=aT�=�#
��j����ǌ\�)������`H�������F�ȟ�R�U\U0c������/s4`���̵�4�X{K��LkO�Yy���6L�}Xt$�$Q/N�ԆKq&pn���V7p�d�W����,-!ګ�����6��居2�w\!2�qC�}� ��>���v�'<�O�'c�z-����$l}�X�ՄO�>�q�6^*�<�Z@��لn�!y!`�p^:>�d�U;$��pJ�c�ZX�ܦ�#���D-KX�S�:LQn:����95�6.!��o�DC��kP�oW�Cc��~����>�vIM{b��?:��\�ʙ#�lǹ��.��q�d��&�d��,�a��I��I�q�(�J�$���x��h��Hd��^+��F�K�p�"� �Q��[�s�X���++_ K�'�J�����5L/�C�ڡB�hw�M�p��}���ʉ��Z�I�L>����<U��ە�r��6�h�,�c]��GMY�6�?��Z��+6�9?R�ݧ�ԧ5��#Qd�'.%�9���z˛/x:��[4��:"������se�����T�@�ίby�h�eO�<4ѝTO �ܐ��_�}9�c�l��!6k�U�0^���61�����ԡ�0�� � ���I���z�^��4u%����F�v��Ԟ؁D��f���P��C�{:�<�Q�8n�ߛ�_Ӓg�z��U:��` O��\����L|I"���bM��7�!7�'韡�2������t�N͟��(-MI,������T�����5J\�0wkx��r�m���-@	B�}Zv�h�����Ғ@��q/\��Z����Ђ�S�_g�Z.�T�P�zM��3,���;k�����@�� C�b�w6�+���{�Sx��R=\��U{�Y�h���Vd��Ԣ��ʀ�0�<�0��m",����g�=�P{�i{�L�*f��t]w'�>����_�˥;����<m�3Xڎhܶ��S��)4ho�+ˬ��#��m�Ȼ�ؿ]kr��y�+ER �O2 u�8�{NR�)xb�٨GƉ��H������8���j˨����Ě�ŋ�	�vY?���N��H�}�gF �Pe6�o��4�� b��#�AFG�� ��Y�����'j�����1��[�=[����KB#�k�1�=����?
.���	:Wb����&xG�W�5��NE�l��⦠����˽d��&�I�rz��{��y�o����S #�{�A��k���l9���_$�X�䃍��ȥj����\A�/��3Ӝ��-��a zن�u�m7��^�/v�PMR6Ww |�V�>H�sh�F��H�K�qq����zh����f�&�g��`�I4��V!�w}������0-�T1�c�Y��}'�H�����8��l�^��5Y��̫+�>o �[�-�uCdQ�p�vI��K�<�X��w�'D�-\��P�����%�͖�+Y\ɿ]��^�u����I`2 �,�$ry�ɦ��r�.�ͷ*��Nd�n�T���WO��~�+Ř_
�X%��"4�n�#f�U�Lr��n�d��7?���M�#�0I��K%�����q9��E#�ZZF)�bXW���{�hK���BUr��ޫ�9�b�|���zA ���6b�1�KBi>�<�t�?�8m&;�  "�B��:�H�H���{��"50G� ;�g���������At�3�.�]�j�	�48�B$}�\F�yeg(@F^���U���s§��U��1L
��U�5`�I�o�'�>�8>ќ71F��n>����+�2�S�YK^��g��-Ԅw<Θ�G�����a�`��	��:�DW�~5��|�2n��X6�"��Ҹ�]�چ����!���Α�j�5~�Y�';zkY���?[���|z%�wf�NãD�&�-Fϵ��t=3,�m�G�;��Z�_���k|"�Wlz�����(/�C�N��1�5دkb;/�.�g)�����)@X��Z(Ԋev�:�AaDi}G�v���Z��ʐ�����k�"L0PQx ΥR0Ob>�_�O@�s��Zc�h�j�	�!�_����h��Z!��u6�CC�
�V��O`�?�KB�h�Kc�� ��=Pt殸�Rhg �<vt���^Z����0�v��vO �k�Es��,\��D�8��K���w��wbw�%�د9���패�n�T����O��LK���/G��K��v��ԟ1� ��qr:Ɛ�@/dH����u�0�����"֏�Fo�htl��#Z�_����鏝����O��P$U�<�	[߫X��CSp�|eR4\���d�1�2/Ȣ�83Bq��ʁ�.o�Z����	2��k�_Hm��0����A4�)~�i`�
N��FP@&7P}��Gs����x�2���]?���_�ƻ9�ݠPu�T��7"RT�X��ر�@�+�ӈ��z�Z�JD9]���ܹ	�G/颃���_VG0[ �=�:JQ���q��˴m�,*��jr����&��0���V��1��|b.�l:�嫸E�$��H �!熦��X��V	����J�Hc�D��U�:ƮC�=��������zL��u ��A�5�b�@j�2�z_f�"�>�KL�ϯR����1�e��P�I�8?:魑�g��;
�r�FK����)FB�(迮;�7�&VgVmv����7�a���]<�5�׻])�ҭ@�K�º�0�������"���W%������d~%�;\��U��Jf� ����f��M��J0�Py�������(�pl�#������������(��~�ޔ��.7��_��`T!D$�|ԓ�5E�.�fM��JƓ��m�,��o4�>PH츬�H�%�MK��y\y���ә"�V�k�4B.���������d�Q�]35 	!d���*/0"�y�Z�6�]C�����Z�fP�G���f����E�%�1f��i�܏LE����|Ai:��3������v�0As�.o{F���\���F��%oS
@\�"�*��d�3O����J�jC�E��j:�\�x?��O|j2ӺN�鸀�<�ep�M�ӵ8��/v/S�����Wv��k�-L�Ma�z1�Δ��+�׭�k��8b�p�f�zÈl������L�`\�ɷ�蔞)萂����/�.������L�Q�bH�<�>�d�=�FU�\�m��GQ{�ң.��J���\;AE��5����R9�-*՗x�)w�Җ��!�`D������)�~is��iMyqҠ�V���O�[���u&�X���	��G2�����vJ���T��0���d.�h�-)B��C�1��q&�LԠ�b;DGӝJ��+oL��cP]�PX��ѯ���eekg>ޫ,���g�����{��q6�{��T�C��X�g!��~������|��8��d�ӼI�� _A�ƇA��F
>�eL1E��/�l("����Eh�#6%�s������O&_���&��`��,�.3���7>y{]�'H��AU��ʵў/����`�B����طfQ\�������qb��m�'4�&���C5a��k�X�_qX�@��
��t���*d�G>�>;�.{R+㱰}��u�J¥*8Q+���U=�Zkh�����3��/�D��d��'6����Z,�s���H�q�'���%�J��͜9��d�����w�[��y���b�BTh�1K��8����d�L��ւ���	p������-3G�dO�-(�
 ���Sw�N�ڸ��_Nj	�o�e/5���D�,p���"����T�
�	�$�'�ʹ�u��S�GMd�
} �\�e��(���VOy	�h�ՙ���P�~�W�2��IQ�l��j�ݝ�E������2��6���aD@�� :<$~BY�j6q�(�5"���K�2"�Uy'��{���DF����6{��̍N�+i���)��ނ�N�D����+��y�覷kxj6V��I������DH9y�5s��KK�/b�J��~[�+1ǁ�n�Wx�6�da<l%�գ��&��}|d���%K(�(+����p����H��V�hdϳ�{���7 Q�T~�
�c�c�+������@C�uQ"hA��%E^�0�t�$���������J6�J��ZE�����m*"����0�
�D��:,� �1g1�ri9`63�|z�]a\��T]�וNX���09O�h޵AM\O�#rݬ�6a����q�Q����弯��4je��tI}��O!�+ӢBA�A�£��b�4���M3>��H��t��a������Ijϟ2��(��N�4��"Wk�E���Y�͜7��M�3fo�� ���H�_��򿀙�F_��hg��=D5�c5(�W�����M�v�ET6I�5�p��YBp��/Vՠ��m�[7�M�j񒄍�8��q%-�]n�*�4T��ǲ7k�k
$E���D�����>;�8�h��n��A�]�b[溗�=��nY���3��	d���]�:�����RJؕ�&�ȏ̟&0�Dc��p��ȹ��z�C���Iٟ��G�鎆-�D(��~<��/=��&���A�J�~���jEe�~��.G���zS:n���}E�D8�T�[�Pq�,6��#��W� ���
�dyüC�����V*Q��R�oM�E�w�W��c�M��۩|���*g�RB!]�O��LC���)>i�]W!
nu��]��>i�$E�nl*î6�L^�x�e7S?&5��Sq��e����_ݞ����٤��+~X�}J�kl2��{��������=��=�2��	h����f�@����h�"p��_�<���Pޘ��m.�eW�:b��G�Z����F�j?��l����Ǔg����T�P�b�!�}�DkE")�:H���Sb�%&q!�JIk�=�̛�-���5(������-�4����(a'Ìi��ڔ�_	�crIxfR��6L)`�0�'�'Ƹ������ݖ�+ܜ�T1���l�=?�C�ԒHIE�j�^�������b���Ɠ�>ג���Q�RS6M�+#fi&�.kЋz1P3��y�v�
DF�A��ͪp���MIyw�^xND���/�����&�-����[*��	h������Q)@j~�1�)�]��ٲ���+C4	�Ӄ�Z��ښZXS[d��������rod@pT$��\u!��F�G�ٓO�[!��@�Gd��Ѳ�t�
�t����%-�KU����w~������i�X��}�fX��I��
U�u�&����mD��<���1}�P"oL��ě�j�s�@h�<��7ۢ�����ŵ$7C��%3�\%���c&u�U�nQ�pn��}Ϥ����O�Q��h
�a�<<чnJ�3��b����8񒥻��Sp�"�XPb3�㔓WŲ[C=�hg*��୥���c���l�nb ����/b��&'ж�D̪o����O��[���0&����_�%@3>�	�}_94(>b�d_R��l����kD��4�&�S,#���P�S�Cx
��F����k	9�Ϙ_���%�THx���-�����aV,�tж�B��^��_�نR�=���t��6��De�&/�g%�@'�D1g	�����������B�b!6��r�ƻ�w~�p$��	d䟤S;�i}dC�Uy���pn�6�� T���R��|Qڽf-�$x��y��;?����ԕ@�>�8��1���,�������E�T`����;d�5����^��� P�$ �3��| �G�A���7��f���U�4���4 �'��/ �L��&�٪kV�V�A�>G$���]Ӎ8��0?OW��-��j旔���;�^r!V���RP���xܳ�	�s��;<����������C�$�o��@���L��
�t�@������e}�^̏�䓼]o��ˬz8�/{�v?��������Y�N�K������!�"�J�nbYv� &b]�C̉g���x\���x���	��&m������1
��ݘ+�^^g�#/h��fӤipl[�ΐ���:���B�>�H{��9
��K�HW�C���:�(<*(P���4�`�*i�Z�@��B �F��Z��5�`�)���N��5GiG@Eځ��U���_%E1,��A��1�����m�`�=}[�
ap��2�=pz���靓��d)'����h�B�5g�- L�3zج�1kd��_��g������Ab*��M�����m-[���P��BV�RS��n���K�Гz��C�.Ң�ݨ�_��d��(���E��z �n�x"Q��TC�QD�����b
zpt���Y�ZQ���eo����S�>}G{AMH���}>��~n����k�V~��w��ӳF�*1�*1:���WRƻ���ڔQ�5��w�ƒC��h�۱N�b=�*d�sv�5Jg�n�����O?[rt��J����5��џ�ܾ�C�j�ւH�����7肶x?׋�Mrȥ�/�
g��P�������=k`x�����֫x��u�@CId~� �l�s\��z���Ҁ{�|$��cQg��R�#��E@T�ǡL�,�٨�G�p���z�R�ќ���qbyO_�S�mM�>�?~�m��V;?��{�^E(@	@5{��m�}Mv^^j?S{T)�rlZ��.��L|>�=f���+~A���ʯ�W�����=K�lCa�3���d�l���*�N/g�R�����-g�k`~���U/��=���t4�zB���\ �sLLU\�<�/f+h9K�R=��n�Z/�*r
���Q$�X�z1�b�ĉvM�N����>�d�lh�����^tf��9-O��{H���x
[�,2W+T���W~�(捪���B�}Hxx���e������P�¥~�8ۼ�$��VUO�%*cWZT�n+v�92���p��[��s�'�p�.�8a,��p"�e�,��d0:I�98�|�,c�*���޻����~����a����X��K���!Nz�'w~���܂�d��e��e��`B�_��|��z]3c��>��q.�_ϒ����<�U���c�O+��q�,b���x�N�r��lv�W4&���O:��~�m��hڽ�R=P�����e����Q0�c��p,�ꢾ��;��ʗ|��Q/����lN���7��^FI�J��<��\>̯��"�ƌ�m�I�A��O>������}Tw����g΋���ݐ�k� �Ǡ���3즄�EB;
A��xb���
�fW?����o�ߓ!�#����{�%|j�V�e}�m���#����Ŝ���N�qa��sЧv�!�%叀i.���f(�R����r�5<ɟ0�=A�|r�b�y�|R+�~�D�`�\2	�+���_�U&�X"�4V���\�,B�V%�g�����dO!up:A���m����XS��쿂 �T�j~��FP��.Tȿ�1�O�Z �7#�c��;�-�O���<�hM͋Μ^5%��/��冘�Ͽ �`2��0��M�����%��6U�	�Y=��ق̚SO���̀,{���AWڽ���ݍe�w���db��/&�C�#3�d�< ���+[f�ء�&�:�ċBE�Aצb`����芷�4��ʙ��ۂ��K���(S0ʁ/v6�uj+'�W��N�z��PM�2._F�6ɵI�g>I�"!�i/�����-;���N� ^x���އ�b�K��2Ґ���0+NG��vRe�#% PoZ���,Rn'�51�"'+����q����i�Z7W1ԇ���Ok���)D�;�,��{�1��^��U\�0n��>�L��uy�!�:~���(p��X�#g���'
��_{;��Wwzl�=	�����"(�'|�%ʡ�vIX� ���s�V��!s��F.���o��4�b��}�3|��[�{X��Vqd�9�%����[]ϋ�J.���xBsZ���Ok��?�< ϗ�h?�>!l8�z��_&O�^��
���i�����o��WllB?��a�ĂX����(�Ja�`��C &����SD�	��^�i3�x�D�ڭ�"�<{V�U��P�oXF�B�
"{m	���x��aW����}RLa�RU!
L��p�ǔ@t9��XM�bg�Jm���n��\S?�2v�n+��%�]}F��
�]%%�0m��;��B�~��Zm�/<S��6�!��J��rL<�T�ly�]��FW�͙�@��u��N�?4��Z:�O��.�wߴ,��$��~�
����85�=�M�Pr���j@�D5����*��k��-�(0�
��O�K4��k���"�[�!��!{T��u���\�_�['R�7�__u�֛��w�����r�Ç
��<p�	�0�*���8��0�~��A>�~1+j�M��j����e�:��6�PX䩥��mE���9L+*��	��m�������}���.��*�Q�b�N�e��h��DYU���N7FC62,��	��*�G���d5
�R��ܴ"��P���֞JT�j��n*Raƪ��Nj�n��N���=q��1��� ���N�`���x@��B}�L�olzW��6���b�B�^��Q�[�zt/:g�lS'�S`U�����˅_�H[�
p*M��)b��G��"^�s�_�'Ks�M(*�N����Y��6<o`�K9$Y㵌h�A�B�ݠ��w*� ��x"@���` �폞H�Hi3��ʩ��S�
�B$��(��i���w�z;�[Pǃ��ug���L�V��=��������;�Z\��m��O�[���/�E� ���	�G�;� NnVp�y���C,�<��hk�8q$�=&�g�Oċ�w����6zֲ�!�<b*EF^k0$���z��K8�<-�y-�
�(��u%P�􀲀gV�OҸ?�6�,'?Cc��E�/E�7��$1�����d#��;�B3{1(�uV�v�:N�g���S&g���-�c�\MR7�Ir,���},!4�=��U����3z��>H$��[���}k?�Cb��������u�|�J��<0L�Ac?;��K9��9�ʚ�N?��W��%��Z�N����R�
ZҺ�_��'a�Bewu0�ے��K[VK=�'�]nph�2��B�1~�����rx��WHe̝�MG[P�wR�ġ1�2ͫ0I��z��4���&9\�&Tsh����8���@V�������A|J���W9K�����x谮�KRĀ�B�^������y��o��T����nf���"�<~pv��BOҶ[�)��p��f(g��--��-�F&��)�Z�L4-�)�T��+�Hٻ�7��*��3z3bګ\(���g��Og�`��0�[:��wW�pRN�ے���2EeWA�&�v�@�y/��$=�t�&e%�󼆨.�T�4X35c��������������8Y�nq"1{$*�:q5)N͢�%/x��~:��ٷu\��[�=r�M��S��fC�&�hr�z�v��u�W��>@�E=�%�� �M&9F�\��-#؆����lBe���F�5S����F2��0q��݁nH�}М����.�d4�����6�)N������	�)u��w������7|�c�a'o4���$��z;�l�V��{�tE���v����]��.��1_xG�z�N �7��Ǳ[��n���i��ˍc��On��&�[��L�k�V\Y=0���:}(:�ޮ*�Y1 �'e�-�A_����c�g�v�I���������.�������\��k��[L;�9����By�ڬ�+�˪G�R9���g���ŋ�9Ͱ�Ј�\L>W��ʢ5ٙ..<��/&�iM�|_�Nq��sMu�Ǟe�+NĻ�:z���UX�c�O�͠��\U�\M��{!�/{�7h.�{�S�a����-�Ѥ�����t�_ �w-�����_Xܹ��gB�ɪ��=縇̖~MbKf��L��r8����`�Xp���G���fP��C�<T�*�k��Q^�OݠB҆���y9�T0�")vN��!DӾ���M�}y�62cͨм��Sǂ���T�~+�mq����2f`yy��6$�X�9���Ims��5w$%5������8���ȧ��UZ���<x�tM���d<��|{��R���
>��x��
��Ȏo4���ia�\ݖ�r��p����fnD� ̓�	���e;�$L;2��?Rpu�p�{}d��C4���$W�M�]M��M���UK#KzGy��Ƶ�A�<�T�	��c/|]��w;hj�Y���E��(��W;�%�k,��- p;��k�	}/�^�?9aҢ`ѦX�U`�'eV�ʣ�9��t�I�F�PO���q�	���C=@�`g�^b�a ��w�:#k lƧ^ #5g0�)�Z��U�)���hJf+�V�F4*	��<)����W-CK�pt���[����X�Bj��1A W�ĝ՗Z���~�}��H��d��ql�ǿ]�1
SH���e'����e�qu��9.gY/C�{�Z��_�������$�Ձ�%�H*K��7j���N�V�_M���jjkigV?�R����%�W����?Uy��k���~3)ޣ���K�lm��H�y���p�U΍�2��,YV�:L�1m���a)qY!��SL�K��ʟ/��\fA�\�tk�T������B���8����,n�׼�D��k�ןe��2��)�F��.i)_�s$�q�а|��g���}齈���Z��_�/�e����g�i� ��޴�@(z�������q�y�_���q~�d�aҿT;���Z���G�c�E�V��Y���+����M|%�V ��>)�O �ݑ��@{=���䓓����U�*��V	4p�>���r��V|v{W۹ÐD\�(	X]ؚi]s�cٟR��|����X�r:;$�ʝ@��:�����̍�X�����k���\��@����A��(l��tӊ���l�>�->�~+Vs݊sSݷ���k�`kl�@�\O;3����?�E&���$5��;Jlc4+M҈'�#�������k`u���R-�/v�_�t�a�����DR�e�I���~(��C�{��&ڎ��v� ;�)=O����2�_�������Ȋh^/e�
����|������8s\���#)�F8�]v,HCM4W'��0vù�E伭��H��_���S���$�T！�C�1�_H���!���D��k��\o�0=����̒$�_2{ف�F�����g�~�o�8����9��9�#۶Қ���`l.d5`x~@�%��5�������kk����Ŭ
Mk�����>hI�4�� �j�(�Ld�gwE8�/Lmn��H�$CV� 2����VibY̽������P�=Q��%DL�g�FN�Fӏ �� �oZ:8����<ݾ3$����_(]�pW�6��S�b�݇��q���#=�hd�x	�{�j{%��X�kK���a������^�}=�L@��G�dHvP�P�e'� ��t)5U�~�m%�gb���/�����z�D�Ѩ�H��!�o��֖G�!��%�d,3bl�gT�$�^�+���LM��Y:<�Y��A�"����Q�V`+W�7�@s�k%W8����k��4\m��h��y�X���{ !2�O9-�d�#Z?�(��O6a.�����!��.�J엎��Ay��+���W{x��
!�o5$|AEDC	�I^����m-��<uä������NQeE�	����IX�VFZb����F1BnF�Kv��w8���J`gǴ�������vd�soOF�.���+�K�ٚS��E\��2�[fr)},�@��$>������s`���Qǉ���q��Z�_u��i`�܎r��[�w�u��p`�D
$\��/�m�=�����b����4l�Y��5��K�]ۍў�7�����)�.�M�0�?�l_ ���3�w�{S~}�c��V�o������-E�6�R#|6��D��̈۴Q��ӗ�G ��lPT�/���Q���
ᯡW�M/����\i d���6�P����#�шLJ��/������y�c�Xk�*�Ͳ�}���l��z#:�I7�3_�!tV8������[ue����p�&�4�G_y��DX1�@�t��-�^�P��Ѷ Oޛ�[KL���8@4C8~��ޱ�R��l�%�WK	%GھLK�{ݨ��(O��:���I=���OS�z���)��e��Q�N��n��um�7,�Sg��ſ.��X~�-l��c�`, ua�tj�eLG�y[@G�����I� ��0���g*!���|���j��R�k�8T���}� �+
�K�����{ɿ	��_^�����&�I��D�Tt߁^�� k�=�}x�̤mL��gʍ�z�Q��9$�{��NY��{�zq���c22��l�����o�J��� \�p�^���SU�'`];9���LEeèޖ*����VW�\�5	J[ķ�{S�:�tHp�g�
t� .*�>�ho�����v��J�Ť�O�(<���ܩPp������r�Ӆ�M�#��M��4��?�X9��}�n�Կ{���{��3����'N,���L�Ň��� x~�e�����T%c��Ȭѳ���Fw�bcO�~�{A�Yx䳎k[����9P�6a㵹�h�$�c�3�0܀J��G����,j�G�k���a��8:�gCF0��\��[H�/N��o�E�/�S��qX^ag�MiF�b5}�KO
�Gn �2AN�/��Z<�тc�p���� �K�?��ORx�4�b��	��:��d^�ή��O=���GSl���4������8�+��y��c�-	vIu��K[��� ��Tʬ�C6�Z~?Jn���x����*�F�י��Z��/�$OB��i�+L���dxEy�#i�����Yt{���E�P�����E2>5��{�4�0+�^�X��
��ΠY�_i�+�jʂ��1��G�6�ż�=�U^t�-�5�f��s&I��c�,� Aԃ�&\4kͦT�J�7''����}༆�P!��2Jf�jr��w3���""Z����ٶnh�#�X�<z�!�Z�[����S����������&繅>��0��6y��?X��F�@V�m������<��~� ������$ �o�O��E�$n�7(ޅ@f檆B���ݠ@c��G*�6���^l�Ǩ�Q\2�W�"��ٵ������V$�z7��3�er�
���'2x\�F9�b -�0����=���ӣw���}��c�{Q��:��.��ɕ�H>��w#�:Mc�@�_+#T[���\<6n���\����MKN�]���j4/6|�⥀�s��m�^���jy:na>enx�y��:�<��赠��`qq����
13�z1!��,��i�tP��~Vݙ�����ÔQ�yps�A\�:���p�&ѓ���c ���Co]EwS(���O�rƇ���ُ{��ݢ��lM�0J}1H��
=̴��~}��A�ʘZiD�-7,�� 5�R�T��:nA\u�ڽi��;�|r�����3�uE�3�=���蠁����m�	�����ht�:����Ώr1��#C��� �B큄(�Zq¸��k�u�g���.l�vį �ݎo�txއ�8�+h;ʝl)s~,@b��h�a2u<T�V7=<�6>#��(H ̮M�L�"g)�`�+CO��b�gE�o�H?dM�8�Y� �m �(t�5<k��L-e�5�Vbׅ&��b	�4ۣ(y�/�������tG������)���\�&<����$�j��Ċ�M�I1�.��F�m���Nu5l�#�|�H�lz'O����}��,]h�O;񜧊Ǣ�g�b�S��^��J�I����Jx7CG�#[Q�Xt���k����d6Y^U&�#���ǥ�SrĐ�n$��i%pN���j>mm���fvU�ܱQs��=�{�J�
D��+H�Y� A�-�x���aC�ha��|7y5��^r��1
�S�LE#�L�K��~�y�[Ҹh{������vV;�R�<�h�\ew�E,�(�8�u��nv�Q)�s�@B��5�q�
�}'��-�
�>=\�=%�ȭb�c�fI'���׾�9bxF��{fƪ1�	�N�{��g���_(���V����Bչg`"���,
�%���:������K�c�5<��q�/qu�G�0������
����7*��(�r[܇��3�~��&���l��]�Gi�n�>+�m�	�Swи�}����~f"m�x���� _Y�e-l#P'%���|�M;BwY���x0�ty؎*j�A�< k����Z�ZȋM稇���M�4���L�k�{����-�y}��3U�=���9���Y�r`K��0�E�Â�>R���ѩ�Z�[J�"ˁE-�ꅆu���]����9�v=7�Q�{k�>����h5�#c{|Y�O����H�cTk�9���W��K6#����9��O�=�T[X5`�?����{�P�$ �I����2\�𭄘� �����4�Q�����W���u�W��ݓeN�^�gD����>*ú���廯��d�;3{Nc_�y� �m�����+�
f5I�;�����:E��߄Qz�c�뤀'~���g���8���>���63�}��/���(����t�y��=�#��.I����e�����ټ��$Uq�귪��*�F,Y5G���l��+H��'~�/8��z�G^����
�d��Ø�8�;yVLsJ��GT�L��"J������|��}�N⮐�w�|��;�4���/P9�(bR)9�H��Uz�.\uA|�����E��J[��$h}OS�64eZCܾ�kE/�
>�#%#�Gf�<g�M2��l���k:�#G�"�2a�ut��bj盓$A�S��^��4��fY�A4��ݣ������s��;��mb�d�5)���7=UR?�3�:(4ᕛ�m����#�٫�j*��u>�5��ߢB+�a�?;Q��kM$�E�#��7i.%G��$��UЁq�]�������Y�6���+�0l+�ނ4�F�ٖq6�k�L>�����/��;�4��L�Q1\��N�.e��>�!20ϊF;1C����J;��	�v�3��*�\о9I+�S�5��M��h�X��bAF��$#��%4�[���M� �=����h�Ez�-ȏ=i�Ώ��]�~��˟[Qv��d��#0���:}5H�To��J=��:q@�k3�X��Hf��A��=9��	/�[�D����Y� ��L}��إ~�T�f�|Z�"\�!å����$�M�#�9�����0�5�*8��?��/:{ň|������$Q.qW,a��a���QK$�|�:Y=�w�\Ւ36����hx)M�;�ۓ)��2���|��neEː��Ӄ��f.�ok�{�,��z�3kby�H��h�mM��L���Q����مWKh���]����u徏��;v+�q�%]WDԷb�b�|�Q�>�p��5a~2�^q��V6�R��������L-��w�<Fe��>�G���bu�&��������#�AP!seg�E��pu���u&d7L�dL"S����];�G/��Y�V'�oe�6�VK:ցH������}�D��{��e����@��@�FYO�ߙ>�� �F�i��BСɯ��˳]��������PE���kǤ���Q�����;3+;R���x<�Ӱ,��h�:�sCv0�D�����̖�M�K�> ����C�5 �Hq6���T)Zdt�!�CL�:2��<w��(�.
��<��_��AҰ�O)Cj�YV"�)��]=�8�K�	�C+��P�*���eLJ��HA�9H����I"~�	�8|IV�����P�ГN&G]��uibg8T!5���*�s�Z�:D�3��W`�xb�ZI8�R&�y@`��̦�Cz�9�������G��s�F�/�]I��c���H�=JE��YR7JA��8
(�k��Y�d�LH6+���{�]��۲��14!��œ�Zl�4���M�R�*y6���qg���h�[�����%�����TDÑ�C��ʾ��b
}�%O�c��ycM�&Y�?bYI6ɥ�u��x�����5���9�YZ6�����������;���:���k�yᕓ����:�>�Q��i�Ϟ���S�����v� �h K�J
��n��`֘Z�k�}�M������G#o�ŽAb��	M��w�Jw}��A��vq`&hʸk�=���{�a�w��4*H��j=<�-���6�*��t?�1��F�ߦ�̂�塟��C�bM>��,�������<efԏ{xpd@��X��a#�<=F�i[�c3$�h쮱}`�[�m�>��޷�IS�㚨��|����ѫ}&BQ��P�2����4�脾�BE�a����(	iB@�t����qr���S�¨��%2��HC�8e��h;_yCE��FC�|�L��a�|󤪉����?z�{�S����
1t<�mi;Y��$w��s�1�^��E>`6M��_��;�tT>E�7|���z*�.��5�z���i�Zp\� ~|���W-)�AD_�2Á3lࢗ�x�}�/��Z�q�Uw_ϼ�ILj��(�Z"�zۚ,�\ �ō��F��!P��{<��rЬ�����x�P�s)\���B�o�B�Ͻ?�;.)&�~�\��OZ�@�spD�|��ʲ����	�z4n�B�D�2b�S���m�H�7�~���Ǻ�;���1Ou�Γ�h+��:�~�
e�����
�t��,���ޅF`l�~*�e�����(���-�X��k�F�āB^puI���p�p6ٸv� lmF�y�������x�|		m*N�j�Z)��,o�?c�>=�gl��o}�$,�e��[��?ȝc���}>+X���Ņ�+.�I����&L���͎1g9�}8o���w��'����Ǿ7����2o#c|t��AVCg$dx+}22��8-�����ɜ�pQ8�\��R���qP��%��:|P��U�}�閦2Ѐ�����w�	�/iI�g�%w#��1y+K&� N���ց�̒_5L�;
�x#"�Y�/���wNY��'�6j�2N���5cb+�"Ad�H�=�o�6iB]t� 0�o!�
Ƃ�kQ#�It�)��L� �B�{zS���Cր���kP�Ά�5:�>�R�%�
��Je\�
7L�P�.<-8t�v���
�`�/2k���
�(�"S�lo�#�����%` �TQ�&Lg����t�WVK�u�c ���R~:=i���eX�~ųa��)���Pt�&<��d�^��ީ��>��Eɂ��K�$�;�`yD[/"�a.f-¸�Y��D�e���U�el��̉�K�ǀb��q�|�J4+�̕Gg��k�+���Y��H�b�D�<k���yt��-)ϐ�w��^����e�$l�<�5�-{K0z[�ҴE#%;!Y�����e�DX�䟬���r{_�|.�ϱQI��iy�i�L�5��E67�u��4m�-8�*�W$.����t��5�Ǐ;�=D� +i���b�O2�z��I ���|�@v{z$�M�.P��sM��;�fMIR�	�c�b�>�p��r�l�Ґ�3��?F���Pù��̨�z����aH�\Blۻ��}�詏RCp�5# �Q}m�C���	�.+�d%Ə��{Hjt�^ã���ʠݜE��8#�k�gi�4�(����#�a����L@|%K?Z�|�]�	h�~4� Կ���N���m�@���J���y�|:(<z�A<Z�.�" ̍�YmG�^F(��f7���#�
t�M>[���]����8�x�
�+@���3��!z�J���_�f�6^�#���S(1-ñ�+(9@�3MJ&�ʱ��ȹ��Z]�t�z�f����>�8�7��/@	X&�l��sV҈�������
NI���(L�j�~H���2AޣD��uY?�:��� y[*��g���=�a���3~-���C�_;�����Cd05�;FA�nU��r��] &�R�����������ͥ^#˶�"QE!Mkx>�Ζ;���v���v�<p�9O;�ixɛýZ-^7�
F>��<�.'#�}(|�]k�!������>AǢ_{�]?i�Z��߉޵3���y�d�R9_TA�4����/�]��S­눶�D�����@����KJm���w9��Uh�XeC���6�xj���5�#!+ρ~�3F+8̩�XO׺��+?O�~?�k����cM��S��*Úr��䲝��	���|X�!��_�~Ɯj��2?0Eh��{2���Dy�{��Z�`^ItKH��PݴH�����T<;l�_��BE�Ck�j�P��*.�7��A���9��R��e~�2�����X�s)\f����e�s[�
��p��#	��M����1^�n�a����d>�[G�=U7������X6� 4���9��Tu�xaG�������f�5���a���xϤ1_>�?[��R���D��d�d��9�|�`�~�� [�Mb񹂖�xc��-Mf�1��<#_�S>��t��k	��xQ�n%�XcN�l�HFf�g9��}�����=��n/��ַm�+�ъ5HUxܾϹ��RrG$0��m��u�@��u2R��>_��E�yH�9E�Y�"�/���@��?�����+\�S�XB�l7t>�z
�M@k�'�T_�G���S���g�ո�ԡ�@I?t�!g�.GZ��L�\��x����dU��?�T]�j��m Q�S�0xs��r���(?�{�;�J�&�Rw��ίv+��N��"��)�n��TJ��W�����$S��c%��Ha�۝�+�)Be�F���l#���w������o(ӣ<��T5�z���n4�,e_������2��'�3x�b�����. |�F	�:�3��=��@qV�
o��:�g�85�N�& 1+���� �p5^H��N�d)BWhj����hѭ�-����I�1���;���Z�sԦ�9*�Q
L�U$�X�1� �g�ɱ�c��	�[�G�e`qhc%�[(��R3��.�;��)mY��K��m�-��+�1�V����3��z�PЕ7�gϡ���x� ]'G�G=�ynpA�6��璀E��v�w���6G-KƷG���L���~����� ha���Hx��3g�1.��5L��Zx�\�E�������տo'��Ɣ�2�J�f��H[
-����zZ\�d8���`s�hr��g�Y!�!�&�Hq��"�)'�@�x��}Ќ�B.�r���Y��d��P�`���Vߢ��̷��F�D����>��w���omV,C����drR(K�iT�򇂢�7w#C�[��6�������F�넠f�^
��q�a��#�B�M9��@���g!���ә��EoV,�h�h���E���3�5ɱ�r�k?���4�Ϻu�PUg��� .S�e1K��wR&L^Q52��R�b��<[e�3-E3��|�v�@��0��**�\K�;ҷ��, ��Q�P�RcF>���YdA];c��iD����P����oy�E��$��F�[M@!��Qzn5��qV3��po92�m�8��V&E3O��W���=�l����d�~���,�I��Wk�Z�(����ɽ���u��.�PO�?�w�&�#��hv��y�rhF��Q;��M$<�`⧐����=J���q>V���8,���8l�4/���k3r���#RG��w�A3��������N�Bd�ݜtOvߤ��#�:7��tϡm
Cm����єG���׿nZv9"N8(ƪ��`j�v��y������G��/K-_��=l�/��^	�QGa������jG;$�[��ܞ��xN6�]5d�)�s������8�<���x;�%��{�hm,����yP��)��`JМ�#����-��y"(���+~HS !/䫑"��~l�L�r���E"L��W�7q�q̴��:;�@�W\�T?�M�i����8#C%�����\��z���[��ڰ��D5T~ł�F�%�2 A�d��	��h|��<�MS��+�q�g�GIO�y�����o>}3϶mUh�$
�$h%c@L��v�P�C�0�K�G?�����
fU�,��V�� �⾗;����\��6ҋT	5�d��٫��ٔҹ-�9����N�ݣ�����ۑ'�4���L)�rT%����ʟ��@@�y~�C� G�]n>=ZD��D�!�9ML���Qėc^�k���K���Kw*Lj���n��\ݔ�6'a�T��\���X�@7�vk�"Y����ް�As��mc]c��ͬ����l�+��`�[�p�<>g�nJ�8"(q��4��Y=K�Q��j�)t�n�F����Ƶ����eC�?����%�:��@�%��8���z�B4^ �_���?��Xg:�����vt �.�A��j�P'��i"�!�󦕾Z"#�����UXfd,����>y>\:|޽���vU ���;�ʇ V�y��]���gx��hg'[�Ɓw���: �6#E�p?��c���!�^�T���[���!O�۩�����Py������e����ب��%/�?�&%U�_w<7�!�7hu^c6�KɦL��}�C��[fS�)ǭ� �.��ҁL;�x���`#�����p�]�J����<<�"�p����Vܶ�~]�M�J>F��$��K�J&9;�w���f8�[C�q�3�����Z�Ս���I�4Di��BLg���s�N9��,]pP~�)߉vy$EA�_��
	.ʝ����q�-u��h�a�}�&��E�����	��%�P{����"��ob��3I���X����Z ��"V��O�uv�;�s����>�����o;������j#kRm�����t �D��8���M��i�A�ߗL��tUL��Wb�ק{h#�z,K�Z`�$;�;�dR��
ȁ��o��ǻ�1g����i��]�#l�/[�*E��e�_ ����!a䛠�b	k�f�����S�+��:�ɀI>�F��dTx�r������a&��Ug���<�%I�m�]�x��?Y�\��2Bg��;�MWͳ~�WG�,���j}L�^���r��[Iɶ�!D�Ub���Nq�v�;���u���`to,��f�XI<���H�eW�ૻ�yj��o��{����H��V�J:��O���q������Ʃ� n�۽9���y�;��d�H+���������Z6�cq ���Yz���fa�qZ�6��ܛ��X˄y
���	h��_��N�਺Z�g�\�nw�eV��x��N�k�/�����1�?T蔾���đ�4�4��&��')�.����� �#"e�������6٘qx�R`��$){�.�>)H4�"�O����'�A�&S`�+�4�����r���8p��V'�]��/��q���	��R�s-Ўb�q���*>)bH����=��gd�ͭ���k Y��u�ȶ�A�no�� :
%��jhn#ZE{C��O�dfl\���	�h��f2�Y�㜚�
������9`������#p0��!����Qv
�n'����mI�;��-X"��8���,cA���Amg���FB���%�����&=��uf8��p2�z�	͢fy�3I�H0'��z�P�)�k�ތXZAX��,���WCU���t,DhL����a�퐽(,)��d���2������⮁�OKq*[��K:�q'�Ƞ<�{m��uV(�����: �W<��4���2H��:�[ڱ]Z�&�6��#!Q,X�O�`��!Sڃˡ�OC4(�D=h���F>H?�N3	��C�����Z���sSa�NX���XDױ $GD�=,��s$j��(3C�s>{�O�j^sS�CNr�!��xH6���;$�G�cy�C̋��0p��(Gp�
�.��Є���R,�Y��2�6<��vY�h�8:�G�����P���󂥲����.Qh�)�h�DUO��Ty�R;��"ķ�m��Ե��S)�'אHj&k�P�z6��s�c��r�|�%�C������[�����!J�ȵ���k<WK"W�M�5����<�ֱd����)�fǏ2}�ɷ�n��Ef,!6�rs��_�;�f�ܪ��2&w�ɏ�O mA���ߝ���	�p����n�B�'�锵K�,���K��,�}˶�ާa0y �xF����рߧ˗@�à��h9 �eӟ�z��N�SϻZ7��3�ē�����=+2� ���c��;�\��({�A�FpAT�j�ξ{�7����Yxv�6�D�z.ᴜ����8K?�� �H`)W�![�(-���ӛ�"D�'�C�3���{mf�Q�yCs_�I��_v�P�ϖo	���*t�}��ք8��}Hhq�Y��
z*�$	���K�����v���`�}��.�U����,�;C�N�.Ђp\�����������=��"悄 xiϷ�b���D���ɋNFe.D��/��3�F�L��o-1���� �<��ٯd�����d8eMF_���6m�:w�Ŷ�H8Ϙ oJO��g醠�|���e�mZ���eR��?�*�fb/���r�\Y����4�Ÿ�l���T�������Fv����.'Z�Q�2 y(��'���	n���Nk~����@�C���cA��,_#^֐�޿�28,'�����%��m~1wς]K��}��?�V:p�iO^��RGZB�⧳�O��Wt�KA�~��茠�����m��U?7����� +wD��2��o\ro�ր8�~r�Ӓ�F32�p�ɥjs���}^���Wд�����NX6���m'�ńre���ςg��Z�kbΨ�\%�����0���49��+˥v&έ�*���{���ðRh�[�!�qD�WYؽ��s���L�����%�&��zI�o��f��o��d/�@�k�@|]X�a]�]j�kL��!r���	31&�WJn�^�!�wJ	-�yzU~����#��h$^�aS�:!&��Sn�o�z���TS��>p��v�,ږ�O�P���w�-H�
U���9��̷&�bD������'�P�q��1k�Vˮ���jΘ�UX7X�PY\��7�$��Ú$93���Y��n��dt�I�*lC=�Y�F^�B�u��@@��$� �l̐�rP||��JK���5;ʥ2fy�--�s3�3�1\iە��I�e��p���t+)E����
�T�~R}T9�0 �0��_��W���)����
Q(<8H��ΆS�6U�0�p�}�Mn��ț9�U��̅~����ˆڂ��^q�4.ƶ��A��"�_T60@gW�Me�����\W��
.k4�I�ϯ�3�-�%�|�ѽ����lf�q������=HPf:;��Л�6^��\X��M�C���R����,�c���-¡���D7���SYh���$�'[+�����AѤ����>�i��጗42�G�7~@#��>��i��T����2�+��:2�!?BsJZ���E%�,cu�E6�P׷�M��C�p��z`�YkcD�����T{Nx��l�O_9,������zA9d6'�;x��J�|}��eHv���d%��L9+i�F@'�����h-&���U��WE���X_�����)��wZr�<�T�h{�^��#ٖ��g���Èd���F��R$��fY[B�
��/p��s5}����*�����.z�g���o\K)���0J�.l������We{%�O(3� ��R�Mz~R��{G&U��[R5��"������ҟ��D+�Qz�n�� k���}��|^�M�<b��\���ф�i�V�J� ��!���=�!L!�4#������Q+�D�"��k���	 �`��­ �D�
��{K�H}���Y�wÌ���E���^02힀d w�����7�G<�"ԥP�-'��e�M2�(u��)�;��q�3tN�K�ʻ3��xUN@{�΀�X�^�cbq׸�>���g��?����'T:?}�u��o.�탷���).������&���}��
a6��v�]%��`���P����7	�,A�p����i��?�S4`�m쑶�Ļ�6J��x���Iu�g�������R��J��334�7>��?�)X�K�#�/��:�z5��#�19Q fZ�ȓ���R��l7��q3�d�����t�Q*	��$e��Y����A���ݗ^T���r���T�?I�x��rM�e0/ݚ��WWM��RH�m}��91��L�P���Fs�uI"�����4�βhM!�V�#_�C0�:G�]V}a��8l�r�p�RG�vۧxxs���B��Zf�N�B��Y��@��H�3��#��g�	����~��+�������c<�\�4jw��OC�d�i$�<U�0H�c�����9�`C\OS\��qc;��~V����V�`���[*�a�Aܰ���W,>E�"���B+4)���( F���G�TR���<��t�<�X�0	d�϶�LZ�w�v���"5�tMt�F��Gᇆ��@yD˺㡬���Zv�]�U
-R���{HN�/[Pz �9����l�~­[g�תG�� �Q��$%�!@Ih��g��r~�|<$Fq�9���PiNB���4� L����-�f�����j�l�
���fԔ��I/8�]�nk;>#��-���;�q&$@��G��6'g*�b��fq�/�-Nc�^����%^��E�]�o�4�SxjG�h�y:�P$` �ʲ�_�������[��L�<`�E(d=��l����^e���x=�;���Ȼ�fX�O�� ��X닠�CZ+:5���8�#t�+�v����+��=���ިS �	;���M
{ <�Bg�s{+��Vވ`��U���<�Z���a�_�nw�4�<�8�:s��h����AۭX�k���]:�z�K��D�~�T�f�!���� ��Y9Y0D�f���ސ��^x�+,�W�;>�7U��L�t��=�n� 9ˋ��L�1�df��<Sü
HSZ����#���e:
")ol�X)?�G���4+��p�@ĒO�`k; ��P2�m��.��2�&�d$UǬ�,��݁��9��]QXa��>��%s�S.>�ey~���E,���b�7}���)H-���]�ǟ�V5�ZeT[�6����2�h�����w�9#�J�Dε'��Җ�҈Nxș�.ކo�Ʃ��7Ucq6���ðJ�&yV��T���wy�*���w(esZ&�I{���s�H��/��ѭ������=����V8&7����D8�4�	7%D�N]�ϒ��Z3��̦"�����ΠW�>Dɯl��~L+�&��x��Sh��-�K���2�m�������bA���4y�sxG��A�h.�>���sc��� u�w�?x�}j����O�VГ�w���H[�
�Z]ـ8��н�1��7r��u��/A��&an�����b���R��E}�E��{��8M��R����EE�V�8��s���#�58 �Q��X.B������d)�MET+����xG���@�%x��A	��-XwE�tC�7��	���amnŘo��	�sg>8̣��s,�%�޲��OD򷞮�2�ɂ�=X�`E�UJgӦ�ڂb�w�h����\��t��R�v��1J��n�ͮ��}yTM�F��($F�H���	;s��d�̤�:���" _(��$��鯛��"e�r� ��q���~z�1�~/�G5�[�$�-�{�[��د���{e�%��l���NC;ca�g!"e$F�Ew��������*A����J���n�Z{J�r�