��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����Mڨ��˳0��`q�M�'���2&��Ȯ�W�4��д��|�6�K!b�'mY�`��L����T#�
���K�oj��eA�@�QL�i����K�H��X'��)d��)b��-�gt���x��~}��>�k�r��o	�l~SJ+f�-io�a�6E�@onޖ�4$-�Í7
P��(����#�'�LN����������(5@1ub��_���!�#��s�m�4�*!���� �Y-p���2�1����8�"ߙs�/��}d�)�`nI�b��8 �Z�S>!��Gqke����fz��"��Bf���5���I&�����2�e`(�2HU�k��ɸ�%�*�[ކ�#���p����6:��Fz������RݓO�Ҋ�mx]�/R�9�.b���~$݋=ҏ%D �z�5{�9f�@�6�GJC0jP��Y��0�1tF��A>51�2�|�=�0�[s�"W/ws!���I�A��ɑ����X��xף��Y΍��y�j�b����C��v���ֻC�,�ڿ��O����u�5̻#p	��]�qV������>��ߧ��7��S$�������������JP�G�V�����ʙF`��&���Fͣ`�
�x��32���w��Ϋ�Җ2�:��2�	l�Σv?�S�Do�X�[h1"UO��L���^���']��M��)Xyq?���L$��*�X&������Pp�[<��+2���z5�v�0����tmQ��!���V_�F��2�y���}ysB��}�mW�0^-0�6?�ϥB��F[�3H���?���iHƁ��@����2?S�%�:
�s��㫃��pS_�g�2"ɱ&Ɗ8���g?��u�t��M��l�̧�@��|ϴ�3-��8,��\����~[	eo\B�TQi�i����~�J���i*�3�f_�?u,����8�V��\$��!q�;ˬPa�)+��fv�ڬ��Q�y��(m���8v��ljEj9DVZp�%2]f,d|�Ԙ�q3�Ȥ&�& QW]M�G8�C̍��I.��)��ǉ��ˋ.T)�S��2�8��N�<�m��~0�a9-��$�z��Ε�W6۟�e�����}�SR�0V�r��n���t�֧u%^�AzȀ����W� S+�|T�ՑcA���礊�y�,�l'H�X��!���� ��S��ii�����z.�[���*b�<?��@B:oc	A�ޯK,��	}~�Z��Y����,f�à��D�W�C��sf��9�jQP֓�	B�Bdи* ��qT]�vS�a$
�5�&�8tW[�EDQ����m�\���~�5��-��6�hvy�6�F�b��i�*M�9vN2	���� ���z����`|wS8�"�+Fu��{W_�Qo��5_���V�Q�n�A�L�A���b9��#A!�Nb
���8qV9��ގ1�{6�d<r�5a�η\cQ��j�OFЊ��x`- ��Ɋ�K/����9�F�:��z:�����rr�e�Ǆ]���v*�7��`p�J^�=A�� jV<�LD�_V]�y�e1y�'�ڜ8��mÐ�޿u˅�?��]�hu� ��\Fh�z/�X
���8c{r�9�\�1�Ɠ"�\�R^_��ݫ�,1��o����$|>�G��ՐB�I|o���X��.�F��B������L�%�C{p��tSn���{�
�}p��"��b���'(_O�F��:k�ȩ��hs��^�࡙�
�6=�-ന$�,���8Bp��O`�JnHG�������^�KS�Y�&x�������Bs���"M�-������%TR8ҿ��p>� =u��n��q�{�ۋa���c%:�-P5��Gs��מ�V`U�>�`
4�_�?8a<}��9.(���y�+:��BX�ґ8)�q������3l[��1hS����Oy�5�� ��f�CA3^�xq�T@�O��Ҫ�#M��)^C�VN4��Aܟ�LO�	�8%v<^���k=08$Ep�V����sq�!���?��ki麇w)1��)1�Bb�%��X"�[�$�6B���g:����#߃��@����Ї�Y]):����>x�Q��������	�g6K���Ȇ��Qfp�DL��)��~3�]4j�E�}�5х(�|�.g�`N�ii�kBNN[ؘ�a.�e{��'�z���4C:���@0���?U�^�G�*Z����^���?�]���$Y��؂m���)_���k��^�E�G<�4L�c-x.�k9F��� �e s� �h�<�zjm��Sd����-�O&�������u����Yj�Q��D�Fbz .���3�]�q8�����V��>
m�}߁N����͒��e���7OSb�Lڏ�G�j-DR���������C�RӺX��}���V;"m�j#��A*g/8ܐ���僎�p���uYN��ŒU��#V�
Fk��h���e�o�	`g,n#�S�
���5e~�b:C�t��åIl�~��z�K�~����4�N�z�}�����>a��3����،ns�9x��4$�D����h �#1�=@�vzi�p�8���YE-wxCW&��Ί�.�a�PS�HߴqMž���ݮF�!Z�+%C���֦���	�dv�6�^�L��
��;y��i�l,۟p
,_�P���kg��j��E�R���24m?yU+�9�I���(�����)�*�Hh�
��R��8����7�.�e:��Ɖ�p��'�0�3���S9+�"wz��R�GK�>�{�<�oL5>��))���`���`3v� ヱ�V�
�G��0��"e�cU����2��pP�
�=Y��<�z�f. ͧ5�e�㵍��/_�m�N�S#I��Y�O=�l�SY�����8�����χ� ��lM*�ah��@7Zc��[0�jZ�^���U��0��p·�����d(��e?�����dH��:Y�դe��Z׺Q�|-V>�qI�#ܹ4�6�e��e8YWU�>����\�� v�����"���r0��]�˼�����;��iV��3e�E��J��<�]���y��.X��)�3s�4�^�7_��7ɠ;�Gb2�.��:`�l�'��f���暱]��9Z)Je�mU,����
!��8@,:!��[p�%JݐE�لE۾�\Hi�HSd����yO7T*�s�8Cu�\�7]>b�	h��I�Yd%>���eF��N�f�O"�@[�ӱ�5ܔ0�҉�0f	��'�)��2��e��Az"w�3#��'�i��?���6��x'6ğ2���� �O@��" Z��J�}x)�WP�Ê�ltvD�8��
a���r�R��f����%q&2C�TX������!��4y��uZ ��nH���l�}�1�t@	+�5�9ёvx�~JQ�!��SXq'��25�����@�SG��S[���tM���Vv��퍭%R�>�h�^��ܱ�Ht}�;��83����JG�+5@غ� ��-[D+r~S K?��[���o��'�c3�fC�L�Yw#{�76�u٪+���+����p'

څ���!?r�F�ĺ`���<���<�t��<=

 SYtSQ7>�Ɋ�wqհ�@�ՈA��"K%�Sp�5�_m��T�<b���4Ւ�˲@oh8����&n9@@M�0�.���N�-S����ʠ�l|���\L=Y(���r=x���W��#�"�54�U"֒_�_�JV�	�kڜ��=2�IJY�c ��T��܆�0�m؏�V���w��Cе�Zz�-��2��ϕ�����fѷ����5`�����}�|3ĥ������`|Fg_rg��_o�V���<Y�䜌����'#?R��*DJ}��u3��"���E��X�� *ʵ�\�
>���p??���IĴ=k$��@��A�Xgpk��*�9GI�VlY�H�)?�%Vڪ}��ǩ�N
:i�}�FÐ.��%��u��J���S,��~q�֐GQg7�~%vSD���mw�</-��^U0����/��u����ƛԢ��|���kFU*����G��V]��Cnr'N�KF87d<�6�vx�)����W���&yg�?.���P}���>��xS�V����~����"j�"�s�}�7��G�3
6`�5C���]ѽGha�^ y��G��1�,�>6
u������vŴ��Y�[��7ĭ��*Wp��",�a��ƔD+#k�-p��lw�}�d\n��q���s�J6�&yW!�I>0����1���hp�s=��m�"�*����Ir���"�zX�G� F����fu$L��2�w6�C��0IHn������)Q��h����ف΀�z��B"�l�`+�����r<Y��	����T���\�i������o	s*�c>���M��>�^l��zW�H�tBp��S� �e�%"���l!1�Yn*��[SG2Vg:_��ۛY�\q1�
4���nx58A��r����^����F�O��%��8]V;wAK����fE�/<��me�}$VL[����A��HW�z�P���#� ���B:c��qG��P�:�X��=i� �=*ȸ^�5*b�WC�8#Vc�wT�0��Uߎ&6I��{4���%Á�r�4IYb
��;��5)�y??�d�*���[YE[8��G�0IO�t��	Q%����8���DD��U�lz�7V��i�W"W��A��.�O~�����ռ+��:�M�~��\�KV<#zR���>8|��zk���5���:�'����hA)ǃa!/K�^�%�?��K�Hhga����>A/)���㺞�@a!�:j���@��� l��]���1��j0�.�����L벢q�1��8�U3��$���*;Ł�
l#
�Wx�l;/3�*F��v�8Ǌy�%r���4�����ob2'H���O���U�|�Ў�XRBZ*�L�a+_��7XO>e�Mm�~يyn{<�����>5�����nJ���W���2f�H���q�)���iWw��� ,���B�����5�?���1�S/��PI�+��K���g�ɜ����u��>�����v %؅(�mYL%���G�� ��P.�q�� 9Əѣ�W���S���Re��?���[Y�ik�������c%�uӦS����偣���JJײ��3�pa���KgY-&�a�$Wo�/3�u�p�0ͽ1��M(뗺
���*�_u��y�P����zq������Y��#>I֌h���|�2����I:3��'4�g��Q�o�tS��H�ݽl��0����r�>�[�W��^?�7k-k��"g۞�RMv)�ŵP��ǌ��T8��IlYq���zt{��V�}���+'��jC�qMC����f@L���r�4�t���Y8L�� �����3�})�/k*^
��=..�������ɮ/)3��h��$�8�Nu��Nxɾ�ly�>��M�ۉ$����Iԁ��������8��8p�ߞ���פQ��&M���r���K�ҷ�� J��� �J��ɤE��v�t'��s�"yϼ�?�TA`ޭ*�L�T`*i	��1�V)��[�
�T��sr�'��dF@���V�����ǰ �70�.�����6�q������6�bT~s�wr�4���!��� �$�z��ʒ��%�7{�}l���jI$�An��iG�F��c�h?�B_=Q�3i;����S|��_N��S��k����K���(�s�����r���}��:}��3���S9�x_53]M��zX���ѳ��t����#��8�g�;���؜��@)�)�cyρIb���nR�+�E�&�^��D����>\�����MU��;%9��D�i�,7�B�=e�^77�|��iQJ�ٺ�8}�2\Ľާ�(�ywؐ�	?r�щ�^�Y�W��d�̧Y�B�6\�iO�hH��8,�Q�� ��}���Sֻ߾�����`����"Zl�����5��Ԏ�����Ĵ�n���W�c|l�ٻP"�8ᔄ�u�|�#}	�h�Aʵ��?UCS��v��=,���j�0o ��@!i���3JY�k��@��#��;�qaH0c��1�w��\`��!}��� ?l;���|����5#����,D?/�&�+��%P���zyO��'��=��1_����V��+6�8��0!%n17|�=��ˀ`���r#��?4� �Q����>_f�+���F�c�_���&]���Yi�6���WM��+�P\3cm
�EF;��\2g���tL ֓��
�N}w����n3!��y��cOaj T/���K�ߊT���H.
T��x/�����A�H<��3-���ؔ5j1��:;���A�[��%�a�<%��$ro�m@Sb~ v
 㳇`�0KR�?�e�>���H������]�7ڕ�QҌv�a </7�>3xI 8K�o�<��T�����_1ܑ�sB$zشf7j��L?ŝ�`��$'�=P��_w�Y%����T5����vqOuoyPu ��PhK��x�Hp�ȘUۆq���X��r���:o���ذ�r� ��iB=�h��@Hs4z��7}`������.uv#�z�R��t�e΍�^��}ɴ��·]��p^��`�m�V`�BG/�����`���/���ш!���*+�bD���Pj��n�Ћ���Amy���J���Zi��Y���%����cv�����p���Āu]�h�c��
���	����qI�d�[e�����bomv�+��G�Q�:���kD	�p�㙭��4 �pΜH�[~����x�\V�&��Im��?�&�	�wYu�"�����N2��.~��9���(�#f	���:0�Y,U�������������4q���k�����&_��Õ�*v%O0��w���;��T�|��n�c����B�RB͔�Ɋ^�N���VZ