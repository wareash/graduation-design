��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,��.��̡�+P�FuX��d-��N��$%�I߽7>wN����u�]��j��ܹ�Ucל�|�=í[~��k�5�P�ؐ��T�5�����#�p"&�l�z�Fr&b6��,���Fԟx�ɅT2n�x��p����Xh	H���9�Ҿ�z�1�� dT�h6��[I�����B�?Oq�_2�9Ӑ@�p���G:26�[�6T%,&'�#JeR�+񸊎2�Դ��E�Jc�������5N�{�����Jz����+�:��G˦�<�_�	�'��k�Ov-��5l��|~+��,�Z��r(?�! WD_����J���K���םcE4��%2���qb�B^���p�G�A�t�\:Gȿ�B�o��Z�l�oS��/A�V�Et"�c|J��%��].l~0Ϋ�m����5u21sR9�?��]�q6�S^p3���ښ�=:Jm���W�����8lO�XR�tɠ�����;�Z�Y���j�f�ll�/����ɠ�����d��+Q�·�fT�ɬn�?�����V�L�!L�Mx>�4��:�!�t��*�㪯�Ҩ�1�P��{�i�x|�I�� NfпL���4��� ��H-L�dL�#f��Cb�^j\��-bS��|%?3�R��lVPy��&V�\-ՓR��pr�љ�#O%Js���l��&���s�<T�����5b���NL��4��l��� t_ĝ>�w�sw���y�fN�����@k�b0�&U��?�l�z�FYu�u����־S�wY�GBZ��SGH5GVB:�J<J����I^O��u�"��R�����$��[��NS���+*�E-$�3���%e���m'4�S"�6'i!8�L2"���S���!y��z'�Sxn�(���y��\���5�UǓ�
p��K1B�48��ÅaH�J)+레���-�7��by�&t\^�d����z�G���h��� �G�]�a��R~�έ7�tj�[b��QJ��֡=XlU�SA_��?��|Z"B�)#�`�K�ư���������?�(�l���(�z�L�,�K�&!��l]Zx�ug��B�L�u$Eq����L������HX��0N�����<f5�o* �'���K�/�ڎ.ֆpH�h�?�
�
A�r��DǜP��ODv�%��+��#��E��2��H�?pD�>Ə��F
�'�JM����q}  e-�����A֛�p|���NΎ
J�"Q���2*s�S��h��&t�ctU�ی��r*m�ƓF�ڙ�_ft~\�ߧ+�:���*�"A*����@�4r�i������ �I�J)T��f��~��enI��������0J��˵^٢���Of�Z���(y�_	d�c�s��v$�ji���K��aH����[�:diyw*���]�~#�z[ntѕ����Q���B�z&��j�ưA�����=����7
��(/�ʾ�r�y�x}K�5���G�y�+B��C�-Ƭ�<D�߼B�.��/S�Z�d��0
�����t��N� ��̀m�3�Dd�L������W�5��"�T�+�_k�m:|_ꊖ<(#��χ3^;����B�xǀ� �D|q�U1ѸhP�%�b�/�yRM[}i�Umpժ��0�l��}7�TD'����T�?��C>I�`�[V�!�R%+J;�L�u�@+� :�m�:4�h~	8��ɕi�H��<{�{"=P|��m����"75���B>E�N�mnjn�+�r&Goz>wW�ׇ�cy��NK�s=�*r�Z�2���Q����c$ ݆���D���.�A�n��ꆬ�U�q[ڹa������:�F��v0�졯��J��s��k!�-����	O�����tK!z7#+�㛦���=1���`�\(׊"l���=� ��lPe(�/�V*Vs�k[xF���5�����K�(t�6Џh[��o�$n�@�a�H@���޹��ٻ���y=Oʢg�q�>/�7b˂��Kr ��./��c_|�?���׾�u�]�Vi+� �0<y���2-<���pM�*	z��༯������yM&3ug�%{������t�`/��yF��������T��(��#H>;֘Q�L	����p)Օ�����Q�Y�{�Cͼ���R��ſ���n�7��w��Ώ?I��mBc�]���,�N��x�M3������ʒ*Z��d�瓸@��&��(�S>��(����^.@2��>䲢�?�o�;���5俬`̈�5��}bOrL��x��@m�ZS^?�b)
:y�L����csv i���2�c�B���xn��aܒ�uJ��$�$�I|�Υ;����\�`tړ��aη.��J�#�F��poM�������_��Oi�\�}-�����-F����'���}3����'H��m3u��x���J@/�I]t�GV�\n��N}ɇE����$�q]u�˿V\�=�捂ɀ