��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� ��<��T�@d�Gu�!�h�����j~���C��P�Rc���FfxXs�� PC��԰�O����p32iXA�t�"�Q��&?,P#̓�*eA�9T�x��0�8nVHAG8A��J	��c���G܂y��S7AC����&� �?�,�	�B�Ũ��aU�P�̧Θ꾸^�����\�(+��F�I�j�z	�Ϩ��y�g�8!�2���%Q���_�m�$�x���b3,B�6����9�@fZ{�G?֔H���R ���o�;��Hd�����������O��3�m.��]k<�B��I_"Z�L2��:*p:߶����aȈuJ�L�_&�݋�w�����j3�����:6���Ɋ=�����e������0|)
m�N�|[d�)��H���ڵE��Jq�)Tꗓ&�^`kC��O bC������h�j<��+�E�v�)��G�i�SN�p��x��Ǔ,�z1��@��t�ܕ돹S��Iເ��8�^x�)�=��V�fE�s��a�3c�e �ɢ5xE�'�fr&��W`��r�E�m�_R�W�(�|1��hR�%�O��p�ʼvkn��I���T;6�<���d�Gt����d��qkcR��H�5=�E�zD�YX�k���B��&+8�w�}��3V��Cbk�9G��3�����h���7�#���J���j���d�]�O�x�kk�J�1�A_��,�&�:�C����+S+�p�R�^4fN���U81�{^��_!�R�q�Da\��p��{��Ox�o��,ȕ����
J��wܡ�V �p~�P�l�}8���KP��שX���B֬ȼ���_�R_�?Pٷ�x��4TZU
�4E[vS���J(R�v��3��C
�d�5n<��"vݻ���Ъ�S~3�YA�E:m��p���o�JP�� ��"�!4�C��,���zO��F�/Aa}��]���b��km�;Bjg���T�+�#k)�s�̥��5�	c<���cv.����XM�ܸ#A����{��k��lJh��#S�[�i	�OO�DUx�h|W�]�7e��tX�%]]���ӵA�A�q�$?0������Uj4x��Q�Z�%'ݯF��v�P�m�j{�;+a���[w��7՝��oeCXq|���Xar�.B�ph�*��V������Pc|�7����ReN�ʴ�����Ώp�0:�&�i6�N�4J	�t!Gy��O�\�.
�Ҭ���{'%�"Ů�ihn{�+�����W��!�����C�d�Lf��zvˣ��!��Ֆ�k��ɤ�jd?�����Q�l���ҧ[�0G���r�fg>��֊��:�LZP�f����Q׸���s�oWB����RQ9�'uם�����i}�j.�W�
?�\��g�c5��ω�T�WB��y����\���۞��r�4'�όa��F�����C@��a�~QG�-4����no�%�~E�MV��!�R�M�O�_���˗ir�#j�s�q���2{Ǘʋ�>Y�����e��dHU��A�D��X�z��c���O�d�,
;���[�`��(��CCꝁ�C�e�d���@}ks���}F�M�6.mY1��p1���ӥs�Y'��V�_� G�VE?a5SC�Mj�����u��\aGq�^�5�V��Q$��-���T�1�u�m����������Z�glt!�<_s�����!����u�TT���I	�8头��)�t.5�%�8�Љ���P=�,��Vg)i��gź�$'_���Գ"|�X��^�,	��G,3e�:5��|5[�`9:��z�s�m�~��7����������Er��9�V�[��yf�J�x/������'��f{�B���H�:��������"���[@c�ݹ�Xˮ�[.���/�,ʆE��]�\�_1@�<>0h�t���&�ӑ2q����D"��C�������N��BFAZK|@�4g\��%h#@�N��ԞAr�cة�B<�a`����x�%��6�!�7���3�	o����!�w���0�lQC&e\�^�s���q�}���=)�����Y��qJ:���!R�)��9N�,j��rP@�nw��ȿ�1���\�� �����h��R@�z�ɆY"|������/)�L���ؿ�w���=��}���	ۑ$���[�0�S��`��=�����f]�98�������*<��2�ja�L�bL�	�E���zQU�K�'������4�^�.�FNJ>��o����5�b6��r���o�����Ne�FP��.�v�p��>�������`����:{I=�	�7E/���%H��PIwQr{��w�Dhܢ4xp��U�@�����81��EU��?�/���;4`�W�]��I_���Ϟ�z_��hxD��Sp��#�y{Щ����6Q�G吕��_�$9��`�E�p�4�(�m�.y���D�lڪb%�����#�g�9�]Dc�j}�*��eb]��׀j���ȴ�E�����
��&�Aּ��g��OU�ux�cL��~�y�&�MF�֧;��e�D�O�:�-��/K���tp-�G(�℺V����󪷝+�\X��z&0,Qm�e��@���ˍ����PcSc
���)�@��_s��1z�U��ݏ�s
Q"G��?��-�A�B�̽�~f}wlUh�{�F0��4jkj�0C|��4���U3
����׊;��;�	~�Z8�@�76ˌ��kbzCj�++���=�������_�C���ON�l�s�V!�å+��Q�����w��R[h�	�y�hpyz!�=;�)�BR���c5�'*V�!o�WD���2����2{:�X���Vm�hLb���ϐ���aը��p�T����8�U�	 ��No�j�%tx�.�ϸ���K~��H�娫�}�߈�^�vC�e��:@^�/e�cM;�j�p�����s�*:<I$>�1�-kE�p+�@rvS=Nd�A��j>@q*"V��Pu����E��̷s�Nd�b�x^�֬TB��`��u� �1_P	�-n��3$�H�$`q/������ZY�ڎ�܆Ǵ�}b������@��R��ꜿ�Cx�w�4���?�!_ ��[{�>r_�!��-Æ�l�T���h��-V�T�dN�]�:Bח��$���}��L�@����ۉz��N���S���6�71���)'[3����@c�͜bWN�ϑ8P!�5#*)��/�������D7�@_�7�����i������h�FV�O�3�ŉ����j�E���vW2a$�s:���#2�Ou1��đ�;H}��˦ʋ�y&x�c����ϔ��(e�!խ��6���KOgZ��G��P ��]k�p�Zį�[c	�<�K��&ߥJ�:e2j�1� Q �]q�`����"�LumSe��q�P+��1�/�ؼQr��s�ė|!WV�ܰ�7��A�� -ڈ����e�~.5��o	�^C�S����Pυ�"5�R���.cC� ���4�����VKc;��Ö����Lmڴ����#� ��ms'w߽fB�}���l��Y��W�q��IZ�7,�vG~�"��3X���z�x�k��i�qe�ur���~��5t�yz@��V�`������p�{j��!Ijv�z��2��REQ���״D����Ƹm�F)U���'{�����T<�y�=,�Fܵ�E�gU��Ph0�"h�hN-�N5�:��O��.Ð��w�VN�_FR-�gn����!]�Z��Ԫ�V����iu�Mҩ�aV�'��έ���GX��q��m�i�v�4
��$�i�9�܏�����i��,��y�T��e)�j3l�	$�U��'���s~��!Oy.:� ��"����1����r���Ye���^�e$���[j��NV��R�6�)��b��/�E5c���Z ��m���KR��Y�>��x��LG()Z��b�w���E�|�^�妃�a"�&�f���(ڎac�aW0F|-��ؤJ�$�I�,%����8vr��Ͷ|j.k^���I��"��Y�3*ϱ�.3��e��}�r#n�W9�M������/I^��;]cM�����P���b�k'�1eYӲ���L6����U`�{��Kg��������t#32<kC�t
e(��	�xȂO�]�4T�W��=07L��qv� �E�Es������ߴɱ�0}�T쬻ޚ����(b�(9x���ʌޤ�]7��1�F?%7JC����0�
��v2��UY*�c8?6��Ѓ��g��rIr���JΟ��Kf����,U"�-	�'��E���QÆ��͘�n*f�f�	D�p�n@�<|�^���8�.n���-1��# �]��>��Lո��Q�a9�i*�S����������@�UT�F̏�Y�K�(���b"��r�4S;cq7����g?���Ů��_4��+:]�a|��
�:���7-�AD���_���L����Sg�<|In�I�}�1P��$��c��ZN�ǹi> �+m(79T�w��節HCOz�����k�_����r�9��yA�pC�Kg���h����k�#v��"{��Ѿ|���*l皛��pIx{֑��s��i��8�?��ld��G�2�SX�Tr���'�@��Rm����ҧzn|�z��F�\���;�,ǎ�LX^�;���������dW���D@L[�7��nf�����&O�s�^hd����S�K���#�I��ىm��g�n���?A��W��#��bR'M�Y.�qrW�Lx3���	��g_�[��Oʭ�г�?ț��XW�v��M+>pJ��x�m�.����$6Q`��$�*6�����8��m�$8����ѩc��MP���Y�<n��FA�{k�xٛ�j͒�j��me,���6�t���p8�gl��d S�v@.j@��f}4O�$�~�'���ߏ��L�`[�r�o��P��kj\aX#��`��Yo�j�g�n�h�W��Dv1s��oǘ��5�>����jF�J)�Ҁ9�d�v<S�s+�;CkЖ*rJO��ώ�U��;H{ Ԛi�:��H����U���H�0�]1��:����<,�,E�%o?��n�5��`Xn�G)���J}s�������?��>�.<��hs�`Qq߈���x&���i�B�D_
nw�����cF���E��`ڊ��p��>h�*Fn7'�r+��|�9���G��D��x�������H�)h��C��zS�×V���;L�M]���y�=J�)o��P�GW�mhŘ	e�I�̾��b�N��,����6�v��ǉH��KӉW�*�E�O�F�`ȼ�=��gLM�^�h��]���ɨ���%jI ��ƥ�؂��wQ��tp�_�0�h|;	���Vd��3�J�K��lm^X��6���&Čr�Y�l#1�v�i�C/�H-c�A��{ߩ���K����gj����1�9�QV"N4�8-%M�2��|���W��C{,Z7~�^�ج>�@�[D	۔M����ȑ^-���[aU]�K����-������i��F
xh���,K�"����n?�����V����k��fSb�"��:�n��w����j%I-K~y�ufwlɘ�S��ܦف��ݯM����5e}x�����2�tL<'�n֘%�i���ǭa�����x�}+D|6 䉫l��3Y�y�0�kh�y�2��0�R��i�����݂)��0����8�R�\�d��3HD.��Ųg�P��R�u,��.(`�J_:��0{'�{.?����膢po�dI���M�j�{oX�?wRa���g�s<��`_�|��Ұ���Bw�E�+�mU�+/~B��C�M���o�d�� 0!&{��Ģ��?�_�Φ��9�ls��l� �sd�v�4p��4 $ș�o�!O��mV��L�$u�	{cVBGP�g����QMOz?OG�[@O��`YA�p�K������e<���U�k渣�D"�\��6Ԑ���\SQ���AG��]yHHSވ��ax=���������v��s�rM��Ys��W��zR�����ʝ�8d�Ŭxy�$�f��6'��co7^�"��e�����(Q|�����@yxd�;�UŧQ%�x�"����)�ZL���`�6N;_6/����zK��ܠL��xq���1�Y�08��C�o�t_4�[S{��|�x�Np���i:����FZgm�8�B\�E�[������gO%�
޵� �$�/������0Ӂ��Vz�X[�@j���O��FH�(dh0�'�I@fE��z���x/@@Q���2E�T�6i���#Vk���B�#�����	��aE�~�D��&$�^��ڿ�8���Ϧ�(m�̈�i�a���b0XsvBL+ĭ`õ��U�8��K���PG���,����oGqS?1&?V��,���dC1������m^�~ �pX�>�t��+��AZ��g���uj��u�(p�ד9��N��c�_�E��{����:{6_����cr!L0YtI	Ə�ѫ>U��d)��7cs�?�@�s:�̪��8Z�����0�
;��,���hL7�����
�լ��i	av��,/Ĉ�g�D�{@l#��yg ��[;�]�y����V��S�J����nvm��{�6��`��E�΅&�<o��맚�����2Z;]Q�	O`���E�:A�Laָ8��fhCr��F�9 ����C��NK��ǮT���ƙ�Q��Dɳ��b�Yx�-矅��e�;�<�WH5P�����rU�o��L�F*�uI��3�#�uʀ�Z{+�C��9��_#��iHd�O�]|��x�'閎q���V����yNC��;\w�Ǉ�ᷜ�ٌ��i2��8���ֈk ���촬��!Bb��}3���f���RẆ�c��W���,��-;��Lt�͈\�P:�5�̕��;��-�2��dH3�Nܚ��e�{tf�:W������ă!�4�[����Z<�� 1s1�=�U]ǣ�=~
b~�������+��
�-,08}�H���S�'�q�����?u��[��W�r %���M^���݃��k�"�����f����8Sn���/��^iZM�r�������%�h8��E��b�c�����[��t�ԏƟ'8�R����ⶭRT+3��>CG�0���h��JXI&Gt�w�:'������#���3�p��e*"�$��Ǉ��@�G��o�ۗ6]'Fb�P5��/�~T��=d���P��0�Sʁ����K�i�~zP�ϸ�,����}�ץ���" [�ŏ)�_ji����>$��u���.��L����)n&4�x� ���ҷ��N4?כ�s�:�f���\kV$ ��,u����	��<n�|�u���tLM��4�kW,��-��lӓ6�(q��U����S4^x�0*��0y|o���p*	<��!��e*׉d�����$z��p}'�������߷��H|I*��ʟ�X��⶟A��X-��>|��8/!�Q
��OH����o � ���"׽�[Z�ؠ(o���s[}�+$��~���u���n��<%V���=x���k���8��R�e��t:����,�}'T:NU�B�:�ѯVL�22 ��z:��x�fv(GC
���E��Pg-1���J�2:�9D���Z��M�.�>p�&$��Sυ|��F!:tn�{�9�������e�M̗�t���33������\�}�L>�P�:�*DS�)�f������lԹ�������i�<�R�b��z�"��R01GjV=��1�)2_�a�s��v����c��r�Mc{������`������)�m������s�#��4�|rͻ�I�@Y"�u�(HN��{=���������ۓ�G�>F���q��5�Ì5���I���%[\6���}n����ԡ�3$BD9ߐ{�vM�RRZ����`l5C}��Ie��W�3 ���6q,���3N5ދi��j���/�mi����V����
A(�� F���*�ǭ�X�l�5I�^MT�s]�(R��m���p�ͦ6�A�I����?�0-a����	:�2����&�J����K�4v�B���g�`�2���"mO]�S�����~*(�e�$�>�����i�����>[��k��f_�m��&����9* ��#�1�wqc\E�Y_��Fo���(
gD�Ə��ȿ]p��Ly"L`L2����Kr�P��W?���Y.�"��Q���<%�6E
���J�,��fȢ��ݫ�*�w�j1�4Os�5�il�v��4W��~�Bu��r[x�������)Qu�9�N�IȜ���ob�:���<(�U�P�Yg�U��)S˒Q4\����BG��^)\��0�k}��K�J�M}�{�������A8N2�%��|�3�CM¸8��(��V٨�<��-ξ�0ǫ�b^��X
4����'�zp�I�Td�t�>WR�I��(�^L�8@��"`ŧS����-�R$v�O܍�B�/삷a���u:�=�̹l�6E�I����ƪ��� LI�\��fN�{�G�����f�X9Pk�N�����1]h9�yz�JO�&�=E�G"/YzE�\q�a@�Er����mM�X]M�ä�=��\�}��hg�*�!D�)�,��g����qxW	�2�}t����#�gK�E�`r
'ҷ����V�z�Ǵ+�q冼�j������S�.:ְ�I���3�4Z�N�[ t��I>�0�nBp�6�i�d�04�۪_p+^����n��DA��U������<k|t�7QMx:v
��Os�l�D/�����hd�Q�Ts���pI�H���P�zX�w=a|T4�u[��L~}1�<���^��5"�D۰�snv�T=�� ��$i&�0��/'�V��\�h��N�Ĭ^��Od���<v��t�w�!�J�9�YY���H�:��&�j{��w��� i�R�}
*��פ=g%�Ñ7HcбY#�S�,�ȝ��"��U�����I}�Z����%m+?���{-�6MLȏh��
Y6�A7@�!�&���<*��eMP3�V]~'zs��+��J���J7���X�v��-ߘ�+�Բ]�8:�
��?>~XL�^T�/�n��T}���S��A+��tY0��k�����E�q����B<9�ڠF�Yn���֕�b7�1[m��4�p�*f���=ó��ys�nԈ�����Ak��B���s
���NBo�2c����+��陈`��������_�Ӆ�\�g�9*�]fś����n�q�E�"���)�{Ű��t��Ƣ��g㫅A�݄Uy�/
�X��G�C�s�>�SG���v.�X>��"r�6㱭�k��c��9���,�N�pw\Ch�6��4dՍ7���OS�طm��sɯ�:�+5D�����\���b{iv�T�Y�p�e�ysfr�x�}s�<N���XAF!M;ic���n=1T�h��L�����"���N��8�����ګo��7�)U�p���fG�;_甿��iӢr=S�����(2���C2Ԉ6=��Z�� �^���0�so��Lڠ�")l.�����RR-,�3L��=��5T�XH�{bj=��qY��҆b
n�/VP��
���� �9��*�	��^Dq.��7i�(k�l�XB��R��'��p��9�&v���qE����
X�ka0Z���zI�[���WC�� Z���a��O*��FH��V��I�WiWC�F���,��JfE��t����qѨ�r?=t��9���@���T�{N�3~�Z�_0�=E/�P��6���ʈ���ř�����1 ��f �n�10�ь�wl�[��}�襤��לG�@l�OG�`�$o�u���߮j��F���Xl����;��Z���7'�WW����r%���6�槌�cx��8���\d���P��5��A*�	1+��]X��������f��0��߻Ҡ�Ej��*����V;��x܀=g&M�/]6b�4Ċ͊�����oP�Q-> �����(-�����e������`�a�F��S,��5���"p������Y��Dn"@�Q(��xL[�߃�Y<�i��R��Ƶ1��er�m�N���d&U-nx��GK��W`�wYZBt��;ַ�s\m�+5Q�!K֭Gc���^�� 5˄�g<�H�O�'xè�j�4|���^�������K��s�>3pLs�7�k�M}�ݲ���d�bE�U��N�����3֟�
�����9�o�x�� 賣�0&���{�X0�"-��{�Gt��{�#'qk>���>l
UbkNW��b#Y�{`�����1�쫦�s"hxF7��x��pPfꚃ�ǭF	\�������	�FY=ʭ}��eT�������8�jOū��(�Յ�����z�L>�,0�5����% ?���P2ǟbBĝ%Y$T�09�h�W,XY��|٣Ǆ����q1�����h� {�٥n���#�V|#��G�j 3��R��LbGؔ�������o��}����ޱ2���R�ļ�3P<%z��>��Ҵ�h�%҅�������>u�xϢ��uPzI�4	�U�b�j�zZ��k���of�R�?�0��io� B=1�%v�A� y��+l{���Q+�L������Fa�� ͠9h �.�v�_�d��C������Cz	tEx3��9�+�l��[�u��B=��+�b�������<�h��pOA����>QGw܋VHѭ�IQx�z��N��T��r�L�� A��~K���ȝ���ܼ��6�.�s��xN_�q�[��{gt�iN��3�z���=�=��iQ o%��~d�9�b~��&`��\�>���7�tk�CQ�yn�#mDas�'��u���c*B�3N�b��$��I�_��S�].�ܔ�v��+�}��!�":TbR<'G_�lk�����
;1��:G����,���dx��j�}�-n)TqJ2�G-�~��f%:,�,Ѽ�c�I���)ʎ�U,p�z�,�c�ƌ&�x�fգ�a��n�
�F�*v��FP�KY��i���
��q~$��7�s)���п(�eh}@|M@�\߶M>�!�#+�M\�)�zųVE�+��Vdo`�9".dn��!w�)����Aᵽ~�=���}D�,=�.��=N�ˣnT�hy��%���g�XՁK��{K��eA�}�RϤR�;�v��Fe�NR��ke Ш�>�b�~8�b`9�p�S1���VY�r�:�ɱ�����"��1Gsry���I�Yb�) ���"�$L5V�y� m�ڪR, '+GU��:��p���?t�=��/�
�#�����D�N��T=rn#x4$�G���{���G:����l����tB��G2tB��!�~�)44�o�\�X��]V�H���54 �g��I�E����D�&]/��|[ʔ�ȥ��˘;\e_��X���cT�5����`r��:���:w��t�X�����R>TC���kv�D�A�Wu]�qǵ�9����l�isY�%�����g���Jkb����^��As~`C��o~�.X�?��5ۼ[����Ӱ���Y����p�������y���R������Td���c�ّ �皸�" �w:]?�oꢩ�0��gZ� `]�~�*m��HPH
�I�r�:pb7E�C�5�v��b�ȉ�B�T�#8{�l�w�f7e��_�$ɒ���ј6+]E��OM� cR�%�	 ��oGt���T�$�ik;���	�����RU�q9/�ٶ�� X�r8����	mp?�#b���/�GG�,gv�Q']����U{��Wic��Y���%>��h�y�����dgL�8�����l���s�]#Ʒp������ �lץ�{�jұ%}�	cAFcd��������N��&r�ZN�H�WD�	��i���J6 ���8J�xF�V��a�Su��Ů���*8�NI#�x���p�G,�r�+���ϕ+O���`<j���CX���]����Ʊ��+�Nڈ��*&-
R���㭵�\jo︈���e.����8k�
��w�LG#ܘ�t��)���ٴ��c`o���m� U��o"`-��|�nN�0�`�u@�r��J'�K�}�U/�#r:�AP�G�᠈X�-1�)9�˕3������hID*��9;rHESP�@<�q���R����֜�LH
�96X!�k��A,g�2���w1���h<��2Έ��{��"�)gϴ=[���|bzq�|�#��1*G��C�#�0@$�E4ݥB&��7�wV>�n�c�w�:ɱ5����j�'�F!�����&�u~}T��v�����G��6�y�E��Y�)�����B�5�4U��}t駰�Q��g��n��MC����|x.�@��˖5@V`���TEfΰwT�H�f�<ї�d!gЀZ�?�e8��Ԛ��v� �������a���Ǟ�g��=P�����~˰>�zS���JDH�����$��>�e�6톈Y�f���4vi�����4��7E�NJ��F �q����_0?�$Q�s�}L`���Zx�lGw�fee~2�Gn�j��Ղ�m���A������R��;&i�0 07x*����s�zgO���>eVH�Րg���Ĉ �0�J�,-Lm����qLX���ڎz�g�*��Y��E��#�����+|����ٽ,p3c�3�ܮɦ�W�����ckū�{9έߗ�UU�A[b���u`c0��!��?�ϣ�ˣ$�~ ����
x�F~	�P*�c��Zl�~|V���=��O9�	�li�U�Q�����g\L3x$?�%e�q�>�	���ʅk�χ���Z{�h�� ��G�V|�)��b�����3�x��#�CN��)	~}��s���?�=9-=��E ޒ��EYG���MqF������N�[���8��n�m0�Q��q������a��,9)qcw�Ζ��
�\�Wq�a���Ba��y���#̣�ɑ�E�#�����n_�h>����%4I;T�zev�{���{�
��)1\"Lʟ�����S��k�C����jb)vVH~���4���-L�����~���s���3�p�I{�D�z��}'�(�S�#�/�r�ro�V�����4��u��譢�����]�!���a�*5�H(��F�g4��1�=R�F0�#�O-g��  ��T,�L@�7;Q�鳘A�@�_�a��ڇF��8��Jd1�^A��#AІ'�����\��F�V��F�Q� �L��QNFdM���82L)˰��w2���V�	`�K:�/���e�M���<�C.<�5bF:���J@�y-œ���	�BOᕯ��c���ٟuR���.���=/})\��ߟ2C�®a4��еc�s�:dG�>JY#��͈�%��lry=��������hH�=�"
[�ʗ&(���[׬19�̫�d`�`
�JUlvbJ9ǆ����E�wT�[��腌)|#�R�E3��R���� {Z�ӜgH��������R�f��I�]@��ʄ��M�����O�m&�E{C�ukS�;bf�_��^�v�������p*溙T#f��_ذTx�E�ɍ�mg�U���j�D�@"a0��?=\p8�i���X[���w��Di�4E���ue��V�VC�� �XG1��|���8�WZ`^6l��a3zA0Z�ړ	��$/L���i�1u��s.�A�cW��x!r�� SIJ�LL(k��:��$p��g�:��>�@���X�<{�c�-Quߘ��Y��j��Y!��Pl�(�
%d�o�8���e�}�W=$:>۸��
�#�?�˫O�P�����|�@�������pȕ�ZڗzK�Ԩ~��������Lt�����
��f����#��y6��(���|� ]�<2J-���+<Z�8���:�5�Z�kef�[�����1[(�G�%��h�~�W���-Ќ�d����$��2��i�����n�5i{��#ݣO� ��YMG$�a(#�UΎ�.h/(o��Bkp��!��W�.�z�V��إw"�����^��d�m�3	b`��H�i:w~�z�޶[�tj�X�Cb�3FF�#~���
Za\7�ʀ�gc>�~Ƅ�5��SQNf��+��۟����i���/�r�9��ɯc��^�H�����E�]VH�$�@�/X�)@��H_�X�gѝ�hJf�7�U@_�%���H&<i \��e�����p�2�mw��N�� :��H�K�>1��~�f�h����9Wy@�xl,ȥ.�w@#VBR����fs;t; ����y-��X@����W>}hv����IGVҾ(1"���7�W�q��Vr<�\�b���t���r;�b#zQ"!v;� ݧ�5+?�t��[�#����%I� ԯ��z�xࢀ$�w5/�ꭢU��R8쏓�����D�O�B�h>�©\��6�0�m�ݹ��w���6 ���4�1�g�b7�ѳx�"�lu(���p����0�L���,42�v��
����9S������*��"��Tra�BR����be�x�T]	�zJ�d��ׁ7q_��;��!�X|MTp��t�ߒB�Rna�L7.�Dt�o�]@0�Ms�*�2���&�Ϯ��q6>8
>TWu��b�܌��@��ɤ�H��v�jS�;ʩ"a�<w��)y�O^{�7}� ~�Dq��ɿ�#��_�;k�K� z0����Z�LL̀v9��?��lExm5�uB����;Y63�(X�`�Or�?���"��j *:��y��� y�����!C���2m������/��;���-�}��O(t`�m_�O�L�W�H���\��2�Ƃ:{j,��<x�"8�"�ǘ��E[�$����Vw�`U��.< i�%�Kz��L�x��9�}���[<�ߠSz��u�oܺj���9Z� ���t���Z���	���1 ��og;eA��Qx�;¢�����H��W��Ϳ��Ar���X6��T�<�U��n���-#D�P��<P���&�Ik��#�n��$>4�ƹ;*]^����*�y�'�W'K���� 4��Me4�`�♘cR�S|�%��/f��R����)�%��M{H��k�����{h1�����R�KUt,�^r�6l:�-x���V�� 5�>�WXOT��k{g� �꨿����'-�tG���_Id]��)�4�p1�L�,���qu���j��� on�R/�����L&���(-9��KU�y���&���+=���V�-2��ko;-�8o���o���@:5Ry�	M�f�#5f����,��BB�k� 4�G���L���0����5{�H�d������m�i�_07!��ć�.����a�/���(�B'����A��2�Ļ�v�����(����Z�I�02�hX�b�P��E���4d�/hq�N��������:��?���L �[��s1Q��v�p�� �F�_��7V�!� ��<[ҼsN߇�w��fe��}���5=La#��=��n~�2���U#�n`�ݾծ�g0_w�/�F|v`Y:U��T!�y�-�$���
��UעAUK��l(�soװ�+��2����3j�2�xk��,����~���.�$�x�g�U�-��(��`D�f^2B���f|Mh�u�F�&�m�[���}���\��v�����Lk��9U�Y>�[u�jqv$��mA�;+-*A߯�J�������Yj�G��BWqao�6ߺ"*F�(P��l�{]Bo>�i+!�I��Yݯ�
�e��{��=�HE��ݏЙ�LQԓ���y�(\X����%���nL?]�_.R��U��`md��`ߚ]�ש�ǭx��!�иT��ќ�q��PB%E�vR�8��L��Q��Lݽ/�,㑬�e�F<[�!��FH>^���h��e:x��*K�>1���/'"$�?G�X�|�)���#�=c}i���t��(K �Q�R�RZ��n�&�N� �z�x^CI|�lP�ex �r�_�i�5�'5������SP܉�Ս�_���=ta���K�+#���3�r���pfc��7�['��&��	^Y�(�c�)f?�qHo��q}��K��C���B��S��1ʦ����Ё��Z���נ>0w����zE�[�M�J+0��	P,���{��@>J�8���w7���<Q�<5��3��`������8hE�C� XA��us�M�@���dO��Ml����+Z����u|��B�P�By�0�|�=m��AF�ޞW�D]�����Q�=<i��R`��4���&��Z�IDJ��#9�qICf��?yT�5����.��E�n!�,��LߝꇊzY�W�7�'<��	 ����Q���n�>��J�,*OI�2)U�4,g�Q��؜(/��l~x�#��4��2��71e�&X�fz^�-C�����!?�Lh@��������خ�B��p�U������c� !r�h�A�d��5��ҷ2+m_�# ���o>d��y{��U�ċ/T�EϬcL�2ܶ��+=\��%�?��t��

���4[%�;\P%)���̒YZ(�Anx�ߌ+4��3�d\S&�� ��H��"T��cJ�Y��z���o6uw��nm\�����	�m -Ζ}���א;�!?�4 ,ehܣ� OVr!pN{L����X`�{�=���g���㭧&�B��h�k��Y�H�gUH��m������Z�B��	歾e\�kK�>g���/��[��!ZMҶ �C(v|�S�)���)��M}V:k�v���U�c�f
�_!�B�s�]��)�xn3�C ��v�.�$> XU��>t�7�W�F3��@�O87�Dc����u�_-�!S�m�~�Ǝޅ���a����wҌ��롡�2�f��w�/uU+v�?�R]p+_���R�x���&@mk��=�+�l�U��Ak��q�1����Aw����;�,nBR}��ƕ׸>(7�F7�[~N	�[BSt:�%��8�H&����]Jf�g�\���<�z~��:; �i��kp�^z�a�u��u�_rQG�T�9�مM��W
)��7b�XB��}�	����)6�~� Ҙ�vF|]����WMKY�d�n��,1h�;s�uv�Csm��Tԋf]���q���5Rl<ݪ*,�9_�=�),��5�I���乹���mͦ���M�0e�\x?@[�-U�e���� _�O{����!*��"g直rV���� ��B]s;5D�,3ooT�d)���A
�y�9sE�u�E�z�(�1�0�}�
��/�X_��?���/�L�T��"���h�5&�J����@b�N/P$�s��} Jf)y��ʷ�#C���4%��~��0 ����s/l�3��JW�xzƫJ:/�R�~P.	�BٳJ�WT��ޡ'ࡸ��B��7��?���y,վԊ0����&��XT(�#���gq�M�[#|��6C5v����`q#
�����z�+��Z��籧����Ɵ�rL�2-��� b��݅;��a�#X������8҃��Q�tv�~2uD)_��0Y��@��+�ܱ)����wہk���U��h��˿��%�Ô"�fV��z*~�H��G��kh�п��6�b/�������ޫ���4�:kc!�����sf�S��3d��f�+==O�ꅴ_�/^�dd�+^t�>c-S�cN��X^�+9�M2Y�쮡j!���E4�P�ҽT��(7�>�ֹu%���9TMF���Z����
��GyVk����b�U�0�C�Mzv��M��7{��2⶞<���I�.��?���67�j��[w�S���SR;'ɩ�,��x�4t���kv��D������U���n�j������Xb��X�~��	��\�� 扺b��[|���,�E���>rDmݭ*��6M�ђ�x�-}��Nu�E�V\��ԍ0lEIO�0JH�9�����(�K��2�ڤ�&Z�!I�b˖��>�D,���^%$dw)�����E������z/�� Io�j}����ܞ'�E�^_C��\��	���hIa&g�"��+fzW^^\>1��>9
J�$����k����LӍ�.���gj�� �{S�n�LF��]�\������u���X!�aP��G�'YO�<rE:d��tm���?�ٮ,WȚ���χ!'�T��<�������!]z�Kė�r�^v28�� k㢳�*aM�K7� ��)�3�V� Vb2����v��a���DMW�k�u�ɂ��!��'��aD�f.=Dy1����H�أ݇��?$��ȱOy�0��.ayZ��-�|/ç���������
�p���d[UqЌ):	�CTWk��ڦ������@j�n��ʀ��P��0>�����M%<j�G^z3r�]�-H$fd�)��{�á�G!�d�ؿa����|
�lK��o�R���$�h=�u�η���rR0�ne�.#?�c����Aℱ3�t�qs��i=������fFB��bm�>榺�?a�\/��_�,���x��ʧ5Ù<�ܭ@��V����G�(�h�Y,F�VjVfO(��<n6��F�+>��z��|�g�̮�Z�g%]�Bo����q)�(�w.�a��IQ�T��r��υ��46�ܧ�ꗠ��M�+֊���{��\X� #�4�K����R���#
�</��u�� ���_�w�z�1�q �nud5������/[%r5'T�S�cN�ϵ�D����!2��U�,�f�˜Ū���}�,��������DU�T��W�s��=�OsuUܹ�۠sD1
rM)�P��~��F�TȖ�V2��"}��]?~���g���k��@n�Ay��A�`~4?<u�q�(�"6��H��O�2""mpv%"e��T�R�����"��p^#@���u�X@�Иv[���P�b#}��<l�_������^.��|�-%'��5)3�u�+���X����� ؼz{����x�����+6PL�5zb�U��G������I�S|,�����R�K���ݮ��H-�};���;}{(�pｅ8-!��wh���,�� �A*�"��!	̡��2:R3�D�V�_*f�9�����CdN���ߵ�~U�2�lA�Cx}^)���}`-�Łj��u�o��:��أ�]PS��kO7���Srd)���f`��T�*�J��$�#��n��&@� r����I[!)��4T�iJ�D&�N��4�b�8�8��O����p\�]����f�u�W1'_����w���^����&�5�x-o��l�S"l.�|T։F���K��VF(?s�	%f,h_-j'C_߼H�����4�-q��
Ǳ��+�(,ʟ'���fC3�M�ؿ��%������f�������ײ8z�)������a_BM��w
�b.��}+Ju�卄�
�_�y#0Y�]!��/z�������T�����q�R� Zl�f0��*�H~H2�����}F�`̤l�"0�I��a�S$'צR�f1A��a����6]�ł�gO�f�)T߻	6���	����`�nܬ��e�,7�g�1zs�m #�tk�o�g1=�