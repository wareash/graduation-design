��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� ;l�Fv1�ϯq׆������s@���'����j����դ�P:�Cb�{�'�t�ɟ�>��(Hw-�u�� !i�^lZ��C�{��И���i�-|�|�I�Dd#����i��	�4�@$,d�������v=�3�A�pO�w�tE���M�ȼ{;��?4P:ٮ�7���F�ڦ� w0=L+=~�&P0q[��^�-\ߛw�T��e�z�"�[S��B=q��È��A7�D��]�!Tl�f�+K������<d��\�毙�����gpȷX[���;ފ@n�%%�WNr5��X�hqҶ�=PY�0��WΈ>��uX�+4 ʿ =�������5�i	��,�Hɴ���d��h�(P�pFtk_���'E.ݷ�T�q����l!�&˃S*��, �FȽ�'(�k���=J�?�>:̃�7�\���9����Px%[�C��a�d�%�}�qyh�!�ۍG��x�58��Θ�|l�zFSg�\j=)霃��f��L�U��!�@C(����U>�RRrT� ���X(�A�G���I?�/�I��"�?�Z��E�T�w>�3p�>����G�FJ`Eޑ^��&z9P4��,�N���*�
;�˰d~4�� ��'�L�͛�e��ث
|%��QLZ��s����9[S��ʝ��:W�7��������gG�^:�6���3=x;-��;
�
��_a���-�V�,+Z���N�69"|����a��tZ>�G�.�/�2�7]�Mg�S@~_m����7�ZҫӁ(�,�	2?���G\�^�����c,Sʴ� ���F�g�\OA6��-+���L�����**l�K��:H�\��B��r�A8��ѵ��1M jp��x���?S��p�k��ʷ8ώsr>!w�2�O���q'y,�g{"�b���ipD�L���#2d��!��K��VFha��_�
]{P���(���*8����N}��^�g�VALl�j�ߖ����6��Ff�'�<=����N3����
�� C3���� K�z�K��^�q�a#�~�F��
�#���xuԇ�#�k��V��z�'�.�����簸�NJ9���ؚ&[�����̀�!�g��j�a�v3��7V�_b� �u��4؉R��c�A�:�$]�h,�~�w�Vh+���%h�R'�4�s��ո��r��>����x�z;�3�@+����=�I�!�";�s�/�_�V[?偠F�������F��6�&y)Z��u���%i�S}�Z�R�"���տ���i�����޹v�]�f|3H\)�"'�)�?�q0,Ct	V����'�C*p4�վ�r�n8�d����V��|� ����M˸"	�%Z�CD���F���]���?��[G�3;H�m����kN*ؙο9Ɠ�B�� ��G��a�c&(�g��L�u2��i4f���8�e��Y*桾o�E&�`�G����"G.���w���9���yZ�?�v�{d6�����؇<�E�?�4�x����Z<�n��~qC��[V�	��N�~�9�X�,����-ˑGC>\�ML������7���c�;�ʤ;5 r�p�Z���41�3����4����	��R'x���������οe�+a�J�=���n6>VU ��2rJұ�x:�#���ojc��0�:�8c�|=k�g��	.OjI��0m'!��<�f2�>�����\F��	��3� �\�����-k�5�y���J�Y�/oV�7�!���;���*l���hO"��v�#�Xf��={����/?��8�
���-�ߧ1�+��xK�����b>ٹ�.e��͏7����s+d7�-:���|5ʁ�����<�ro<�<.|��h��*K�Gɧ��[F�j6�Տ�?�/�o�ͥ��!����C���*��F��(�b����µ�Ta�K�ϟi-�O󥍑�x��BYj��E���CEw"��sB�H��\ �����i�g�0�iV�}Bh.�DR� p�-��	L�T��>����C��Nܭ~Th�|��ȆCY�V�����o���qn ���[�_@f���P(��B\��QW;y��Dc���d8d�9$
��CC~����+����}V#ɐ�'�Rb� �"<03E�vpE=�~����M>*�8\K^A���9S�R���a
r ��dds�]s�al�0�C�,�X���*�R5��I�j��[[-�3"4�Ju�?��"uQޯM)/�#&Y�w���?��zx�j1�~h$mB��{�݊�����D�􍣄�B�4-ٞ%jž9Vb���xw[���q���{yja����18sk4�b�#v�0�M0Q�Z(����,Y����À��δ2+�=RJH��
�������s4>e���}��۫� �@Z�rJcV�)B���ŦG�D˗ch���u��Gv�`�@��ڟ�O��37�����I�f�!��1CW�t�%n
������z��vб͊�S���~Q�~
�ڟoX�LƘ�֜�`�����V�Į�J�@�|$ņWM�6S���Lkw��4���������H�cIq����Dꏂ_ذ���x�����F��7��jP\��lBg菻�"?���Vk�[q~R�3o5O�]K��K�_Z/lc#�n�9mRf�����;Z:���`���x;`+fV*G�14j��/�)��ʈ�T�)~���NR_Yª_orױ�B����yפ��"g���)�7tx?r�����x=�zNVo��=Pބ�ou)t�@��j�׳�~�a]��:sbg�� �;�q����gmG�zh�1b��n.W
�v��%�� �&���+Y{~^�t3��4�8���sU�V&���{�����qc2�dw;��鉳�ې���w��tQsub`uAA�-( �]��U��J��SzU/ӹ�X���W�@hg.-Z��d�CH�@�S2E�\�퇃��X*eri�e�M�WL�؀���{_���LH��	6��~<\�@�������'�5��K�cM2!R̺(Gb���<] q�����M��i;�e��zq��:��j,q1����!I���5�5��Ɉ�:e<�LG�p��	��s>�je3�J�MD]��Q�������{��@05E�5�xN���,�>�Y�t�	�³nb���j��=?J�KBJQݽ�Tm����?����g2��`��S��抵Kф��g3�nr�*�+���Zz�eh[�AڡZ��|pp���Ƈ'���TS�� ��P�7$CI�e	��-��. I*��,l�1"
�M5�^���y��Z�ۙ�i�MO��kN���-Z�K<V��S@�w��
&C�F_u�}}z������/"��:)�r1 X��b��vd1+�ސFhf�^2�م�����vC7ö��Cž7����hz=��翰�ח/�ћc��Q��8�Q]����0�U��r��ġ��J^
���hO�lX�)����5��J=�O[%V:�Xn�;�����x�Q��Ɂ�=�Cr�?�gH���@!F44~�h+�4gܺ�>5��CU��Ly��S���X_��9��=�a:ºiw`���_P)4V��H˔M�AXD?��D<o���}S�tE-��
�L�kZ$�% 2�~�٤��xM�n��.@@�܄�N��z��)�:��7��t���@�5�!�$�����i
�C�#��Wv����3�jEA�<��.tҧ�}T�DD3f~��ݦ�x����%���� "\�gh{��hk�V�XA��lb���G\�K��<D���|m�|��aw�~��#���C�S*zP6���+�@�ЙY�lh��e#�M�z���X�Â��2j�
O���s�J*:��D	�NNb�����j��4�?k��8yӫ��U�x�z ���'Y��o�R$ d��b���=��mS����js)�'���a����w�^����8sQ�� �5*>�J�����l��uM���4䎣��r{�8���8�u�����F�Z΂��H5������1��j��s碶q�`����j�f�C)�����,S�w���
�kρ���\E�SIe�^��9b|Ξ`<6�A���Ě������E@�f���ۊ�% ����=��"|�PF��	�=T��GW禮��H��S�k�����i�o���H��M���F��Gat|$�!�zUe�E�t%����4o�4�5weqiZ��1p��[ ��^`�_s>i�-�4ְ�&��nS���~�_��o���8�Dա�����<�[����]&���[��E?�xc��N7m�U
{�54Nn���Ȱ�B��Q�!1�xmH-����� ����X(��성I����xє5���k����@�X�T%�+u�g)p�"�Oy�Li#ƶ�w���#k�\%����рs�?l��`�V��ey	eE�ܠ��M;�{�S���EM1��nߢ��!H?��#P�ZpK*��\�-��UE�����F!�Nh4����+Ҹ4�W��'W��$�I[�)��L���@9�]\�z��"1�N
1 ԡ����UT�-��� �}���m���&|��|ăN�vC�[�7
:���	6���#��4݃D#��r���eދ�g���j�R]2F˒�%E�}	�J���X�wUM���@�=P���1�x�>�SpM0�Z_���ǝ��)�d�3�Z���5N���jF���A)�����D��F�tɪPc�f�b����1e�P.��(^���G0����6�Vf�2��s�:Uq26ӽ��EA��"�W��{���rؾ�мq����u�1'���㬸z����]+p ��=�����跰���g$�A��*=C�%��ǭƍgq�F �E�$��'p���+�	�ͪ�RՆ������Tih2�.�%`�6����za$�f�f:� ��\�^s�+�xnYf�!�9�a~=�/�*ES��*���?�R�^��(4����D�o��M�o$gms�j�_�j�o6
3+&�l�����ΎhGiz�.���!"�o�;���vRJ;$�v�׳�yQ����ks^��bD�yK��-�ˌI[�a��l��P'��9�,9!Ӻ<w6).��%���H���|��u[z�`�36���m&|�/È���qt��P���>߮姹<��E�Ɣ<k/zX&cD�~��cХ�������2��4i/ž�Б0+�K�c�����M�K�f̖�+��-a~.�t$��eb%����{Sh�T��F0o���.S�t	?~��錀bO�=��)EyW�-�W��
M����)�5j�hm��e�I�@����~�?��k�N�u�k��;RT4o�U5&���e(y�fś�S:�8�Q�����Y�%q'7j7W+9���|~�n/�B z#w[�;(|e�j��٧��������+H���瘭"E領���F���;��-DU����3dI����Tx�&��ϧ(��?���W��:��<z%!I$�խ̠W�N[fW�s�v :rš��:Y���(���ΰ�.�b��B����X�!>ؗᢥ�ص0�^��ˑ���i=��t"��u u�C�l���J&4�&�d�U-m��֍�)r3]4K�v^�m}�L*	�^h�E�����4�-�b/�h�ٴP_��4��|<�b��/Eܩ��2��K;���bP۷��$�:k �FS�bY����mJLc�LIRe�^T�ʰ9�ߴ`�i�ǡIˮ��TŁ`U���u�W�cxG�.^�DH������<���l1⠵�a��|������:ٝ߳�%�9��g�.L�W�E:L=ZVҶi&� ��S�u���)]��,�v8�Z���6I���QW5^>Q���g2�R�H*l���M�it'7#��y^����mxץ�)����$�����Qb�{�'���)���E�3B���A5��4Ib�X��pg}�;k+6mB�H
�ruq�u��ޅbl��kW�+n��9jYBc�M��:��o+��<����gE����Z4�
@���Z�Խ}�����廎kH����j��s�K�=)��U�)��VBq���ՙ��!�3؝A��k��������)��fk��E��z%U���X^�Ei�1)�ח��'B�j'ƹ�bh��!�\�u���Ǉ]$���Qҵ���]�T�8�;���c��Z2����h:6Ⱥ
�.�"���BG�#*�F�>��JT�3��������=�D��s!�j�'o�������:l�v���)$2�S+fqj �]k���e+���sF�!�Rhx ��A)H�7�d��|�=�4��]�e�"��p�m�%D�b��&��](>K���6��{\��&�]ބ�wD�
;��E��Y���J��މ~�곩;�5qz�T�:�V���Br���Іl8z��`ů[|Aܱ��#_���{1(��x,v��k����o��d\�a��~E�.�\�E�^�B�#�+~���7b4���Ģ��W?Q�f�Y�w@�D/�N��j��d;pG�p�#d��16��lރI'�/�ߟ,��?��oz��ax��.��;1�6�6*�[�����b9 kk��]���l��L�'�~���3�p�\�]�dD�|#�G�ҥ\�L�]��q)]���,� �l,��.Β'xу|��j�$B
�̂�R?���疟B�ٲ����Ω�P�>���X����w�#cc�C� �e�������U�����D�BmPl8	�U޳v�G�$�ظ�Kg��ƪj�w�����>^q����Nr�[dM}3�f@V�z0�K���Y2^�&���l,-�/���;`���5�����O�e���ep�X�2�g�]ym���vj��#��_�#V!��N�DMלH`iC�1F^M�U�ms�'M\�G'�Zf)�y4��RJ�`��pޅ�y�NB(�d��L "�DY���(tZ����y(�eH�k� �ؗ���`�"G����*ӥ ��ϡ��E���͛�h�q�S +y\3O��'���`�5�=l�-�wvpC/��\�*�#�`5�r�����~��/z��U��Y2��f���׭��V�r�%ݞZ9y~����&m{?
�8�BL�'mҙZ��Q��"���q�T,R�������MBj����b�k#k�G�Y�8��7Z�py�n���/�;����;/�-2��3���
i�pe�=�d}�k�,���In��#�,(�ɣyI��Y�6s�x���.�U�q��i��Hɉ���c�5�b�OC���5dC�R;�`6�S��kvl�%9�8�k�Z�Ћd�v�!a

�&)�qt;���&ZGOg�jZ�po#�K�	��˚s�6� �Y&j�{sipM��H|<$��$���[�7�Y����m�	GfL�{�
4Ò��߁<���W;���wK�lx�,��m��~� ࣹ�gƅ�ֲ��f�{u�W���l�m������Dg��\������]�TQ�U��ѪF�6�{	pb�䚈���P�9P��d�Ր�q��x�L�Ҧ� $�0�r��Gf��rAjd'P�u�3�S'`���x�Q�n�P���Ml"�R�Yf^���ȫ�%@p��xޘyy�b����3�V�>��K7h�T��(T,�WII�q� o>BV/d4;1��a��"�@�ü���=���:�_����{�_;��ޖ@ʾ��N�J�M�@TZmF��\I��,��vc$�t��}kw�*(�r3u��r���Э�<]D���Q�k�CN%k�y̑�5��^�`�Qs4ߴ�|�w��]�A�ΦF��E���.����r�2Yk[��^w~Eˮ�x���C�v�+�	�U*������@YO+���웭�u�q}�݋.AUK�,�h��jN�% ��	GZ�v&L��.�#ÝZ@%�x��|D
"�����P�����xi^SO��ߧ��z�/��푙�w�2e�+�ֵ��}0���a� Č��b��*��N��ϳ��п0��S�q&�]ʑY��K�����[o��u�|gtp0Fm!�\�+�a^2���_���]Ym�����l"5K�6�0�@}	+�����Wdآn�����:�vSs6f�%���������A��K�q���ѳ!�p��5C[�e�2�y�Ď��F�^|����O�n�LZ^c�>H=�ޑ�dͼ�x$v(f��,2�H!�sQ2r��6���b�mwLy*�?��[:-0_[d���+A���Of��֊,��-)rh����ԁ�Z�;U�a��^d�t�	u����{ct�Q{�=9�Կ��bC)�`�T<:����[P�3ȇ�C?���]J��*��O_��:ñ�, Mh��#�?1i$C��/�H`X�0�x����P�ts�i!mZK�=i1�l���>e�$�8�A��`�U��t�߁�K�P�g�����Z��;����Ⱦ�O��3���x�74��6�!}5~��:����3�	q�����e����,��h\��k?�au�}����4�Oft^N�0����o�|XK�K�����rӐ�rap��a|iD�T�C�+/� (Ϟ��5/>2��v�L�
m~��h�
`�*��1V �0__�vo��Ϗ�	�'h���|õ� Uyی	����q�i�9�<�8Ƈ�����+c��Au�=�vp-��k6�4dЌ���IH�4>yS�Bѐ��c���2�@�[�Y��}B�C�r�i ��,��� ����[��%�Wq��uT���F*P��
��!��_��P2�K�n�Y�b����l?b�@��� �RQ�H��wa���?��[�����e��bЍ�c��4�6��Bd��	5@�k���X6݄W��>�!h�.�UEc���Ӫc!0S	����'��Z�y�ٯl�E�-�ER2O5�t�? o��!�@���G�s�x��.]����~�iR611_�!y�N�k��?3&�LӒ���� n����NM��dr�n�BG��Vq�Sw���;��1u<4�l�o}{an/Dj�oVe�.N�F��l��S!>�n"�n��L0��c�D�x���n����W�B�LB��T2������)��W��aP����PC�Nnv,J`��Eq����g�'�,u�����Pq0��֌���#��Ɛ��c脨�H�n�l�z�o�7埄S��:o^�F�F~��(O��/�5m�v�d��?��zv�)�DKS�R�3�H5Q��*���u��䐿o�m.��?ᔕ{�5vxVp5B=�T<�Qɏq��V�,,��r����D�/���S[x)�����ђ0;��U؊�vr RIudxu�%{�T��^�4�rQ�Y�S�U5p�A�S0����pWj�Wkx:�8���	���u�+_��������70c�q�àf�U��#C�ֵ��5;�ي�J�̏2�}�N���BzS�I�'u���h�$��SH���=���8ޢB���.Z�8-��ΰ�m�� ��M3e�J�H;�u�ب��{!��O��Q���o��4tZ����2
��X�H�7���%���0�ˏk6��)jH��!�������{�>W��Ň���w^(����>kpOi�:c��=��)�,��<ԁ�-ղٮM乑�'�n�9�p�ɠ;<�í��D�T4��=(?9T��ua���2�C�s��LZX�+q��Ь|�o��;~�Q�2w��� X]p��F�u<
�f�I}�'�D��}�	�t�� ����O��R$2
�ݟ�����Ji4��[�]���GWK���@�
�0x���oN6�]�V�#Ҵ��)L_��'���f�mZ=�K�r� ��q��$�~-����<ɉ������y�E;1�*ݹu��V�:~q���Ҧ��#��ye#5��ۻQi��3���T��� ��.�6j���%���Y?�>�j*&cA���f|�(�(����H8�X��x� ]���x����ݖ0L�$��%����;t{�#��ɏ?�q�*�q	J�_��ʂ�;2�"6.�=ė��ы����׋���{\Q앺$��B�/������ݼ
������o����}=��K@2˓wd��ƀ��I�C͸��3��Mi��﵊%�=;"�d���R��;:
�.�^������T&k�ݿ�_NH��3�e'3�u�Z*�h�yZR��ns�