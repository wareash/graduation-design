��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@���$U[H_#�/8�y��,��F��`G�m6f�f�aiI`������tC����dl���=eZ��^�٭����B�FYĸX�G�����݁�]}~�s�cC�_ �c��2)����$�a<��d�6�q��tӏ�ˡ\s�$�L���Ÿ|^*��g�@U�*2�X���2��^�:9��D<��;�h��É}����a$;��몬g��>��W��iv���o�ăN�G\\�[�4�������W4xl��0�;O���V^��@��l5f+��\�&�7F�CqϮ�Y"�� C�T���/��Ƹg"���l ����~G�_y�kIe�+E�9�>Ǹ=�oWS�|���WV��P����������L��΋I2�G�r	y�i&�l��vЦ5�o�#����T�WrkV#��+�ڛ����C��ɀeG31>�����k�\�%�̶�@J�%A-�@�'2�}�0�΋ha���RN;zy�Q}N��5Z��}L���Z��¼�1<}M�����g�) $�8��Ρ�g���}E����G�@).�b���L��<�1�~:�~"�S��Y�p*-��^(Yj�����k��=98VK�ϲ�=�Zhy��� �#��_���c���~���YƯXrh"� Sao�%��Ƭ�;���cE��:�<:���6��E����Mr`2C���L�g.�T�"/)(dAX �B\\�xG�� ����	��r=�ى��x�⿐�z{�&��!�$�ȠC���}���?pEp�����p���р�e��Tu�M�@(���v6�ɥ.D�{(��Ķ)B0�h.ˢ�ا--��I�OtQ��I�ǧ�b:�ot����'�� �AvY��ɲ��c�Q��h�v�z�Fo�6$�ǧA��h�;�X��?F�4�E���j���X�Qd�i�� �C���¤T&=Ò�z#������z?��:�]q�����'Ca[q���?]6;��TO�c�����"{�K��ك���u�Rଽ��^S���8+���8%�����9o�[��Z,I�i���Ⱦ��aPw���ׂ�pV�D'ƽ�s���0�m�%5�����:�p���YUP]�+�qhw�[���(��5�1,j����>���f���eׇ>z[aࣻ�l�lU�E��|�R���o(m�]b��A��������_�p��bhy� |K�,�QT�¹�]P~�d��~��(�h�|Q����v����V�h�=�z7y�+�Yq�۠��7�YӲv�e �҂�d��e��b)M5� O�@j$7=l_����8�������t�d��	��s�u�뼽��'�|*�TpX���ѫ׆C��.^�a-��V|#��u�I�ˠnY��=8:9˺�R4)ϱ�M�_%����N�NI�[Q2�c.&���6G��ҏ�������uc��I}����� E-���z^=]��W!��)�ڬ��;�M;gֻY.��ھ �H�L�?�26S�#��ԟ�7ލ^s9�D����i��J���ވ�Cs#�O���i��	h�-5𬓳�����uK\�ƀ{��z��]�1~��/���lѤ${\:��=��+�z�ce� ~��sbӀ�~dS����+�D
i"/��ʅ��L#��N�!�1	�-��j
�98��㨑����K_�LL\�h�ĸPSK
nTÈsPf�o'�.����;Z�dS��y�/0>�mT0�^�\q�J�=Fh:�7�?'�V�"Ԛ��ܸS&[2�W.*mE�����컉�.����F_���7@,�nA�QQ�	���Lp�W�W0 �
���}��q�1:k]�L�i��`�]O�T�߳�%-6>��k��u���U��B�ʰ��{"C��^��ޞpp��`��	��Q5�����"��}��hW����5�'�W�)Oap,(�$�y)�]w�!�5�Dv��_ϫ�2IuE�N+s,ן70�?�F�D�h?���q���&r8�
ډ�Rt��s��GK�����&e+�/��$�ny�oˤ��(b�:�V$�C��؀i���5����!7�.���2�(�L���HSh�ŧ�����eC}��f��n�\��E��##ޏ�������AMn�f�y}�_̰\m�K~��;2��$T��4��h`������֍�ZF�񌼧�p��Y����J����&�s�gڪ-Č���-�fG&&���:{22�V%8c��nP���[�!(X$�X��R>Áw�(؝�ow=>�9�T䆾���?�җ������Ia�UU/P�NSmh+��n�P k���ڞ3��Ҟ��ki-'�k�y�-��%�ƈ�H�����I�0f8}q�2T����o��)��v����|�E� ��!�Z�Q� i�\'�>��Y��8+��)��2��m��SII�����������R����/x>�GZ�[U����}A�~wt�L?�/�l���<��!Dl��c��1�O�:��)x���r�tf��	�Z3�"QS����hoY��*�҆&�)�b��������R�{�= ���o�HZ�c�7
%�t��BBB
 y�}cL���W���a�?��P	�ІW3#�{�h�����],�f"���V}�S�A�>�����x�:�7z �w���Z��v���h�I�j��������uB��i�n7�����1�E�ao��ˍq����3R�A�`Rg�h�ηw���Wn�Ax���	9�:����e*ӢP�=?�x�$L�ϧ��j��J����IƷV��<��k� ���=��MƓ��s��m��}�{��#���[���I#�y����۫2��ё'�����������m�q���s������) �#����	$Qs�V�o��*�&-���o-������^�xf��c����
h�GB���k����n �D�L�����@����$q��Cv�?]���JM��"�8`4��]ΰ�-V��.$� o��T�m�ꟙmBw *�u	o��B�(J�1��3Q%X�d$3�Fz3;����s�[�h�A^q�N�2lk��C����Ϗ����(?�h�#� ]hM������f�Y�H��%�09�0�y��%������	a�����(-n��:����/S<.�Clz�E���˅���/:���C�r���G�i�x�<v��Y,<l�[����v.ُr�-����j޴��ѵӔUݜ��/���RO��n��@������1Ƽ6���x=x
@6��c����;�j�r�Q��UFt��9�X��&#'�a�*j���̦T��#��z+�*&�8ʸ䡶Ep��x�D:C�7�8nᘾ��xٮ�2н�d4�5h.���s�#'|�^������ia�|�Cഅ�%sHR�W�⣕��s��ڒ�P�l�iQ��(y�u����-��^څZ*n�z��"�� �g������R��hK�qiį�TP�Ieְd�\�]sl�owI����8�ia�e��G�AS����>�3�$�M�=�:�6+�Q�R�&����յk�J����P��5�֍r��C���.��oh���m${�K�/n���ZAL�kU��4�M����v�����w^k��m��zw�P�>�:����=>�o,�ꪩ�~.jKw�����|A��v��� �j�2}e���fՋ^�_�f��C��h�k�2�~C²��.��&,[x2e-%�Q�[��5�v�gB�r��3{hV�t�H�rP�����*߱
���P�[J���j��s˔B�Ug�GaI!��8��Y��vnu����'��b�eC���Ű_�-�q�:@��$ m�K��j��C��&*�̾y<Een��h+�eY�Px|vz1cCKj ?����!�g�_U$!�D��
���7�̀�K�h�#��^b���'-�V��-Vf1'��d�A�aR���I599������1a�����e6����f���TE�	�A�&�W�NB@�����2��I�Ĉ�� _�9�!��ޕ�$	���8��a�X�݉����-/m���w�&|q���LbB��e�uӟ����d����u�2Κ7V��l��h.&�/=�]^�����e�<�����j��]�G�]3)���~���ܾ&�)��`��?!H�� ��ŁϢ��O�`j?'<��v��}�\<�NI�@*�0tDP����)O���g����"%���k�H�ŕ�2)f���@� ���og%���=fM_��&I얆�	����9����ᧉ?��n�U�H��?A��l�U�z��|_B��������]Rя��G#?M��T���s�=��R�2��X,�]"e��i�����1��5X�	�K��3�B�G�$ϋ���y�n�����F�.��۝���_Eb�A ���r$̈��98aH㤋9	p~��Ⱥ��$�Mq��V����n��D@S��P�^�B8ܻ��`���#qn@��VS��J]-k�q9�̅� 3R9`*�1���D���&�W�����^�Ы�����F���Qa5��z�N>�H*ԧ%��"�}�|^(�<$�����@W��7w���%c�˫݆
��؍�JKsT��Y����(�V|*	�V�s~qd�Z��͏��Ţ���i�p��tGyC��{ǔk��D�r_��ݒ�T�<�L�v�-��\k����=�H�&�y��#d�:��ZﳽY,n/u	�
ի�r�
�Qx�q��N���@����8�/��TH$ֻ�� D5B�m-ϵ��$L�����Y��m{��^�A�PE��Y�T�����Ϲ�j�^G��Q+Y@4&UkEAz��_m8��F�T�=f�H�-��%�v裼����&�x��Q�qԭ�]\�<�OM�2h�E�������]�1�vzD�l�����X�	��0y9xe!q�.u�b �Zc��5���J��7��6�&4u���Wo��
����bh�S�틄�>�w�0���":	�c� 
k:�|�V�qEZ׮;��.�u=�2�b9La�x�iJxB��X���q�i��	�<�ƃ����mw �o��NN�gD˱&%ti�a���C٪��r���hȓ��+)�	�V���+e)��a���{�Ӕx�$?���o�b�P��|]e-�Ð�a~��*j����|7��#��7�Ij@Tr'ub�T��lXvZ_��!C��J�u(����D��ZF ����vH�V������OJ��=���D�ߒ�*���+��-a4p���/t%����~!�>R|jef��� �ҢV�h=	g@LI��G�ˎoAL��@fS�X���Q����h��Z9�I!�hޮf��g�A�4��4�d�\����D|n+��!�Jb�Ր�s��$E�����	�Q�kl8��hKʡa5��[��Q� ߧ��fۗ'e^bѮ���u�s�|'+.a��� K��+��ׁ���p����+Jh�0���R#��b��2�53��_�r!�x��D/�}��ɺ�¸"�&&G�;�p�OSX����j�J�n��s�y>#�'�n{S���׫��:ԧ5�2���OD_�ksZW4R����`���迓�h�t3�I.!O�Q	�֖[.Tg�����8oX�6��w�t�`��H5D>#H�-B��G䀨�3ɾ�� �>̙�;#��y��[FV���۶&d@��t�0��ɖ�4=c���~A�z0�2��H1�P���9�
��ed�ew���\�j�SkTnK�����1M�F��S���5\~|.J���Oh���2�}