��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf\�|Vv �|�
�����W+i\�d����;o�o�[��e@[ġ�%�#`�G6D��v.s2s�
���Ϗ����1����ŰOy���f�˜��G\�'N��)�b��؇�>�j:�~��@W�/����*����)��T�vw�,��)¶��s�;)2�"��v����v/���1�qX�T���.��!��Y+��.:1&~x�:Dy����mƹ��Mz��1�V���B��n���t�l��q�����\2���=._c"Dك�X��?��N�7X!wI�e��^�-02�<T�۟ۨF�Uucn�{�KNe�x5�!���\UŢ%�hk�G�|�D`�� �%O(���]����Sq�h���1�	YR�Pt�ґ�?~)���'!QkW¾�z(�4xY���t�.T����r�G�G�qC�3���<�;_���Ah�3|���@�lG�ʎhf�J��g�3R�(���Nu� ����8�ږ�*z��+����pjw�׺��f�(@��Y	��=��I	V(�Óh�2�JKeB���.�&%
�Ѱ窮ɗ�vg��x�����֛�հ�`��h��&L���^�b�A-�����xh#�3R_����F��G�ݭ�fS�	�(j�`����?�M�2�;�<'~��Sn��*L�,@g��o��T���^^IE�v0�T��!4.�פ��盞�`��X: T�> e���4�vꩌ1
�����,چ���siO��M�΀"�q(������\}O �( �22����r�#��M�Bf"
W�"6Z�Z�wC���-u�+������;#����?H���~҄uW����Ɨ�a�[+v@��E�?�>b�xA��������\�=x�����NF<Eb�ڕ��c)n�v�5�����a��%���P�x&�M�P��(�r��Q����u5���_���+��@���r���ꗤ���¾>0�!i
lZ���{KQpP���nXF�rx=�=��m���K>����r-���-�h��˴�N���$��/�1��iEe���2��I#�SM��3����W���0k�� Ҙ_���������aØ؆	ct\�z�'@��Pc�'�ӧ�T�1���z����t�C���cbyM.'��o�����W�o�N�OA,V�[��v4���������.����F9Ce6��d�_�Y���w���\!�O4?��h-4s¡��?W�PY�c����e��#�0���5U��y`�K��D�r� ,���I�	����bs�����6�\�+����X���Sĸ�,�^s"�Y=�AT1G'��L�Xح���r��P�UL1Q�)�f����th�`%�E5t��(��+�j$�ǌ�)f�����A�w+��Ĭ��C�8�$����%t�j�7�kjRx���Ig<Ԙ�s}x����A�'廙���QQm�e;�q;r�Oך��ϯi��z��i}��`��Y|��y���b ����Jq�=�����o�~�ss�:�q@�n�"4�E�%N�[����{ZK�`n�/1�)BC�۽���s�2��"��=�A�5��e��<i(�V)��l����䗎�J�>���#�-Us�5�_��6����Fz2����o5�i\*�3� ,�A������LK減�
�3�p.�1�/�VI�)��YQK�h[����������Q�"�����J���ieQ0oU���>��ׇ�YsG۾��v$���Ҹ�ոw�+=HP��Rm���n�d��:����TD��B�p������rY�V��Ku���F(D�!��v�U��w���[6_�����qp�Ui9-uc���d^���
AӍ5�c�Cr9�/~b�f*��E�m��#(8�k��`��t��sQ3�ž��,oi����?�Fݟ��A��t-C�)2,��-t�U:f7���Ä��)�~N������o�%	�"�|�Rh>�<���RvZs�X�SI=�1�p!+/8���.)�3�uw-�JPIU[�W����^�p�}���㱊}���a9�6vIP�?f���ܾ3�[f{P_Eo�2B��_�m�冔�Щ��-�]ᤨ��6F�6�NX<_ŕ{4�+�5$����[��4��ʹ�#0�j�r|Z�D#5�0�ow�| �;�E�7�>D�O����#�����-��dJ&��zYMf�	숺��6�{	0�d6$�&~���OfWװzڝ�1bL˝���T����U�V�*v05ri�v\p��D���u?���tF�)��n���[1wW����${0�ﴏ�]a�9ޢ��p��.�i�c��`og� ��٥�\��j��$��In��V��}���4�� Ω�ڑ�Ѫ�N�W�|5P]�6mc� ]"E[x�چS��O�N®���i�."�m��Z���KdD1w�2��I1�o�G��n�� B�VC�v
�g�K��a�Δ,���
%!g�+���ЈY���>>O�\.F�d0�3^�b�j�E�:fFJ���݉�ȹA���"�y�����{!�����;�
�^;3�]jCRZ��<�M�ǐ�7ȶp�i�8_qxm�o<�悒�sr+#vJ�u���_^ych�i�,/�؅���4N��h%	e�3V�/VU��^�w�j\�Q���p�4;�G��$Bx����H|���u��Kg������I+X��Ԅ�+�ͳN�����
F	C���|�V�k�^�{���n�d��etGy��������##si���upi���Jr�A��Ha�"�$���Z�0tw���kt8'ðh��� ����__5zɐ3μ��5�y��36�_����a'Ɠc7n���2�U�P$��e���`�G�9iE�pB��s��J	q̉�fޛ������!т{J�th3W�h�4��'��l�-�L�XhYP���j�t��o�nycs�IUЁ"�:�#�4R�q
{z����@	$�n��~����Y\Տ�Uí'����n�����!�"��΃'SG1��$~w}��Q�;��˲�����/&9IH�j�!蓔K�2�[��Y��>n1��|ߟ5J�xj} ;G{���`bP�^�F�00�W#����5H��V�'�֕�;L��UP|��W��8fK��ض��x��-#�-��*���1����\i?��M@����?��.��!�Oɝ>Ȇ�D�zhm�3����"!lu.�?�k٪ݳԿ�ש'�<� ��c|�	ԡّ��Z���1�&�Ы�fOV{�;�b�W�������)�4K_@��6-i�9�Kã��9N��1��C�t5k�/ae#&X�j�c�ڿ��ߊ�K1m��y�w&ˎ����/��tf��2�'���Cl�]�nN�_L�I���,Jpn�]_����?�=>F{~Oua�̫X�S		��S�����U�8��D��1�W�"B�����:"2��s���� ((��ۥ��ʑ��m�'�]<�iE!>�R��K��)��a��8��-Ҫ/ ��,F�Ȥ)Mg�I8�
�"^Kwg�o�Q��,���uSq�ι�Ϯ�Fi"��C��q�����kbG�@Y��g����"��	�1�R���}#+���J?�u~�+��}?�zs,
�5�4�O��az�>ᡨ�x���A.j���M�2 �����=rT��U��p�	�tYa؏)s�A`�%`���^~K�|bYr�R��� M�N��λ�O�~"̼�8��Twq^?b�.��ޑ;g}������oow������NЭ��d��ba(U�j�������y�4���ǲ�jTe�0���Q���-�vV�rF-a�w4���2_ "逅�]�� ��[�6��^�.͟��`�A+�o�:Y�*��4nP6!T)똘.BO��.C�q=�p�ݒP�j��ri���l�}�-�v`��S���W�]�v	�IV�f<�r���6�V���]��y�c�i"�ݖ�h��3},��-�5���M��e�+��)e���]鳝:l�$�ɦ���Ug�b�3P+�	\#iǢ�����V\�x��*��'PºEwWe���$fY��e�Ϧ��Vo��+#�g�,�p	?��E�j��+��t�ӝ'���Td�r�L�"�����˪��_�"�?�����(��U
-c�x��rPM:΃��9�U*#~�;��`qo��2ͦ���E�NA��DM�[����|M��Y}���Zk�A6��Pg�a�i�2k�L�>ʂ�i�QE���%��b� )�;����y1�(��>�'�w�T�eL��%��[�.r��A���4Y,�Ҍ�0O��-	�Ri��*NLK֘��U��@Jz�P���Ƣ<�+?�:(ؽO�
���)�>����K�ps-9"����I|� �{���,9A9������s{�����n�b�ڝO�g�xP�4�-ˋC ����94|�
ƥ9 ����9!f�_���1�J��5�{h@�9Jf�l���
�tgg �8�֑B�ڂ4 ~��]R�#d�����4�,��C���:q�z���Z^l[�3*p�·P�|�����|r�$kàGQ)�d�Ԗ��Y�T7��g�����LK�ƇP�̗��XO3�zn�)Ħ���r�91�S�`WC1��Zp�8G���_�f�G2�"O��ڞB�e���5܇�۪�3[3ZZQ��u���"ނ��<�٦��xIbÜF�@}����T\�,;�\��DX�_�����X\Tק�2��2Az�f�:��|ڒ�/���g�@ �w-oq�0��b7�,�U�����z���0��Z8���,J�kb9�=��PQ�����oW=,Z!QG����Ð���W� 9㬬��cR�7:�yʠ�U8��~���I,�(�pl�-|��� (��e5���N`ޔ�����g��%��_��
Fz9��͂�*Ā��9��S����p�͠)�l��9:\o<�\ٜT�h���\�K��is��_tI*��H��Iz*�6`�i��l�=5��YX��ڔ�;�9a��p�O����-�!^IY�7���q�'��W�;�	�;J�ʩJ"��O��E\��t�Tz^��>��F|g�{`1����Ce�T������~�������������U��yT�A՘ʉ"עnw�[5HY���t���1�������Z����􈉐�f��V{̍�9eO����N�����/3J�JuQ�|dK����굃Z"1D,a��wϜ�p)�c� aH;���a#��&�]�=ų��#j� 	�${�tP'�Hm{�N����3p���9�/�Q��*2���av��%�A�'�j�P�[b����{y���\w���r@����1C����Q�Q�3Uv�TKBC�.�Т4	�&�*FV�G:2��D�cpa�f�	:��&�`��6����+n(�O�Q7,�5u���0qQF��4���sٱ9��������+!]��m�M�	.�J��q��q:@�p�ފI��G�B�9GЫx�!������7�Y���c�eQL�(�d���0o?X���9�N���+��`�N�F����E�!���k���}m'D�E�n6BA*ҧ���uSc0*2d�+G�Uo��Q��z6����/���S_nHN��7Q~{�-��4�_3�/.̓�/����U�T�}�{ r�Q��{E��/ c�]����sW���	���Fi����wL���|of��ۘ�Rwsc��?�.�܌��
�D�)
��r�v���^�����'h�����{p��Qqm�i1;��r��i�ۭ=N}Zź�;��?C1�����dc��[|�.?((���4&�ku pg���Y_lDq�|I")0�HSz(��Dv�K��5���%��"�&�S�k�5�%!�s��Y)�U��]�X�j�Fq\���1$�2�֋�Eg�|]�R����8 �e���qR)�iBNc 慏�E�>Z�'ٶ���%�\hｽ ���-����P��c�<�ZfNHa`x�c�`���C�A_rJ�<��s��z��� �jj���y[ھ����������{ΡY�售#60_9]�����N-�8E>��_��%��AK�S��^YI\x���f��êB����L�9�Qtؑ�ٗ�
�P����x곶��^��dn`H�����Ѝ�A��ʹ�躖Mߧ�+Ɖ�t@��K�#FY"xop[O�}7�����?T/���6�8�-��	����]�ƣ�*`^:�9�$���!�_{���ՆI��Ҭ�N�PH�I��T�d�q@�&���kv��s!�egZ�F�C����%p�S���mD=����t��	Bl��"=f�J!*�^^���}�cg�V��[��v�?Fn�8�g�D�7�0u�qek8� ���N��(C���4�1����"^0s B��1-���i8{����oP�(����*��Lk^�: �akB{X)r���h��'*��m���/�`��$ս7�"�^ ����ce������=��9v�g��5����M=;C.gI�aY����_�\B� �K��T]6ς��S@	!� �%Y��N�Lډ����P���[�vI;L9+��GR'9?�*VI&�	38v��͓�p�>�՜�o�x�;a��I�s2��Ȓ�ʞ��{��1�}N����t��d�ε���Ȕt�FG��o�����7[kh®c-�ίHy������Q��G ��L3I�(!:�j��x9v�.��ٓP2 p�õ��Z ��;��A+!�lU��т���0�m8/r�
���%h=hԎ�W,���z�����
tI�#���2c�_%z�vO��)Z1��T5����2��'�

V�̲�j��ծҝk��B�7G1#+�B��@�����;Ha8���A���=-$_K��)EE�@�����֎���ۛv�n���Ԧ���f�N@S������E��1Ä�/WmvʂI�(�8D����}�n��XF��8��P1�&���uj�z��d�S�@�]�x��ۭ���C5]h��	�����~�k�ڒ�#�3J����o�DH�8�O�G��u_�:�42#��j��g�,k���R�w%��Q����M˫�FE4P�܉������4C�:P�[DyiA� �M�O{�A{1��x�%�#��{e����2��o!�ws܏���p��h�@��/Fh97��%*[k����PF3	��Z  	�y!Ô(^Bo�<']A^O��:A���8SlϏ���'�g7:KI(�
�r���cgQ+��9�D7�[v*l�)��(��-8s>��u�����|�k����d̈���-�)<tg*�x����#��D�R�+��@�ޮ�ʆ�{�K�
`�R�	�c��$�[dO�m�[��\�V�?g7��5� �L�ڂ�J�2�+��
�T�X�I�h��6�����K�+@끶\5�&���Ԋ�*&l��;=����:N�n�S(L��J29���@G����,��E�ET��>�K�w�VE��"Rt�����	hިA!ln��T^p�=��,���)Ļ��ȧ�}k�u<�|:q~��D^�ų����e$O�2��F��1�i z�.UOĈ\Ĳ�cS	 ��i�N�i}���
�ֳ#� ��l~4��X2�%ۉ�'5�q�FC<rl/��ë�6ޔ��?Kh���a���5�/^j��U
�ma�.O��Qd!v�Rh p���>Z��_E�����n����k. 3OT
��S���?r�~��}�k�_��8�ג~޻�b��_�W:�K)*x�	}��jL�η����7Q�,�3�J���I2�X�<����~�U����b�sd��>;W~{�v�DҦmõ��'�@k	Q��t����F��O:�u�Lc'�濯6�X`Z7�g$��NR����������o�������,����þ-hE%^�c��c�􅟼O���*��=�؎�(�ToH�]'�/��t�G�	D�`���q����,Im_	#�VGΝ�}S�J��ܱ�Sim�|xa+�9~@�6FR����T�f1��M;�و]`P�)��mo
я.��÷`6 ��g>A�_��N�(t싕�s|{*߄ݹr�L���`��϶L�]�yuR�݃�+X����%`ݎs�>NM9a�`�l:��#�k1?:j*p8��}�'&JŖW)����+���3���_5*ծiI�6��f�AG�!%���/+I�?�*����pe?�;�Y	��T�0[���
j:=[+7��t�'�JK����S��GVlÞ�m!Sz�B��mm���d�y��3Ⰶ��]�n�����X�U���4�q���,��u/P��}V�2[h?9��|$V[�*U:��kebꯊ��a��B�w'�bNVv��.���Hq� ��گl�!$dB#�On�-����y�X�'(�S�y�\9��c����,���C��Zk'�Z�|C��8�	�ܗ�^ӻ��m��fPh�G��=�ڭ={^f�S��ޚ�>QC�R	��x}�peA�	���<��'�|0U,;`
���>rW`-}hUɈڻ8�0?��m/�v�e*����̙�L@��/0L��B�A�������H�P<SpL� ;��h1��D��*bqwX�����bo ��+��� f:L`���=iG�_Q;�e��㱪WsM��|
u��8��u�����]���ړ6=C7�
$�Sd��6�1@�Á���e_��8��bg7�ķ�3z|f��t�z!�qNl��<'b��3s��`_ɪ�v*!B����S�<A��*���rj�;	y��ɺ���������VY�a$ʨ��r�?�*d��J	�)��S32�VL>�(=��z�'�R��!����lI4L4���z��{�D[�\��g�ɝW�d��(���K<��a��9��V��6��f.���\��w-��!"G����~5���C��*����[�L=���-���Y�t- a��r�J$�.�t �Ý���
�{ʞ;x�9eP�`���C��lm�f#^��UA�ع[�b��&��J��c.	�j�<�&��]�Ev!=t���^4�c��Ȼ�b�r_�p=`j����1�$?eɂ֢+��'��߰þ�1Ѵ��To�'L�;�����j��3�>7Z�Hg@Mvp<���@������ŌC��,NXg��J7z0m&��ʙ��� �ײ��F}u��)�f�ez����tŚt9�B�a�R����&YVz�۱�����ן��?�8���:�]m�N�� 
U��s	o�:;<�,�L���t�.1��؊6��,5�]��K���i�λ�N�Ѻw�1$?��H��1�j�l^۷�9���7����%�sO4���P�yy�tOlb��.��x�+~Bj�D�<l�Z%��8��R�/L������4�5�𛀘�l��4�y�ķ]�#n ��y�a��F��h!�wh2���x��j>C��>j��+���Yf�V ��$��E���/�kn�L���������
� Wa��7����(��ϑq�v&M��Ѱ�j�Z���R��	��؂ھh�HSj#���26!OW��LhAb&������+�� ���E㉸.:|]��A�~o6�he+fu�i5ᫎ���6�4��P�_^r�W��3w̶=tsZ�Y:��y����~������F[QS��EWܜ�8��l�ڐQ�\�XYEcbug�ى�[)���$Vx����I�s�ꯆ�؇���Aj����o��R���ol�+qy����F𷴊Y���8������7a����f����#�&��'����PQ�]oR����O�m9��*Љ�}R�g�E����vQ�6��C��l䭃S���B|�a��oY�J�M�{�<���3�>�H&P
�S�a��7J�J�k�f7��o�8�
n�0bͽO�)Bp��'F�|��55޺sg����[�ְ�
$���3�s��������A�A�j5�8�Ê����۷9�l�U�K�P��e'h�tc�1!�f�.�7s����İ�mr���&x�hQFݢ%Z��=x��s���4���옅��؞zfY6�5�d����{���|b�jh���$�I�J�`щ5����0pB�$y,ZɂV�T��ؓ���4�ɶ�e�$
���������Ps������>׎�6ܑ���")R$�r��5±h�2��\�O�ڶ��F�d�e�	��o=Ū�����xZ�A��i��J���z/zr#6�㕙�Jx��7n��/G~ꓘdʴ���+R1!�}ds�f����� u�aܯG����U�ݠ���@ƕ�K\��ކD��@r�^����4��^���:�E�El�q��E�P����1o5̺v�����v7�S���l�	�\B��a��z@�OR��M�����WȔ9��i���@Ӗ��G��fv�0`���X���S�c�o��!�)f��x�'PGx��������ћ˅��Z�<����AF�{̑�����4����.��z�l*}���:�$�-	�T4<�=)s��V%_S�<Ⱥ��uz�Ѻ�p
��ڒ'�m�޳����ϽM�S=´)#���NG���c9�����q�'�����&jDʳ���	�%��M)�t+2_ԟ������P&�4�����v�q���EE�sd��G�Z�m�7�@��m29a��Mc�78=A3�y��C��ղ%�7k3��C�ԄB �#x���>f3��h�)e.�ݓ�M_��Wt��S�W�Og�?��>�����O�ƌ���8��t`<L�+
b�^���"y4�R�!���Wn�F�@Y��@�M%��ym$�=�(�?�4�@E��x���O�΢	��T�Y*����7Xrj���4��*C��oe��	���5w,u�u��F���N�Г�"b���<%33�$���<��O�g��J�68��2(�Ԏ�J+��L����������FĮ/�d�*s���N�ݬ�y&h\�`�xO+r�B�A��gŨEbRj"��|4��e����#�����;�Jh���:�����W)���eѺ�=�⤜�n�Lo�JJ+�L��\�z��-��_<�߭�ü������ݾ������8���0��E��>+d������K�ܭ#����Y��so"�[)��`�EKB�[�x�t[Y��_�>�b�]S"�-p�PTD�HS���������}���~�����WFe{�����Y��;�9q ���x>�� C�:�]~⏫o�W���A�Gj�K�C���$w9�M��
���K��E|%,��U�\ŧ�!��l���=`�R;�<�I�1:K`k
�g�bxP!~���B����qs��}d������*42q�!v�Ȃ��>O4�Eި��8���T�x����� ��1���6��AŌ38�M����tq(
��R7�2��+��<�}�����6<���s�<�n���䕘�bte�&�P�������<��5�e��'��>�����lþ�c�\�:a�<F /@��3�_���Bf
$��`� �b*7��3�˽5�u����`��JuO�e
���͐�����v�'�0*~{t:9����y�r���0X���W��P̬���;��PC"��@�E�ޮi��O�����.걙�����K��G��~b�1C�R��_h�M�!L��=�c&����䈺8yf��v�]Η�AE_��!��i�J�2nm~D�²}[���'U��� �MI���4�}�'݅�۲w��K�l�'JszQU������������O�J�K�pIɗ�\�J�����!O�P��a�R�c"�?R��q����)B�m���������ZA�!+E�8�O���,"4$/R�*< |�//*�ӝ��!���J�@�l�4pކ�5l��iR;���	�y+��8��86xCH!V���ʋ�+�Aw�����-�߀����e-����ߢ��_7��mW�I&�0�V9�t�`4��1�.�B���q�T�?�|�3�3L����@�����tr�+�xK:}<�߻����1q%�	t��U���ͯ�OY���%�1_�[�КL��4���� ʸ1d{������.�}D����=�iJ�p �j?`LN�Y�~����������w%`D�;d��j��e$��Ab[ܛ}zA\�O��ў#� ˂/�C�{�Ȕ�W�&�n��:r�i��������rx�Xȇ&GC��Y�*�&x�殯Üҟ�˿n���05�����T(ܮl��H�^Lq��������A��φ���j8-��245�@��큩�!F�Q֌b�uFO&�tb'��H�O5�7X�ٗ�7b	I�~d�_rX��X�i�|�7Ќ�R�r�:8$��j��8�q��ɯ� g��}��|�C�Tu�pZx��䠯�LoI폕��=#Y��g^��(�e;K��UWꬑ����0"��K��y�&��
�����T*���������%/�4�8��Ѧ�La�R.�����
�r�mϊ^�S4QD�S��LħB+#7Ɠ�1�E�����;,s<a /�G��I&�f�fj��F6٦>ϳϒ��~Eiv	�ĸwg��*PZ�7K�Iª�=m%u�z��o�� "�<_�u�(�PW:Xz�i�܄eYu�ǉ ���F���@��@���᩺	��i�D#��'�c��{IӘvK�^S@;����t���P�|ά}R�EJb�%����?�#b!dCbC$�6�M`�%l���F%��l9�QD��۫�ç>���zY��U���%�5�i=��L,��0���/f�00�S��D��ٲ��9�,��tDh����<����h�}����f3�e]qi����4�r���{���#�ϱ��۰�i��og���єw�����, Y��1't�*��!�0�扸��ޝ%*�F��t,\5�`�ݴ4���v�F��
lc˪:h�A� ϭ؉<NRya�0�}�Ws��O���(ltT�A��Z�CA�������TM�R�^���N0|/�,�������f���r$F��N��P����s��L���/�N���,��r�`1���*6�nk��%����y�d�J�a6���=V��j�Ėم�{���@�������a`�dӴ�����I��g��T�/�>#!�^��B�K�2�9v�:jcw�yj�B��!��K�c����^��ejAV�56�����fI؉OZbtKt;t���@���sKM�p.^��W;��ky���N��l%�%f������$�%�쿙OV< g���郪�����{����6������ �������l*,U�M?�#n��=�Ds!�����s���r���\�����N����7_�Q$q_m|г-6y�ڶ�o ������3le�ѽ%_ʨ������ܣI��U�8��S�W�r��_)�%����S)O]�*���1y��I�qgF�Ԙ��Ŧ�:��/|�����YR�X�L�K��ak�������q�v.T���s��٬��H8G2��ч���] �(���;�e�He�	�Ħo��;ʌ�Ǯgl�C>L���������,M�5����+��7��ǋ��_�e._|zGϣa#򁐂csa΃΅�6�1jI�N���6�L��2����~�8�ic���RS�36IWR|!�	\������I}>�Һ����ǩ�M"��Ab���&��v
��HՈD��ӏ��ZN, Q>�ܳ�}�ӄ�tc-i�ǲ�ݽ�aS���1�'�P���\��\2�Oк�L"�NS��%o�[���_v�>�h}>���W�ĥ�=�Nq�Ň�/���&�Q`�I�v>��z�~���^t���yb����n)��93onn<��y	�)l���)=��]s�:�ԋekJa��ģ��JJl�`wD<�����YxW��d6	�c�����s1�Sc��N:��۔q���Ӌ�v�#x�)���ځ���?���S�z���cG;��&2[,l�WM�r�&D�|��P4�D��;��b�.��y��\0h������n��b�T+7�oY¢}G�/�� ����`b�����T��t�\��(ل��A��V�K��T�K%'�)�&:]���8��tpV�>�Z~�� "?W�a������|�)�l �d��[Z��x/OiD��Ȗ���ojU���05�N����&�v-TjB�,��^��/��у�~ �-/e�#/�dՉq�2\q_i~X4F�C*0�h3�H�w��$tu~V����ג��*�!f|�����Z8��I�����}	����%�վ���#o�3�3��T� 3KN�W�2��$2}�~Q��إF��]qܔ�L��
Z�c�%�J��\���vhJ�Йff�km*^�|J�>L?�4�T�$�T��r0�0�õ�h�(v2f[Fs�~���K:R��SR�.����X)G-Κ
��<%��ތ��BT�x�����\��MDcb���"�e6�w��E@���������m%������%�[�����e��+���L�BI�k�M)Muy�~,�Q���9\e�%������á�Y�����%����"_�����Gc���J���L�.�$m��7x$��yW�M�z�2�1���R�z,na��wj�B�1'aZ���/n(�D9�.I����vY�s�+�-���()q���"O��l�K
ͅbM�Qa�l;�\Q�����j�G�Il.KD����%�y�e_Z�W_8aE� ~@s}�sj��]��VT��hG5�r�Σࢤ�v�~b����6�6��ꍉ杸�ƖP��ё�9:�@�W�$k|07ԑ
�g��%�헫۫OEM.�D�69�c8��i�V#�3��?�aD4��Cp.t�XY�K�{���Զ!��͡�{NDx�M	m�=��N��ܫ�R����	L������>�Ӯ;� ��45E�5������cI�����p��
���4�ME�������9��KN���3T�y��=�-,,!!�g�Ga��z%{$��D�ٌS��!MNU�R����t�k���-QCJ�PQ��(L��&�̙����\��ļ���m�e?��}��`
)�Z��-��6��(M���*�o�`�����O������5QW�;��@�"���m$�}ی��ɷ��B -��$X���K9��J�.�~�
ra��XF3QƊS�(d��|:RV67� ��3�v������pB�TE��.�����[iy�z�ç3���#�P�~1띶�������S��{������2������jsq�����������9k��.�����d���lW|����J�-�X�>���ϳ��(��O�@T�w�%S��`Tw�y��7����.KHCs��N�R~���͒4��H�Uz��~����&~�鷒QFx�Re����A����\�Ҷ�E���^�KNYГ6<�C+7/'i=���xL�䝊��Rc��"�Rِ0䂿L�8�ù{�	��Y�U'#~��W��6WF�X7EP�y�8���I���yUB���뾷)��)Jȷ�߱h��ǐ���)�79����P�ęYU�ɟUp6h�U���u���$��ɬ �����X9��G��G��c�<v��1K�p�4��VY{�R~�k��[&P��.f-���npq}�H~aB;0O
�{̳Ϣ�pb�O�v8I���``��sU�(���A�z����d{?����_�j��+
f��q�%X��=�	q�w_�2���~x�莴��I�:�m�Ȣ�r�黤j�=x=���u q�q5b� ���������������qa�+@���,u�|@9�z��+ia�b�ߟw��X��P�sCY1�khK��"�5�}������Rb�Wg}��O�I�4?fOɘ�Os����Df�ο"t�U7����c�����Bc��=5��C8O&�`an�m��H���ūܦ����	H[���:����̶C>�3U1Y12�[w�b�3|1D�w#��	�m��?h�[>�
�f�����P������_f����C�2P^�����PA��~�ޯQ8��Mc���NY�pBf�>Q�0>ƴ��:,��g���D�儔M���9U1fV�B{d�W������,��>�
5���¨D�@�ڷc��ψ.�1`Y۫<��k��t]gY#\�OG#���
Q	�H`f̐��Y��q�٨z���Wm��/��mʹZ/2J�,�T���O��u�Wt���2hWd)��7ԍs�bըx�D�>��ŀ�X�I?{�w�D����W]�<NM��Vg�\v߇V�"~�����w���R��!r�3!�f/ʂ�LF�~�TH��������㛔��b�]������o���ȭ<��>F��/�]���H�X���[\N~�Ǆ7�ȱ�Z���F�J�~��6����@&r{�iZ���0Κq�iQ�j{$d�/�*�k���t왘wCT�#�u�;5v�|��ZԮdp����iD��<M��-N�iDfK��Y�c��å��e[��Ĵ!�ǚ��ķce�^r9�vH����T�F�t���ߡ�й�k��L�j�LE��:�J�Rt�8�_���޽+:�ZE����YL;���dJ�q��C����%���hL�w��~{���-#.z�=h����lU���Cg�%	)����.Z]�H٢�H}�" ��%�'���x����Uv��'^�X���Z7/d.�?��H".�P�"�a�m5GUO+'�[u_G/�dA ����)���y�\��v1������.��n��oͺ�	��z�\<RK�1�:QU2l}���Q���oE�o�߇��	oL�&�%*�g2��o6r�}���`;�y�'7�'?���5.[{��	�7�{�R mO�FT/Ǵ�ƅVTY;��+k?֑)#��!2n�7�&�T�i��㇎P���Re�&����N����I����ھԣO����OP��Y{{�Xp���a�����e�){����������ń�9�@]_��t����oG.��b$ss�Rܞ;]0dj>A�<����N��?I�"��s�UC��%{�n�{�wo����� �,�wq��D����&`҂��r�Y2�����w�DD�0̐��� ��d�e���U�.��A	6���������m�C��1Ϲ�=�"�1��͵A�����~���p��Ǌ�r�+���J��		Co�-�mvF�,�@z��6�/��
NnV���泊��?<���$��ܮj&��h�H�'8[O9�����O�ոb�Å�S!��:)dpI/�u�.�&�����7��(Ӹ�9p�6/�@���`�w�Q��g�ί�Ė���, 9۫���F�{Ch��R����ֱӮ߳H��Mv�F�P��O��|g�F'Z�5"�I�,��������>8+Pvv{�=K��|��6�@�t-�:�����,����t0}I@U��6���U�\�56�H�7��N�/	l��A	ض�����&U1�� Y�8�qF2��2vR�:`wѝ���H�v|~}�DhHM���2�� }8��ab~$��"�q��j��ow�}䩤��v�L*�lJ��P��3⛫�X�<d)f��%�eڢ���O�_�k��@/g��Y m�S�Y\C1
̫ ��㊂k�<E�O��n?�n�ߵȠ��� ����h{�v�t�3n��Mĝ=�R���7��-B�29N�v��>��#4���ӒR��Y���OM�ܬk�b�N�xǇ���[I�V'��ĒW��UY30,cJ��)�^�SH��1[J?��s]�@�AGJ��)O�Ѵ�z�f�vz�m&��,�Q�Ov��~�P̔bQ���h�X�_�H��Ig%n'�O-�
�'��?.��H����ǋX�- ��޺PC�
�-���<����?ܗv��U���/o6{�>�������N�0�u�Xx�ר�z�tG�U�k��h��W����ץx��sf�SQ��k;1��H2n�㨉`�'�;�H;�GmнS� CU�;L����:��`z�K���vH��x������G�~�jv�&q��DR�`��ӌR��p(�Бd�t	kmH�?�R1���c��Ϣ��4��ai)�?a@�v��/�����^M!�d�]��N��u�Ռ#rR��+��iK�x'!��C�+8�ڪi#�ĀPb�\z�#���,�K~_���`�;<>S^�
١�o���	�]9M�}�n�,\�1�\��˃���tt��*�������>��},u��G���3��Q��Ӵhـ��z:Qp�u�Wyk���d��;���T84\(�ҽ�~p��t�\�g#�㟜<��W{�B������4��HM���[;���� b��a��`�$/�k��Ä�\��kZ��V��a�[��뎞���^�;�/�Y!���0w|���{��Npl�GU��A[ �pײ%� i�J�(A[a�%�^6{�6� �v�gрfeApЯ&Z.�c�
�pp�Z%�8�c����8�S@���W�gzd;�3kH�C�
�Ӏ��_�R��jr^�;jG*�r����%X��n�e�%Q3nx^٢�=I:��i��b�<R����P��Ǘ^�� �WK�(�,[?�C(�'b���u(>��H��$����m��h���ʀL�Fm5�6��1�6� �������w�YsgjN)��h��tPp�7�=��O\k�q������r����l�8�vo�Vg��А
��e�Dc}��U7P�_5�$�vQ��@����eS��\^Sgn�m���Eg��k� �um�_��-/����5���t��s���s4*�����LJ{��Nd吪�������R�(�Ǟ�y�R�A�C{w�2B���:�ov"#�!4�3��ݶ�m� ���3. 	obZɽv��qk�f�f9�v.�
8��P�]�P�nG��D;�D���*�ۂ�]s��)E#��B��)æH�1��C��"��e,��)�7��^6
�E��셲�Xj?����<sƖ�g,�Y����3��� b�]��a��^$���Y�E#Β���˸���0����Y�T�`A�, 7Q�pl;<��dt]q�����5+}���
g=Xxր�Qy��Hn&���(lCd͒ ��CK��خ�Ա�jQ���v%��AQ�Hk�=��R	��*��������_���&��\��"�I��Y�Ʃg���Ϲ���-#�,]�_c2�\�f-�� ��Y�hQx*�&�������05�gO.2�KpuA/��]E�9��b�Ͼ��S׎�jj��%i4����a!�b^�N����1oX�M���x�ѐ�=��|�OAPa�[�&0$�I5]�K� \7�)�V�w)��O��ΰ9\��KQk��8��s<��S�弯Ń���M�;���T7��K��9�m�SS��u� �:͉IhQ�|�s.�d1:�׿�v����*���p�9����Qk'%غD��⾾e�5 �~<��Lp�.ؠѝs��<V��rs'
=��V!�L�<# ڥ�^�]L��BT�H�;4�N�,�q�m���@3Q.����&�?OK���xݘ-��UY���Q�����#����
��~�����NvA��0�9��킱n���a�&ߑ�������:Q�o��o��e���P+1���i/kO!��e�6Ќ�i�CAف ���3vl����T� L)��Ȑ/f��S��1o����K
?����]Ƞ�I_e������&�~T�ri���J�����kF���/iNX���<��qw#E'�K?2�v�Y�ї<�VE�#*HXD!�T�mU��§�RLXQ�I�0i�yl������[�]��껸]kQDGΥ�@c�Q�DoNa��AC���񟕘�Q�b ��m�+�]�A��6���y��)�a���O���f��0nk�w����$$eS�w���Qn������W�]�A�<��Y4tN1�;̹;[]_� ��E���P�Fk�
?P��;����o��=��$�·�a��U/3