��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jåا{�\�u�?߷�dn@6�zf��r������;g��Q�uG�ӂ}]����p�^��-�v�o�;H��j7�_�q9��{a�<ɶ���y�ˠɸ͏ށ��&�*G�� \����BQ��^���ܚ�dfk�
y�J2,7� �N����O�x��WMj�� 
s���SG�J� ��d,C/�^��M�rD�d睅��ץ,
RV�+���ǜ<��)��m�eaJ�<ɋE+!6�`i���tT�`�J�Kkίv燞b�ƚrQ��Ǝ�]�&�l�	�R+��}��ǧ3�{�P����T;����v��d}Jcq�� ���w�����ۍ�Ē�	�eHa��p�E.�g�������BK�� ��(�ۯekcи�/�Ơ���w�R�Yzy����J���p���uUN.���;Y�I8��s���c���h�*�k���vu"�d��?���BĽ��ofh��q����
����?F�;�]t�cn���]6�5"�W5U����V����*g�oq�q&� w��a�.RV�%bpk��>}��>�_�r?��,��ލn��b6*?�`4u_�����nn~�r� ��rL���1u��#1L�钴�N'd���Z� �R���ۘɸԡ���B8������:�qt�N� p�J�:]��R��H�Z���/LJ��&�̾څ�PJ��j|�z,US0)���sav�{��Z`R�{�P+�OM���5#zM'��;s)��*�Z8��9��2�l�X�.0���W��!�"�}�K3���J	n����&=���9��T�� �"_ݬ<�u���l潵�m�����D@�냒om�È!w{3���3�\/9(� ��K�����B�)�Q+n3�2��ۉ���,n&S���a���/����^��/?�g�x[��o=q5��gث�d� 6�����S��ւ�f&J�q$�R�3�Y�v�������yI��{f=���O�8L���Mu���:���]~u�Y8r�+W|��'^PX�x�N��o�.�u|L�k���j�=\�7"����0WN�tK\��5�2�,��k�wx���r2Duh�fG@ӽ��l_m�B���2����6�j��Z���n�Y Y��7�{'�j�Y�`�2�p����
��mzl4�z�$��l��x���yb5@�7�+w�C����Q�N��T���-{ȇ_v�=��hK����9���������%����_�K�%Q^x�G��.a�L�g>��!�H/���U\��T��������xƈ~�9T���h4P�|��g>9��i�m�.�Y��
mz���7a8U���%���Hn��@�W�ӕ$��h�c#+�Ȥ\��juX#���O���rV�e��w���;�)���R�y>:Q�T�Ք�Q#j�qѸ���+��w�1�~�{G�e��J�M�Yš���-�r1�h�A�͛�|8�#������扪XN?�3%^�8���T1�t�<8C��I%ha��pܸ�H��EY+�]n˲<��|\T�A7�=���+�l�㟖�f��b�q�z���
���d[�F��|U|(]��=���l8ۿ�;������O�@M��	�CG-a
]�iڽ�����f�����U	����#���CN_�W_�(C�J��\�X�#*�Ʉ���$�N����#����N���[�<Q*`�lM��]]���8�̅�:����`�F�(!���waY�w��X��&r��c�j�Ϲ�n�AtE�ܰ�F�Q>�4�gO���0���%�F"�va��2@�4Y5O�
�F%��Ԯ�IҪ)4n�P׍ ���;�D�[�1D���L8��\R�/�S��i/�=7v8�0�3Ά�Nk(~�e2�E�Ad�������m���e��F��-���&��9V��]��؉]����_���Ó�2�2�U� ��kq�[u�S���xe�hb�t�q��ТB&���D���8(@�\����D�
�p�����0�+�j���eL�2�fl�s�Eπ� @HW�?o��V��1���> �{9�CZ�(�Oe��m�����@�o!�ZW�����b���Ċ��@)5��4��к!Vװ�����Up��a��v���V��);�b*���{�C�.s6:T䢆@r'u�؍9,6����&�i�Kl+�C���4��g̦o	K�C�>�W?���mIW����;F5K3L5�{p��䜐�t8_
�6����z	�gn%�bR��M_�r���:=+����CY�A�h5���2+
��n��l�ͬ��H��)��Ԝ�gj��"�<��M�l!^rR�v$��R��9�S7wM��c�R|�h
����XeU�#4��Kr84��zJ�0������҃���B=&��}ĥ�����ԩ�(,�g��
�q�Q.��[����B)��&-��^�F� ��:wd��#�a�a۱�}���8燈�- Δ�4�0~�]��P���E捬M4���R�+	����݊=OJ�;0w��l���=X_��p"�	�M�)��F��C��|�^�z3��{����7�����թ�F��S���U_�����'�\�����FS�-g^�=��{�Ix�U=Qt��Fg�;0c�������~�/ʩN��K�����{dX��!��N+�v��׳�����<��L�8�lض��Y�]�0�&c�c��Sh'S2@�x� �����g����v;�p Dw�j�3e8TIy��������f�	,d��9Bq��9���D����_i���Z�/^����� I!-i7�S��+�g=d=���4ekL�^Y~E�+��G��׈�@q�
M��;B*	��[�9W&z��"c���T
�En�[Y�>�(u�B
k1��J�8]r��:�x��밾�AU��FW�B�Xk׮����튑��?�������ϲ<�����"z��@���]Y,��gWb�j�����=��Hk��ҔIC��$Z��)�>���ذ�����6�W۳E���Y�P��� ���*#���ʏslb�� �l��D<����Ʊ'��d~���$B̷տ�[�{�RRVփi��r���~���F�;n%�t	�������hr�²����0�=m.v���	+���0줇X�/�6��������)�BҍѝR[ �}��Z-��).�+������Uy����iL9
�!�52'�hýEԭ2�"�0�8�gh�3~��1^k���2�;�;s$+�}IG�@e��Ƽ�XOp��l��Ġ�� _�wq��¹^^�'�Z���^�6|%,����9q������\.�򎛘O��X��;���Nƫ�_�'e��O�g�8�Y4���N5��0�D� 2~L�Yj�
B��F���I�̵�@�+�9kyl��PM fs��R#0.
¼WC��������"��^#���8zg�`�U�4B��!�y^MU]�+��owSS�=�
����K��̂�E]���rU ��p���F�a���l��β7U,��d/-W¬t��pDqGuS$��
K-@����Dܹq���k�!C8�t�����:9�(����&����Q&��c���X�Ky��j�E�}A�5�,ˈ�!]�Ҷ�0�b���X�ۭb����D�.�7�2�B�o��T��'�F����M�E�H]�|�Eq^���2.�0���
�6D�N��N��6��M��9eF��;���(���pZ �<���d2q�}+k_���В���5[�2�*�1�I��_��k���z�z���=b�c}B��X�?bT��\68Ԕ'_�QOҞ�$���8��Ѭ�^;4��Ϧ��Y$�f�G��< ]�BN>�А:{���>���œ���Q�Š�W��x�D	��-)�3�:�0��S� �����$T�	�]0i߻�>0mu����zh���ع�˺�<|�ݕLC��/N�D�n��'ig�is���{T�𶨁#�(��`XI�Gm�3[����B_�"�>�"���:e�W�+c�Qf������J�g�t�kPnԩ�g�hl#���tJ��Je��ʀTK6�_��|��ƫg�ي�^Uf�3����Y���ߘ>_!],�$��J#/Q�*>��4��_��ch�&�|R��TXa�@�].�`ϵPE��<�:�Qk��ԩ����t������5-\<Y.=&�{�`�����X`�ʎ��O�
Kbv�N�Hl��	F����I�i;r�0QB)H�g�MsP�*�d�R�qS;;�Aʒ'�o�u�	�T�W�k3vI&fd�W��=Iv�ќ�֍�H��ַ|��SՇʔo����g���癉�:H,�`{�H[ X	Wk�ьI>\tPP���	�e��?�k�,k�Ӧ�t���=A$@T���(���ܪ3�0�vw1��x�ԸT��I��^ecN����,��8U�����Kl�z8�W�CW�����y\)��B����z�fؙ[�1,�F{��B�\M���G��0�&�K(P��OF�}_��a��<o�����q�R�w:V����P��:"�Ȩ�=��D�}'�R�û��r��{?]��o	�R)V��Ú�9�e�Nۜ���_̙Vrf�H<I�R��+||�N�)Rk�X (�ɖ�"a�����y�u�A��<�FF�נ�-F-W���sh�#��G���q���lއ����o�q-U�ӻ���+�2ƀ�-����Y�q}�G�'3-3�IuӺ���H,��ΌY�=&��gA29ҀT֦/6��V��t..m:?��|CVO��EX&o-Ӥa� 8�+9N�]����L.D���sr�j��{!�C������@����ڭ�Gh�+eE�5,:Ѝ=�x2�Ulom�1�Th��e'l��ad-�?:�r�̆(HD:c�ry���j��lڳH��%��08-N�ٕ�^�u�8�rp���tJ�"����@�Ym�H��TЈ-�,�"w��ߠ���/6�=MO��0kY����]�������H��٘!�[�K�S����{҉�~��ݪgUh+7F+F�FL��8*(r��d=�0��'v�|�߳/�9��]��ws���{s����h 1x��������'�r��6��5�����36��V��(�<u%μ7W
�[; ����ac_�J뷖E�_LE��Б>�1�[�ՍY~O����AH>��3N��#6�CS��&d��_f:�w�ݺ)�M�e��V'��ن�P_M���[)�?N| ���	Alx��E7�M�09����fp��̈́���U1=���T��0����:����]� p�U���۷7}���+j��CRxِ붻���I��G��h�b���4]�H_k���*1��a�^n=�������<�L�+�r3`�Y���I�Z!�k�{==���C4��]H�b��J��6���=�!�����@)a��o��#��%�BQs4�N�1���E[,ɪ �GQ��?_��y@�cY���M�bq��&�&�P�_;$���ڵ�������m$nX7�͊O�\Xl����M��O@:#`�T��&���W�W�o��xC��_G���/Dc�D2u�aTF��������&�GsS�B�ƠA!�c눨����piv�z�V����)�ۻ(�eV�
�7�H�$Mj.�'۪�݅mʇĜ-~�&���C1:`A裄~8�Oo�;�Sr�`<Ji��s3��\���]��ڸ����|�Y�F/�(p��x�0�F�'�d�K�]��'/��Ƙ�T�$㯜������q�Y��ӆ=`6r}��7&G|&��>�A&����R����(��N�r��hY��ڐPb$���(:��.n���9i.�^BGz��纎�^楓��P�T����E��謒��u�O6���!�_f�c��c��s��̶��Mكh1$
ja-��u�zV�n�G��rqzs7���̑�1���LT��84wy1WE�5���$���U/s`�Ű/��*147��_X cq�杜!+�e.��`�TC�ak���\Je��߮F>�b%��Q���5��=�������6G`�[��` ��2�;�=i��ϗݧ�/�m�h��i�.��+$4�ujq_��5�Q�����ho��3�#����!�o����;� �寇</[/�T3���8x!�<X�K�D?���T��u��V�� .�cw!��!�Wj\�3u/�Vҙ���P~�����	� �[?˂^�*@�7�/N�*�$���Z�Pٲq4:6@[ �l����U���_���\S���#�C������/ tC��֑4�2�}��6w�e��y1�
_�\(>��+h�����ih�	B�(�0pt�`�˳l`}#�y��u��
�(����ӄ��E;&�E� f-| ���1N�Y:N���]ط�-ω��h}LF��yW�+��wk��U'�Ϗٜ*�u���(:\����d��
�[��M��x��@����ݿ��H�ʏj1xc;���i��V�A}��,5z"	{tL�
��kx�c]ώ�y�	X��U�#�ֽ�[�ؾ�3Ԁ�=��ӌ�^n���2�f���ֱ"#�10���̭�����p͞�%��kd���0�?��� �ŝ�0X9Jr��,~a+��y��M_7�_��-Y�vS�uh��%�/�;U~ߊC*t�҇�t�k��z�n_���x��Ɣm.��>��J^�I 
V j�Ke���j�+����?���V"� �'vTf'���z��`�]LϠp���q�vv/�-�����?��n�T�	��ʈ���(��9B"��VX���ma���b�Ԛ�$�C�`"�4ǈq�I��Wrȁ��0f�[**:�����-�QJh���W�Hf�����s�Ax5�R�%�BDLGߗt������h-���/��]��ޭL�=M�,��m��ʕ�U�^[�9�o�C�[
��A�n���]�?�4���V�|I:Y�v�z+�t��^�د����(:�×C��	�.��v��B���S��A\�Q�Fxo0n+�y5�͗�o�p����}GݎDz����=����i�tO�7�y�������W�
M(hF���s{��7��� ��@W�=�${o�_�ĵ���~�A&}��"/��"Y.���9�ӏ�G�f�cߦ����-C�QbD�G$΍й������~Ԯ6��p����Y�EtT�RFεOf��h��k��zW}؀��ڭ��~'��EƤRQ;p�Bi*D�[��1#a�����豽�EKa���9�U�V�y��Nh�9�\��vs�y9��3`6�ޕ����	�[ܯ�(�&u&0)U�������A}��sO���?�n��u� ����=�4�|}���;����W��-��*;��F���m���R
���K©V�[��B�V䏣��PT�T}��yA�CAy���Xƈf����	�H�e���(�B��kO�$3�0�on�ௗ�䱘�y��1@�W2O�D����8S)ͳ7�F� Yw`|1�H�w�#�T�q�B��H1������9�S-e�K���~�%������K�E?�@]��E՛�,/pe�\�3�z����Wmcm�T���'�E+p� ��,|�ËH�������8l]MVȌ�������YL	a���i&=��K�=�����z2�m��x��}|26���e#�`m���	L��k����������q`d"����v_+��<9U?����Y�(P�(&H�2,S>�� ���H*ݻB� ��j6Sr�C������ύ��Hab4�3N�j'��2f�Go�a�O�z+j3�0�����=9q����%���f�f@m�����?U�qt�(8��Ƥv���B����>��c��&㍃SN5��6W;�l��hx�r��j!-J��H�,���&��(�N-ʒ%� &�zG�Zg�[E?܋"�A��ଛeG?�����m�4��T���GA���������)䤭���f	J����V�_�'1ou�4TK��*6�`c��_�$�,{א̗�.��ct�%��q����}i��ΐsS&0+d�{�]��]D�ѫ1m�U����U%a�f͡�t]��u�4��b�$^��cE�\���[�������~��}zb�M�W���b�ۚu�v.Ń�^���'��N���K�*f�'�#d����n�i�	��� _��3���_C�Ն�Ŧ7�-�Ј�Wc�"Ēe ��B��3GٰU*V�V7���������.O��H����k�� M�'^�*���?��w_��=�C�2���@p��5��La�-��� -0#e�&,4t�w\�y����7�p�
A��%:��jJ���_��q�1� 1��f�5�*��gq mO3x=��H�2�HE�!��.����g]���Ewy�-�[b���E�b��@��`����|����	rv&�^���T��]�RF�w/����g"G�
��?��R�r7�QX���r?��#,<;���["�ة�m�o ����ǊK��Kx�X�<�:#��nsm}"w�G�FW���;Ք��g���@����m"蓊�AC�Ɂ�-�Gvc�>6�j�z
��įe5�!B������z�Բ����Ϊ��������Ȃ��-���\U̯�zkL���B�K��۝^D��v��j�K�
��l>���r�S}Ԝ�U��G�/5��ؖ���G�Ki�v�8N��d����NCШ��,���02���������cJQ�c�W!9�"녚:�`�%��Ɲg��*�7m'8�j�4���y/'po�=�Et�3LLF%5>b�ѹ����/�B5_(�
�<Y�;5k�D}a&�%���zbB�Jv&�rU�$�!>�2C�*���N�ʤ�Bq*f����ۑ�"�n47���ʁ�8��ݸ�i��P<�^���T���)��7!�.DS|�]�~�ǚ��B�U�˧�@Ў@�5m�9�Z��3��ӓ���h�l��Ä�t�q �Z缾够�F�1� ��t��	��HO����H{��/�5#�%$֎�Jb%77� �z������ ���h�2�+��}<,�{��y?N�H�0�c��D�ׄˊ�gi�}e�h��U#�I���̊�4pe�i&,Ο�_x�W:�Xd�����zq�yY���c��&�9��J���>Z�I�����d����@W��&K#��\��^���֙�8wD`A�o�K~s�w�@���� ��A$��Dkgz���`�7��Ȇ�o!ޙ���D@�>�Te2b+����a����ɩ��]�4&��k�/W>�J�@)�J��/���g���,��MDWg�x��������"�/���&�3KP�:bbΛ�DW>�c҆�?�{�	�m�2=]k%L�����-_
�����t�$1<(����̱V�Tj�{�3Y:�w4q��_Ns�Z�(�I���tX<�E|��J��kq�6�mM�������� ����i���bR���K�7��$%Դں
���	\�L3�7�%~����������|�Y�+9sBve?���6͑qw~N�s\L�׳)��'z�ߚ3 ��3Tοb��g��Qc��Ɲ;��w輮?���Q��,�Ju<��&:/`]ǋCl$���|U�巟��HH��T���ڑH,�E�9��L�>B�c.���.mT7"�p<�kL�QY)V�C���jQW�_��q"l��
|�#G�e�ǚ�#��Ά��+a�95�Eb��V��Cv*zZ*��X�YG�	����/��S��R�
�7Z91���5��~��Ɂ�#1�ce_�*O!̳����y)��s�I4�f!�������,?Wy��.���O[�'��Φ��"b9�Q��R�Ȏ�W�C�o'�C��u��Ն%��A�,dX��D͖��Ds�^�0�p�����i��F~H���[���\H��Jl�<Z�\�ч�J���^�ոV�_����}�
�-��0��Υ�� !���zp�_����o+`=1�h��}�w�~"��͡�ޡt���noVʛV���;S?J�ɠy�d����H��^���:��;s��k}夒ܛ�� ����J8�D�0f�aq#�c�ئ;��Y�3d`���l�_�/�6țM�暜ê+e�'!�cL�J�]�������n�s�+^�x(�Zk\N�0����e��A������O��ie&��N��((�����'Kg�u8{���:���X�L�V�*B����V�$�n��V�@�r�q؊���J+izoD�ЬC~�����2&�9��Q ���k�&-����3���{B֦ܷ��<3]r�ˮ���+v:���K�{;n�f^��	����3�^7��ؗl]7U/�rG3����ѐԨ�����K��sc�����]�-:�QXK+��~��|SF������������u�Nf������a�ԝ�E���O	���\6Jgdm�bgw���M�3N,訬��1��p�h$$c.TN�(|%����l�ޠz>��PQ�������L�����/���8��DὛ2�^��᱔�Q/J��y����
�XS��4��]g��( .3�شt"t���Ë�����.Թ��%�g�H*�w��5�pɏ�Qo'��P��%�8xX�g�p悢��u��no,H��U��� �\狯�M2.��]�.[�zAn,s��Z ��ue��w|J9s_���0���ݚ~zY���uK"�P�B���}S$��.�(���z7P7�׬�y�)b��Pu���)_)1#U(I����{�qu\f&a��Q���d��B�^�I

p�+�*��~���#N�o��;�c�v��e}M7 ��iA���)��ф?�&%E�������Aj�P?�-J����O@ڌ�Q�:%�;l����V�x����"GN��׿��������|�Tr�����V=��;����?6�1QpЄ������OTI�2�#���sKp��8�&Z��̣z.+/����g�6�PuLȶ�$����U�تlQ+��h����pV��qU�ݏh�J��9�����	v� F3
��3���/w���aIh�E6,� �KG�G]u��y1[���׭U��M`��6h�:>x�=<[x93|Q�5�N�jo����TI�'���?�wP?����T	�C	�K�df�.b���Fu",ci��ܴ�!^�!���՟�6:gF/�����Z���h�㍀N�R\:�#���i���M<�����pg�ΊDE_����؇j��0Ұ9=��ᘵq�	�k�$cЍP�O���4���)��ߐu �����*
�P�]�D�8�b��A-����U����~�ZX��s:�� h�{/�8�f�DP�%����՛#��G]�]k!����[L"p)������AMp�m=#��|�7~җ��[>��N��=,�A�ʈ��Dń�}���Wi�����a�晻qα:�5$-J"Q ,�*2OA�hF`헗lHj�����29�����T�6��M73y���wc\2� hQme�T�W.��k�J��bn�f�&��g�K.V�Q�����9J����zSr�"�9(?�fw���r."Lvnk�n����(̉��2G�E�[�;8�*/V��p3�>��q����3$����Z C�pT{8��.í�*�3��^B�r�,�B��7zf��A���+{�di��JuD9���ˁ�M�ɑ/L��s�xc�SZZ���
	>V`���N�I��e�MOќg����<ix�x"|/�g3:s�|O�b
�<��h��K��42��1f��)�C�l����z�[S?�<kL�35�r����7�f������繊�2p	s�G�w��l��`���F�r. ��kS�������<�~��kS&M3��$#1/��4b����C�Kj���]a��c+Y1��������.b �*M�f��Dm.Z8�P��a��v��Z�L6������L�[�'��IN��J��y�|�v1�^�<�]�A����,��3?s�Q ߽��:ק���\%d�f�I�k��Q�~ڶF��s�����]�Еg� Y�#@ �Czn#�<ї��m��$w���=@֢fm:9@�L���
����]H����P�W/\���6��p�.�A���0�qBt�{q�:GP����;Cl��Vࡉp8I��Bz�*���"�P
Bb)�����>�wn��yH�7��Ҫ��Ԓ�,"�0�>��Թ�St�p">�*nTk�(�9�3F)ҭ��2�VRe�PN.L�m���u�e���_������)x��ka\SD�)������a��NcvE�z���|8<p��&e�X�~Ρ�2�G�UsA�1��'��8�j�m�<P2vC�u���]&���IIϛg�o-�pۆUZ)��+�*>�R>����>���9�Z-7䅘�#�y��Gn���ՃfG�j��/�~�X�~�{G���V�JO]�� ����+��xƅY�+Q�2zF'�s�M
�9�ϱ	.
&���{m�J|��-D�ƞ���p���ƺ����Pt�cD �Ĳ�*�Gӄ�V��=�Y򡬟��g'�up���Qo*�fK�)�G{�}=
9�˭��:Mo�r����2�,�^H������bTd)|A==�o�{+��_�K����!8�J��v4Z��\6�Di�~�9gp�Uԡ��Z r/Pu3m�O4f܅O�an�i6�yW^ϩ�	V�E���|�Q]�e�(��6�hY�v뿕�yÖguE:��ʸ�?"X%$g�b��tb�#l���w5~�Sm�MՊ�������c���ȟV�<�I�h$�ύ,�e@[}�Mq�_(]���z8�Z �M�����u�ݱܘ�gT�dY�y��P�GX|!��S��Ƭ�$��ED0�;o��~~i<BՇ��_li��:���0P�I���t��������Хv5L�˶���P���V�^��Jc��09�%Nv%< (��i6�S7��yK�j��(}N1Q���P�	 �����E�I!"���X��)��V�z���&���"G!v1���b�I�p��s���'�m�@p�3�|Ġ�Ԛ�T�� @�����~��;	�p��j�#�x��\9E�����TZ/>�}c��<�bM�9��ϙ�u��l���v8"2v��MD�s������%�>\�s������z��*�M&��҂�n��;d
�Q4k�Jm����#C�r�#Fg<�#?��4���z�x�4����6���)��}7����n�F���C �v��j�t�w�;����Qt�u�?��"���WWٔu��Q�dh�|���0a��AF�u����2�����"���r�PG%�!��)O��H�b,�����W!\���;��D��o������t�4�4��ez��5�3�2�\�����	���zL�b�pA�+U5��C��F�#����c�]�� l�hzV¤�C�w�����C�#%ß��G"C��������+���n��x��̧��G�b��k+��:� 8t��0�]�[�����t��j��5�"�ow0�D�'@~�\r�XA��論S�c�"��Г�E9�}@�����R����BA��O�o��g8�I7T����5�u��s-z�Q:��X\��k)�YP�1���?�9^���ɚ���uɹ�)!�(	->J�-zxVQȳT��6)�f^}�������c�qP6���I�Pm�x�dĠ��$k%5�wZ�`%co耄��pW`�"�_���FL�4m�0����_|����ƺ�xj}��,ݥ>��ʳʨ�e&�;�oO���w��ϝ��=鈠W���ځ�z@�������3�L��J�&�la���P���Z����M��g�]O�P���힦ފ}e�� �����h\%�1��u��U����RaL��7I����DrM��#c�e�q�:&�[d�{�����B����̗�,#4���l�c��e󋦗zc��+�v:c�%�����@R����V�n���/XM�����������X�)��qlM�o��r9�n%���zTc�솊�>B���)خu*'�s>��R�!m�;�.b�V�e>�^���T&�մ-���Z�>EhE���2XQ:.Ay{��?Y� �n.ҟ��U:Gi�����Os�/=���ϼb��?��c�w
*�pw8l̎��Jʳ
�ԞNT��}�u�C�izʠT��~D�)�'��B%8�	�Mx��	s�#_=�D�<;,pu�Z���3.9��(���C�N����N���@�y��
lV՟�'��9x+В�3�����ov3���b�a��� ����Z��m�+q{,��=V��
�]�o�A��n�(��OL����9���m)S�ˀ�����������K���<��`�'̙�[�20*�b0�P�ՠ#�_ː[h��e60w��9e9__(�mF`mhC�N%?��k�Ⱥ�SP�f����,�8 �]g�_�+�bE�<�5��#3GyJF3�.X��˽(�+��}��*�c����?�uŤTA/�w(�O���3U^�. ユ��:�_�ć�@�Fpt��U��ז{���c@�}�ӧdW ��
�է���2��,T��	09�z�}B-���Ng���{I�Td�K�&&�N��[C��f���i	��(GV��|~1��yM��Jvz�3G<+�������E#�[�Ph��TA��ܭ��ׂu*�͎M�F;���H>h���܀0�����cj�cFz8*��=�m5������7�=���ݻG�}�y�q�'9pMN�\OE���_����h�B�� �(VI���g�\	%���|�<���]����D�,��1��72��J��p<C�s6��U�;���L�+L$g�x��z�!�����cH㪮d�7��ej�zXV-qC$E�HI�v��5�2g-D킷�6��|���Y�Z�háɟ��֡�"�3��rlx��kB��Ε�+��ݧ��mg�_��@�������֓&�D	�\%��4��J(�Ǭt�%J���?���ֵ�����S'��ǀZ��ج�?��J�#Z4�}���(�
Xr8+z�{_��1I�FG����ψM>L�kvDhc�| 1�;Ќq��p��OY�b�$�*�+��Ed�e2�4	ղ\^�^n	�:�� �����7K�̋�U������tV�2������-�O�/���R�u��X��\v_ ��0��M�1��8���@�#����掗�pW��!����$p�(;璖S�j=��?K��'��~u������%��)��vC��ɰ э�Qq��I�m ا���� hOD4γ-T��Ed-H&�sm���w4Ψ���Jc,�.���C؅�4�:�R߸��z�-{��G�����PWE��k�S-������!��7iS��x��Iь\B��[<IZn�Ed�
C�6O߾wh�Bx�>cY��|w��$���q�wfL�zƍ��-�5_�w�i��m-B��|�J7VX����7h��'HB����f_g�&â�f�2�4�y�_E�38{Ru%S7�<8�CH�F* k�[U�!/�$��!	T���̼�^�J]�[�^N>pvf���ŌΝB,�#f��`m�dfu�tH�-_�X=�ўA�3��5���f�ġg��.p����H����x���>f�E>�uJ�NsOF�C�Ƈ9~�����4^C��$�p�8%�*?���
�Q5����O�<�]��Tw�0 z3�0�S*:�_����J�}��>��'I�@7Hssh�)\�Ō�fc��8���)�	(�|�Gv�QJD0:�QWj�cs�R!����b��i�Yke��m�ڤ�q�w���s#Ƌ�S��r�%��p;o�2s�H����}������/TBqXp|���
�ub�8��G`}��z��
�j!��$��0�b�v����s��zZ}g�(�y~�R���["��f|��mņ���:Kp� �n0f���v�.ȯ�̯|���j ���|����&�H#����:����G��(z���?I4�l�jc+�t�M����٫J�3�*[����R�QSq�����6��@_݊Xw��^L��*�p�5��8�:
A���lg�֕��7w�ߏ�ɬ��
k)(e.��B H͇��3� \"��6�Z.�#Y��2�,�������W��N��ę��k�F�N��e��Ն�v�֑��O� �X��o����:}c�	j�.k��o�`4+� �"E�,��/8������vn��W�r�Z!��]�7, Q0�Rt��F���j�n�+�St��y�3T�x���E�Z�(K� F�d���&|=U�r�h�	E,�w>��J�Ir븕�zР��[N���)�[������5</�D.�g�ⵓ�EU�z<��W�Q0*��:��`#�*�v�c� �~oz��I�$��S�r��s���}�TK�s��>���KLI���@����.�\���՝s�1��W����fiɁ~���^)JObbAR�� �r4y:��1+9C�f]�ޜDe|�i�^q7���Z`�&偾��2����$Up�z,iE�!Y8�2*6nk�4+[���b���YD�M=v��v�V#O��?χ���Lgs���q�Uճ��.m����j�us<�e��79?�i�Ä�Q]�tZ��vDH8����t:�֖bx{
�@���c����E�۾�{�)���`�ٙ�nz
!�̼���8Wr�b_l
�z�4��w��@��#��"�r�Ŕ<{/nS�����`dd��8���!�ܴ�7�?����|w�v���kh��'��zz���8������-�@�Q����c"pX��J�.�R�:���JC6yZ"]�;w����fb��<�>��&�� Ձ��"�����%zXc��4ou7�ގq�HC-��2�-�H�g�U���̘�WBDsKFw�fE:����U��QvG��ƜN�8��D��z���zsj<<��D+.��T��f& ����A.���� E�܅�ӄ(�yǧjr�5���6btQ+���l��L/��iM��NT3�����@�/O�qK�t��+qM�p�s�jܺaw���`R���E�y���������S�;���j�ā�j*U�~�ԑ=/wv=0?�E�#+ja�����[g��@eN�(�|ˮi�����|E�6�r_�W�ޭM\L��T��V����ĢZ�3u�̸L��i�q�@��,���t:f�>x�R:¼�D$���t>t�E���S�8t1!����~���d� ��vuS�����9�Tb�#2�ZI���1%ق��t���Y���f�E�H�ύ� [��'�⮼E�N��\��k<��²f=c'�_�R���״�U�?�@=|���4�C]~FL٣K����s;,[+���Uﳔ65����>�/>̨eG�~��6Ġ�����7�˔����/ �5qNb��!�'�Mi�IH����y�$
�\��M�0Z�d��a=��e���H��H����d�Q�w`�?�4]������Ov�x�xUg���e=�Z��fy����,]U����4Ů�y���V��\�_�^�JCG���
Y͎����-�G}[ڠ�	�ɣ}ٱŭ!ϣVz�J�t�.�� ���������:S��*"�jo����Y ��oee-3{Bp�z{MP�ӂ��'��1���3��}_aWt,ں�H⇿� ���V�!��c;C�
�pͭ�]^�<|���U��gW4�Ta2��<F)���!l��\��Tr�����I|������0��c@�^Vk����k���; �a�j�/AK���5<�ާ@�݆*ڔ��
��8�ㅑA�9m{~���;����[W�"h,��v��N:���=�Jl�6�ӕ&O)U@զ�cJ�5g���Z3��ۀ�H��$�,����9WB-RE`�7��y���F_/EHג��X���D�sJ\��!�	�����	�H�e)"�d�u�f/�/T�6�½�Ͳ�&�wRn��^��,�~%>���gW�vw]���0�Ա\h/b��J4���=��K+�\��Wb�ِp�����{T_�����^�\��W TD(�;�#Mw�ׄ�ub������D�:�<_ɒ^6DwϤ^J����%�G�}��Y杯'sA�a��n�!قx����̦�n�d�{���A.+�#��y6V ���{>p���rTlm�"4�`&�ٲ�,�R���C�~W�a��1N�����_�(u5�p7A�=7CU�
�5� �r׊����1����f��g����&P@8�_�T������r�T?6��B'�	��ǅ���T�:�����l��V�?>P0�KOt��RxA��*��$I:?�ՠ�~u�l@ĹG�*��&z���kЉ|yI��iD�	��7S�+���H���f�#,7�8U�7^�q�kuyN��������. ��[�Z��o����龷|�x�yG!��ƜGhK�������Z�n W�������H˼)�������?8OG=wׁQ�����'�.f���Bs<�F	���	�/$C85�*�C��q��%`
լh8�)iњ���+'͉jΤj=N�%(4�x]��nA�ї3��g����=�u^Q�����b�v�f`���B��r��˰fL���R�]���+�k`X$|Y������mH���`�`VX^jOr���,.L?��w��$Ԛ>�>M(�E����"2��ʑ�j)�� Yo?��� ����t�D��ӓNRDX��|��j��������	`����'�$eF	�\P�Y[��۪�ק������ ��ׅ����c`d�ɾL���F޾L�bS���dn�G��%�^.M$2�ؤ�Xx{G�+��K.�"@�n[/u}�xß���e/���v,a������s��`�1��]��;�@�
_�g�ٔ_G62��*W�w{�3̘c!�h=f��N!׾��qoА��5���iU�����l<p+�'�7�E���fMFL�Qw%�.`��q��,v��A��I)����h�ۡ����kU�A>U���~?�KM��8PK���q��xpF*��1]��.]
�f�@�l�GK�W�YГ�DB�_a�o3z�|�[�A��_I$�
+�������� Է�/ޒ@S^��
�fD�,�Ʉ0 �|�0�g��i���"D�TT>ٍ�t"����|ٵ��.m��u�q��/O�p�ު����g9�u=�ղ'uN1@�(�%�Nk��to���v���U�05,�v� ��'���#�0%`Ȼ�]o����X��6/��a�i�����A&=yTE\��"&x�� d�R�`H_�	\3l�@�7�V!�Q�!��?`�7����T�6�<T ��� 9�fC�}�8X�������� b��lʆƂ�=����_��"�]/�`ǰ<+�;��*��t�����g�&������Q���l�B���i7��∧��O/��6��$���A�v�Y& �d���n����%U�(��dVh�?�>a!8�J�r2���B9���;���e
�"F��l��<Y��C
��5%��ِ�H�����dsB���֌SPe80�ۜa!��b���+��툆���z�&��t�7�*�d�EK�-D@Av��H�{zp2u����t��{��HI<�Y<H=�2�z��*e�����pg���*����I���EV C�F��܌���F �
�����n ���BcD���a�U��D-��/V����LO=�j�/�-�a9�7T�rK�qx���:���A���JSI_�� S�;{obѕ��B��X��R���c'����hP�T����z���b����hRB?����n
x���3�Se�>���O�GEZ�� 4��O/��?+BDR�?�hE��ڱP�y��drv�����)���*��}��l�a�b�]�yg�2�V785��c^Wvu��
ż��J�$��ȑ��n�K�K�)WMLX�]T� ���gq�����Ѓu ���Q����e?�ؠiB��
nl��A[
����GD�hf���vJ�b�X3hu%�P5��1�Mё꾌zzh���u�K��vE�R��i�� #0΋<�@X3���]�bل�T�� ��8��m���Vv�1����8�f�h�(�z��A.�b���A����'X�#Y���J�<ou�C��ق3Y�&HFgI?!�N�q����I)yv��K�]{�x�`����j!�sW�9ô��w����E`�K�
�$��}{��|̼=���}tN	��q���.&W�:��<	ԡ��ˋ1/>�	���Î�%�u�R��
2P ���|?m2'����h}�$�e}�ƥ��F4	7������V�QBP��G����Ʃ��X��tjpIeDm��ߢcS�~�fҎ4V�o�B����SR���w%�u5�xۮ�>�߱)�I�dQ�b}�G]ݿ�4ZZ6� s[YL� �����Ό���	Wx������C~݃6{'S�ƜE�<�>|��/�F��On��˹Gz}�u�{;��'� �S��Q��\�BR�0��4���}t(�Uzj�1?��d6N���&�K��3�/v�\n�U׍�NTT�<�\�&H
h���&��}�T�� ��"�hjC:K;؀����D�}Rix�JFm;�>®�|p����/�
#��ûx��v�KOegr߄�,�6��>e���5r|�p�//E��i��hN��'o�
�EŲ�#dB'g��`p��|H�h�5^�J�
(1�X}�:�hm�-_Ə�ϖ�<܍N4rq�Z;��XG������7Fڕ����Vx���De ���$k%f�}1;##qw{���)�<.(��LV�/"�t���u��ؒ����h�]d�����4���{��S<�>X�l�g��c��t��m{qg�g�a�h��z���j����T�G��I?�qn]t��I�_-����9���N)-�X�s,�Wj����BFz3i����FG��LXH���
#��c����P��'*Z�JQ?d�fYc|M��b~۱N>�5G��S"憤4�4f�:�s���������s:� �4��C��ύ"��lv�z�������[˭*7Y&u
���}�9imݲ�kخ���g/�JT��Ko����2�(Ge��#ߢYe�|�ݙ�aJw�C���~����In}�	C�؃���1=���Á�;����)(�$��/�o�V���
P�WM�E���i64X �u��>�IDE� �������R	g��6�i���)�V��p�L�	ѵX]n� ]JA*�E@����7���6ʅA�(y%��'�*J���έ����kVM�ٶyU�U��f%��U�h��b�(���c����i���a��W�+<NV���'��_���ק�Z��m�l=�&�+b��tW��2T��?�
��?Ӯ�͋�d�%l��O> �s�~;�lKEZ�V�ʬ��|Ƙ)����Ȯ`��!oD=�7.�5Y�4��:ǚh�f���#�C��pR4*�;���2D�(�+�~����,�z_r͸.QDT���!��*�����!ń!�������rk���]İBd���˞<��<��s��������j�ױP�Z��!V�Hj��45U
LYZK�ZrH�{Fa�\��K�9Zty5l�F�~�4��v�ǘ}�����{�p_�����=j[]YX�ˍ��5D<-����0=���u^JPE��E��?�W�� -.U�ģ3���|Ul� �ҒE�	<�Ll����*�x�:���Wf��W�7�� ��1�`�w2ڐ+���:Y=�o�����a�HS�9��� �f*�+/�u�w��Cgȋ�~,������،� �I'0�e�ڪ�5@���۳_� /���Ja��݂R��3I@���2�5�;��r�іiw�HǘS��YIK	� ��7M���!t��C�n1�E�)6	]n���&�/��ߜn���"��*/�'0S	�� �Qߖ5B�so:���`qJ���K�(��n ��#�_iZ@�*��U�=�ˉ��[�p �3��[z:r'A�a�K3���+}�H�� �^����rj�&�j���p�2�*��txJL�G���牭b��q��5������R�Aư���l�)�~��Z\e8\-@~KQ�i�a��).è���aӶ�æ��Z���~�gVl�5�ӿO�E�1�R45�mn�C�]#G�￰{��]Q�D!8@���`t�@���l�ںP� 6�E�]��w���[�s�	� �}�#����K���WR��L���𓧐H�ɀGT��,\<4�Z��C��Ȗ9�nzff�u�����8��",Gbƌ�>�,���Q�p���s�YT``4RU�	�%(0�]}�/V�c������!\<�3���KB?a
�e��/��GM[.K)�(Rj߰�(U������Ie��9�1��?5�e��!Ҿ�}h�|�"o�L$���T�Xp� ���v�G\TD�l3KJ޶��B�Qܓ�V�
����Y�g��2b��y*��S�y_�y8��rS�x<A�~��2�;�2��wM�@?D�a�t�V�����:���vj|�3-��<f���!N:�Z����m�&^��D�6��M&�@���݇��L��8��̈e3#��Bc���_?d5v���qjQ�d��a,Q��lS,�Z�R����KY&�72�i��_��Y�I�b6����"��6|��,�^z�xe�%�JR��Th��o��>-�����}Z�
�T���Sfwޢ8E�)e6HO��};�q(w �ٙ~X?��m6�����4c���?���\�$�B��ָ�X�?:���h�����tS����=54��b�7��Re�$H<]z��a���N	L��L���N�-c�hk;�y����E#W�5GJ�\���:
~M���<��"ל��\QY�_������t�z��7��*S2.�O�̸ ��|u0�������u�E4��:�u� ��U��	[�� [n��������*��qE-[kmKCN ��k���=�0�4E��-ȂĠ�ӑ����­t
�₶��|.п���������ٵ��	���A�<��r" ]K�U��)Ҹ�?�św�l����
�Ĳ�.���bQ���Фh��լ�A{����b-N�WT�4�)}���9w����[7
�!��-Lڸ4p��36kd
�*����G�4�����r2�SX��{OAM$|"��5��б�0¾�4zm ���w,��r��4r����6l)^�İi���NC���Q8�������<bp�*B�S���v��|K�2j!0�W������� 瀪����!�%Xm�����S�e�|5��p@K�==�}�#5�{��� �I�Rx����( ;���jh[�3�{�w�L
�5���jGK��1���#poܳ�Ov>.W�����.�&�P��V�urf�K�ӭN��s��cE��*/�R�8��+S�d�7;�.�<�/H!{@V�����^��(���;`���Ʈ��u�+��
w,{tڻ#�K�����z�đ��o^E)֧L��8�����Ζw�T��N�ڣ�ŧ�����S؉U3�c������8gX+TFkQ�I�����8�Yj\�.gZ?at�7Ć�+`\�?�UGA��%)s�rd��\W̤�auG"}(Q��~����|� �hk�6�:/, �C���%b羊�ͅ��xqQy�cG�7�G�ӹ�J�a�D�d-<��n�v�$E
?�;~�k���K�$�A�����_���K�Bn��-�x)
+�"���/妣d�;�x��\f��}�0���\Zf�x�-�NMU�� �S�
�E����o)>`�;b�Ї���oS�I�{���:��撫��9r`5�_Y]I��QD�K�H�C�uױ�+ 31f�0|�7�O.k;�b����>��vq�{��`]d�d��*Q��0o:�D���J�w5��by˿�P3���^�錴%c-�T&���҂��p=��z��jP
�JIb�Z���Ro�~�RJ9�Ǡ����P�:�?.���1�;�F��|Ėh��|
:|��>4�+fF�HV�b!�<��f�Xà&�j�ԣ.�>Y=w6��Z��U����D�����+����'�3V�l�gU��aNjGv�>�G��ܦ���c�߂��'�]�zB_����B��D���J���%�:'�Y(_2oq~�,x�����P�+��������`�$�}���$��fda�E����=އ2��FR��U1vbM �T4�[��+T�b�c(��0]�B�d�9$�=�:���y�� ��%PӍ�չ�I��{bW��U|6ޛ���М�/FD,V+
��A?|��N�k}yX��s\����a<�@#��i�'�CA0�1���� jH+я�75���_(l��ͶG�o�
r]��)����u�������{�JV�l}ԡ�h�>^(��իR����0�7���k�u�%�� ��aW��b~D�v�+5&�~)����MIh��O� ��}�<w�w�Ѿd����E+QWj�s�I*��@w��[�zxʰ���ȝX0����=�\۪K4�B���+p��������R�Ԝc�ŹVӪ#FXa�2�'����;E������q/Q�*Og��6�g�-v�q��gA!����Z�*��(�z����4�߁h%���g�O�˯�������i.^��Qͤ8MsB:�cj�2|>����A�8�B��r�b?��r��c[��+��.o >��fpi>!�E��L��}�HY���� *,ܨbur��<#W:�o �Bz�z>4ܴ��=@;Iw�.h��=�'y��α� ��(��u�22ܯBf�4>��N��� �,W;���G�j�|ȝ#,b)OX������Z�����C~R�'M�`��V�>.lȻ�n�� ���M������\�� P)}�C���m{!��@��������\��a% ɜI����0Qu	K�W�;̇�@�Q,�Z���B��d��U(XV�yV���^l���#�pd2�Y[V���A6��1� ��-����M���cA��w�����o�=C��;�޹B{�r��T+���*W�>����h;�zb"z��/�0��1�&-GQ��sW�A��TOr�OQ���yD�0��Ub;t& �U�?��Of#���e�������h��N���Z�M�m���kv��`L��j�J�GG���+?Ā��H��f�2���CD��{�_���b@�3J�.��#��
b�n��T�fPWS�u5>��d$�����C=[s,Q9��S�dV|�M`�^���UzT�2lm�&����Rd�-6�����|%n����/�C���i��uX;�����;���F����$��͈7��Q.�y��^-����&-�! ��Ɇ�8�]��H��]�!�?ȏ]�{�l���y�ͮ(���e���V����}J������CY!2�`G�)��+��X��j?H���N�������Y�=��!j=�YƱ_k'�L�}���G����d`�U�]#���!*3�0+�K����%�ի5N����.:�m�Q�sPF�ou�X����CXw�
��[i6U�f�����2�S:�����͡�O�8�s,_S�z�Ts^X*�aM%�"qt<WY�,B��V�H{D<�n�/e�ƎAX洣UV�ȭ9R� f@�x�>���r�r3���������<����MN�0H�J�<�Q�5����
u��#�Z�lA>jE�;;�,�M�+�8uOK��ˤ���nisѥ/�s��h��v#LU��9����"�K��]��8��hO`�϶�:2X6U��Kb�p�W�����8�	��Z<�4���'~IPy6�_\h�Dq��"��z�{籤��|�'B8LwDU�����R!�SsF>�f���@��
P�Vgn�16���ɢY@� ��q�Uz\��$��U)!u��E`G�Z_��ӿ�u��6$p��_<��y�]�o���������� ��y����=���t���E���ci���ꘕX�x�v��-_��\���T��;�2�LHŝ�9Ai�r+2�Y�ι�Lh��[�4X��T��o]Ř]���k��/��e�Z������K���W�a���nG��A?�&�O��/�jz!�̫V��r;,_I}��_s5@.4��@Y��@���1>˄#��?����Vp"��˯��@&$�ˈ
9���#?Ū`�	����{C/?m�o�w��E���J�]���xiT�>�#r��9��{2}�Z�u탱2�T�I��t7=g��p�e?�`�Ht�w'L��|(QZ����hY:,�>*>��njQ��k*���s���JR*%g@z�}����V��C�j`a>m��ZQ�vC��xO[2)�LZb�I�������<�7���ح��������L�'�]�'��l{N�B����>�,�{$�cl����!����h$�������^����Ai��G�����3��� �:��lr�Ւ����|mu�F�n�.Ռ�p�8a�D����yxas����$s�A�V�EΕ{�,D�OT%�0���m�b��|��,;�U���,SUv�_̻�GJ�"FV��򧶵��n�(��B6�ss�58����0/�Z~�M��[?��ng)VX��"X)�1چx���T%�b)�7<̯e��S�i]��>����Z�j��(�i�@��8�����t�.rO$r����}�xY*
/��4����cb��zn=¢i6�Z��L~�n�Q�ϳq�y���~����q�w�}x
"��)�p���s4��M�[|�Z;O�};�v���V��-Z����xS�  ��)~�T�[j��+��U����P������z-y���e��������O��<���l�C!�c�v.�mDy�B~����F��i��?y*_�o#=?+bE�,�R0�n�ȸ���z���朾5�qx@�Ef��g�T��k�O�q����bx�]1��Zh�/1_�ײ�:^g2�<��1xaT+�d3�Jw�	�-)0[a{�c-����ӓ��f�z��$oCz� _��u�����O(u� ��x*ѐ��1쳛�-MirX|jE/ꫦZ�X��^f:�����:�i�bF7ǉ��Fs�Å	�	u��s�[��yW
�f���nO@���VU����	� ��_�\_16������ #�4B�Hc��)4��O~وؕ`�����p�"嚻��ت���o�F+��;�-�?�v�ܗ@ʂ@U����7�u K��a����;Ńԇ���>L<��gw?҇�d�@�ǾY�ս����¬Q��΂\��i��J���x�ʧz?��yM�25ze�?�9>�a��P���
P�0�-K��n�!b�K`�9d/t$�-�wSu��H'8HS&�?��|�e����E�Er�T�deW%#4�M����>���/���j�}ɜO�Wϴ.m'�T��P��������͏���B��D��}���	~s�.��JO���H+$�R��W+$
01�ŴC�<uĬ�+{Ar�pΪ�hZ*�ULƺ�2�<���ԯv���k�6T�g8�&��؁��:e�3�������\�o�q(�s�^��W��SCW�a m:�ި
Y�: �~!,F3eYs���/�Y���TS@��	v'N�6��Q�xG $��(,S{
x(��!µ���RH �?�`8��� ���{���v�[)�`F��!�f?5�݄�FU�F
�)u�{����[^��s��@�n�-B�<%���Cϊo��ؠ��,����>�"��W�27�z��Pk��Ĥl���ܺ:չW;ST�)E��,�����6�-��o-KS#E�0/�r�M�Iz=��ݰ�6�f.�>,[8���(�N���癞-��#���L��U��Ԑ<lu�h��\1��~���I��o��Ր��zE��N�j��$�N��]�^-��
�S$w�o�Ed@�ut��=�����5����{��謑>�Y�N�|+p#��5M�]nc�h��Ű]��YvM�:V������9�U��g�	���Z��z�A�EY_|�B�\�_�e{��>���c����&��Zh�݊�������}���'	8(�z� �B#p$�ʧG�%.�O,�n�6^�|8�6�d���)� ����tB��y�'������上�r��8"U�LtyQ�Ӿ�t�	O���鉓�s<L����!�h�t��0kjQ*���r4\Ho}9��~���~3�O�R���/���K�+�E���� S�����Ƽn��J�FK؅`/,�%.�sA&��8k�U�3�yw|���l+��l�����`�O1��PY�-1��pI�?b��`^��lN&�2zX��#�G��۲��vF7߿��)"���s�vox��+�t�5i*����o����=[�9���$��M��,�Q���(��� ��R���*ɚ��@�a~��=��Z����9��2������7��;����lN��J��sg�����o�E Dү�a�8�yN����E�TYVziOi?��ʸ�ၹ�^����.�r&�����:��>�t��^���a1�P�&*���g0Sl�C�4�}䂃IEƐ�mo9����������\%gD���}��Sr yM)�*|fh��������>��݌���6`��o��<n�j*NEC��!A�4z�Y����"�_ٻ����m3�	_��a�Պx��߫��
�fWKR&�+��&pqw���i3���=ͼ����=$	<䲨2c }ol}r�\X�pl�T#[�"��ŒK���cQ�C�|�"��C=�=��j��E{E}Z�a���p���c�!X�D=�&�d����|'#0H�r�'EA�1"6|G��,FIy63�%��%�\�n��[;kT�fA��(�#{E���%��]ptAI�T��2������t�^ D�Q��>�^ϊ�^JS���NWH��*���҇\5�ٗ��n\r���kn�H�4d5k�Ǯ���z;e�y�;�#|S�5x��|���ױ�N;i@�l�Z"b+����௚1ʘ�M�J��}<C���U�O�Go'����R��9�h;��w��<n�v��c|�U2̣q7n����~EYE�����D�����N{�O-׫����w��9�IK����d�|�!���j�{�7墒��!Zִ�5;�H_3�;d�/x��6'��e��{���`}���j���8�q�Of2�<�m�����;���Ѷ��א	l�a~�]�:(t�	nϫb6���c�//��r�*��+{Ρ��KW��SZ�,h�m��*�ַ���MP!+G{���l��\β"�p����4�YWj�Yʏ^Iơvr�L�s��y���M��+���T.�y�[S}8?R�G:���#j�
�ɧ���9��+�r�L��jI�H� ����v�!�\>\m �o5Q\����᯿�����|>%�����]*1�����5)�Xj5����WC��Q�d�>q1��]�, �P�Eѯ��=a䰿A�4����2L#�U��ܣ�1#z|�$mu�[��?|X�C5!���c_�I����UCWGĢ��I>ޭ{H}���Hju�'f~@a�����g�(t[��#O:9���QuB�����9��5�}�P���!�ڎ}�U�S�N�j��V�~�Ż�K!���(��N��t30��1o{��L{^4�%h�<f,WI���"�:0<k��	���5;�0�kʒjC�N��$|)�$��aSt�S&>��8 ֡7@�4�w�L�g�XbzЫLp��ˌ��1��q�Y���")F����o���toj� �ߪZY.�E�lU|��B�\�*��^՜T��gE�yR*9��B.��ݟS��i?��x{�_�}aP��)�V�����4�D,��۩�|ާ[7�/z�/����^�y��$kt[��&��L��)���vLO8�zR���ݚ�j�g�G����E���ǔ�o� ��2�h�5Ԙ�K�(1Q|�ô��v�b�!7�5��}��@�3��$�?������ό��:!.�7]'����?e�K�P_�M�iw�Q+�8��j)t%U�g1-]�"��� #�z#{b 2���k-���
1Q系��'+��G����9A��`��OL�6�@���@)*�f���h�E�|�PeJ�6��^ϑ�����l8��9�]7�F+'�O<b��z�/����d��6�0+�S�dm.wRR�`�������H�f5P�ɸ��k�JM�����%�%���`�;~�!0�����+F^K&��ԝ���R�����4������i\�=�T�P7YɃ�M$DȔW� ��.��!/D/��
�z6���A��)����
�u�ԫ��e@0H���dj���_f��U��U�S��+�m���������wA�d:�U�h&ӻ[BS�G2.���R��l�}��/uYY��� Gޤ�/D�͓������'t"+��ǖc��T���u� �^�YJ�,�Ca��ʺ�Đx�l�d2-��-�:je+��q�V{nUa#���J��ǩ~o�xL�����B�E����R�����`�xS�� *u����P�w{MƘ��"�[�b�$F
��-���oL���&`l�rcT?�L��I^9��X!Hϋuݐ�uZ(k6�7$?��r��p�YɭR��Q%g��(�|��6�׋�1���^��9�y���p����K�]����,��ז���p���z���*��'�+�>DK�Q�s�n��r{&\X��|�Q$�	v�@-�yu�H��uί�'�!�fiv3�k{ʥ���3�+��w�[n�G�Ov����dZ�G��u�G}*���j�}r�v���<ʛڍ�ӱ�|�?<R4�sg��B~&�ោ����g�`��?���0d{���a���"�`��˼s	Hv��}�pF�D柃8�T�i0����h}R%�)�S��zR�;�xƔABp��TZ�(9㣅5�M��V��o#J�9u��/&�N'NZޘ��4s�''18?X�i��h��%~�kE�����:̏�� R�������87�����3EA?NU�2��)YW�&[j�.&.ee�@	�x���W��ju��T蜰�k7�
�Zb�[�Dp9i"KG����p��b{��)�T�����i7�_Ew��>��f�`q��Iv��Σ��IA����a8d;���%	v�.�:%���2�Y��k!W�tt�u�h�`!�[�I^��?�=#���̮����if���MוU��2`��Md�qB�gi�CB/U1�P��[щ����A�AW��%�T�\��`?�0'�{g�'�0QƠbq���l̛�U�$Ǵ��bŚ������Uܬp��pޖ�'�r`V��ˉ�`飏S�i6��R��s��/�ަ���U�|�^ӌm+�J�����@9�Q�Bgvh:>`�҉
��Ebvm��W�~!��qe+rx�W|+m�4��J]��I�� �/���o����MP��MT�̿�fS����T	O�v�fwq� 5x�����;t\2��=zxa9��X�7�Z�
7���rq��X�\�u�4�,�w:�"��HvC����1��N?Mj!T��4*e~?:A����͑��0Ahg�D_�I�**?Ш���~���]	���ɍpi-�t����}MI`!Nx�'�]�1 :)øR^娌��@�3����8�a�����T��8��\�m�B7��QyB��"���k-��`�􀛪@������}H��E��E�o0B�L0�zP=^ﭽ2&_{*�����&��=���G���C��V	z��=��ztճE#6,@�NT㻳���{�9���#/���īJ��S����|{�Ԋ�y�C�vF�~c�C�G����$�y]�Fg�gLδ^��}JM�����~�ʗŤ�U���MrM�*�����e������ڵ	���a�� �R0>���	��s��_D��Ts����r���Y��s��82������^��Q�Ɨ	�m?d�;~��0J� �~���XM�}/��,{��=�#�5�d��0n�Sƙ���a�6F]���P^_��d�jw�#��~4�G�H;f���w�����kD5��+�.�hK�qmVj�+T�d4�妢1���+��TMq4�jF�(��	Si5Ղ�^Aё��2�6+�'`I$BWP�>Ae��Q�p�Iф��.Oa哴���P���
��Hm���R�]��0& R��QQ�fFBM�ZoB�[u��r�퐇�gI�����J���	6��؞��A�P�G��6���?���ye%��v.�x�"ȴ� ���
)D�+T�g<f�(V���cu��u���ec]B_��w^��P��y�=�f0L]2h~v=3��=iv�b.j�Rl�ȋ�÷%���{3���e*���+Mb��#��@X0�������q��/�&�ax(	$yX��phw�9��äMp�W�Z�Ro�-�w�yę�v�)@�ئ��󃍘��?򔕈6���k��h��A�"b��.u*w�Vd����U�R�)�4��Kđq�ҡ�ؕ��$+	R�S �YVyfVwƉs�K�{B	{�8��Zo��-�p>3g!ɥ�*���%�b!Փ�G��b�3Ŗ�.��&	���_���1+j�u給{�R��ۧ	��h�H���;�"�7+������><������L��߭�I�	��G�\���+��sA;�O2��G���;(���a�8{B�-���k7Vm
�,�v\G��փ��R3#43/�c���O:ǭ�d����F�;���~���gV�z�~t�XV��s/���rq�4!��M딟�<L����D�5K��0v���}���Ve�a�|Ee�4}�i�e�t���Nʍn~�D8���'K����s�7��M��n��'�0hUSb�lZ5�M��q�KQ\�L�������Lc����\�弫��~�a�-�xh��Dz�ꑩ'2���`rV��=f� V���/�Q)�T�澞{�_��3:"����2�?0#����`�Me���b�թ���~��h��t���+$2���#�+v�!\x�PE�q�YI���[� �gA�!�h��&�����.�I�A
�q��c�qa]�Q�a�Ҙ���ڻ�eN1�G2�ڂ�gi��2B�1��~�wk�HA;���0:|X�	\]kD�{��G������ To �r1��Y��?�HHQ���4���a1�����Q����X�x���У՞Tl�8ƣ�W�ΧdkAY%�=�8�٧86{��O�V�4 >d�m�!v�!�Hc���W��ZY� �	��W���;�ӄ.^�K������ȭ�^�����r��@�O�ښ詟���n�Ɉ4�u�c�5ʤ�K�5X5���ah�ȃ�sg�毰���YD�������a�^W����w�w��<��
��ێ�JkAP-���3�l��t��/�
\�18�-d3���G���z7�tխ<$���>��QN��uw�J�mt�5��F17�x�A|��LD��w�!�l��gKLʪF ��4L�4�������C8�c+>gݡ������i ����[���:�>P��jh��P ��zL
\��oi��������T�6*���ͥ��u�*��� ]�TS�d,��į�P��8��<��������\7V�q�X�,5v��.FW�xV�s��
�[g�DN�o��OZ�\Ih�a��&rWF<H������S k���G�h�@�>A�9[@c�J�Z
��1�vQ�􏃕M��M��ŕ�LHc�ovһjYK���M>E:·Ə�~VkVx[ܣ��yN�H�\b�.H@'e~��#�ŝU�������,-����rWGy���2?�����`O�;��k��Bv��~�P��Uh|����fC~n/�h�c��zJ�b{��5��0��h��X�=�o��P���Ú��S��������	�����Į b�T\�T�,4	��s:�%��m���<SU��`�x)G��f�lߟ����-h�W�6q��Z7����0
�Ȥj����'�?M>��~'D�o'u�j��+�=�~���_��<�q�[1h���I��R�>�B�w
yK ?�N�b��q0 �,�3�A��g���T���h}p=mE��v��̥x\m�HO�n�^/1�D�Ȁ���uL9CN�x� |A8QT�%�}����:[7)y�.���5*\���G���8Y�[���(nM�l`�r����9�I����[���G�N
�$7�Ē�11k��jq]2o_��I��vL����+�`]27B^�GƦ�lB��}�T?��OYXTy��� GG�F́č�b�c�%�oe�n@����]���Q�N�u�9)Ȋ��a�Y�ְ!���0�E��L�kNL�{�u#
����E�Ѻ������K����9p=R�Z�EA,&6I�]�C-m���	m����T�W���E�T<tJa�qtC�\?�:mI�QJA��n3�9t+�Y���~-�а,�F�Ud�`a��`����t���{���%"'�DJ@͔οU�6ˠ0.���n>�և;�`Z�\[�������B&(W�֮K[ן�܈(�L�1�� 	�4��P%'ߋ畭%<)(��M��J�i�e�J���ҍ�v�T��@�N6d��ᖠ(H!o��I�9L�?#�֠gkțC�?G�p�1�jى�q*k(c[qx4-`<9w����B<�It 3{[Z	��3�Xi34��|�O���j0����t�Xf;,��S�&�P�I߹��Q(�@!�9a{	�ep���������p^	����xSAW�UU�Uy#g��v�p/����/�x�^|a}:nS��eн�k���,M��f8��RP���2��?���Ig�����fA��e6������{:�#VM��ꏩ_�kZ��� ��?�X׭�������ˏ޽U���U����T��5����e~[���$�~�&�M��q7ԱcׇF_q7�?	kE����`��QS�@(�?�ا��vO42��Zu�ʨM�3��!6;M�*����J��2r@2��$���Ίϭ��j8yrE�B;�,*���d�3>�}�N�|#7$숩:�d�a�1���zWa��U��BϘ�������,T ��\���+b`��4p�q�Dp^��c�K_T���PN������,F�#r>��g�[;�f4�W:O�D�����c��h9��ζ.y0]�h�������G��C���d�|j%���y1�W�Ү}����e�oTv�|�p��	Y�RW�0�����0@���U�4��FRbA�K��s���~mÏ��]��	��'�[}'7p�	f�l�=</��jp��|�9��ڇT�j툛pL��Չ�6�+�ã x��P�,�dcf-y�T����ǷJ�lc��<��70|��<s������1���1��A�8��UQ@_t~�z
1~: dvv�1�.}�r!�+�m���ه)��_Yڨ�E<\y5�ć Ra�&Y4���*]e�,Q��ָun8�,�NҐ�W	����:��s�s�����L�w4+д��	����!��*zyj}a��<ݛ�O*z;��k�:fQ״������`T��1��Eƚg��	��:zY���;��
� �8��H*=�p���1��Qi6���*A����t}ʣ�z��i�����T�78��v���Ac��/*ǌ�,��1�ѻ���q6��o_A��]�?�w����cՄ�7atˌM-���E.Q S+@�MX��Ji�$Y30�����i30��)D��K��޿�7�E��I{�R�$���@��T���MnE�4	���YA} ��@t������{o�Z���͊�*�uU�(ou:�N8ڑ�,�{1{,���nj�c�zͳzJ�b�Q�s�d�2�]�sVS��+�о{5c$�f�2����KUX Vb�]{��� �B�7��}��l{AV��d��[��1�Hfy�Py0%��/F7h�MG�k��A	3�.���m����@>����(���e�h�~�m�xd�5�^+/-x���:n���E~?{#�ZM�L
��FuI�#[(!Rj%l���[�j��Å�}C�g-,*���~�UÚI�� �,~H�6�T����>�,��R+"��^<��_�.����GB�W5�X-�9��_�V~��j$�F$���� 
�� ��>����=�3��FE�<`R!HLC��z�3|U;�V�y�7�Gݥt��lD螪Z�ޕ�0.8, �x�jkJ�������J|{p����ς��X*�}g�3���&�Z�qt����z v�k���at_)���]F\�P���g��QO�T�z;�(K!�q=u����G�#�8�b*��ќ\J�{��X�
4A�E�O�g�c���\e}��4��B[Q���hق���4��GE�יX!�o
�11�/�nb��5�\�V�r�@�f¢H�5��;eK�q� �_�A͑�/��[�M�V�W.ᾌ�G�5�X1���+��N'W��"�h�]��G'<1z�Wߧ����&+٤�߆"���*UT�_��	��ȇ���}��%���ck�޾Ǳ�%\�\OJ�� ���l��)�.��q��e�&,����;<Ae�!y �1����߻3���iF���)Y���)�}�m��<N�
�2�����!L[��aw]	�[#!\WAۧ�����9g�@��u�oWky��[��Jp$��r�������p_��T4%� _3�.pz�4@( �\�8 vׄ�;�C�i$v���)y�t�q0tkh#���ok����#/n]�ɝ�ly<cp�Κ��8����O�z��G���9�.�lf����<�gY��<�|:���ȕy!`m����V��ќ��jb"T*�Cy��P�I�)�N2����NH�v�뵌	���F��Ƙ����ec�+\AEQ�0�X�+uzM�`5�����R���5�ZV�4 ��FZ�ʫ>E�ޅ�{�1��؁�&���pu�o���Y�P.����%����R�؝ap����w�v�$���?�`�u��-0�����ƍ��C>q�
T�a]��[���hoz&�������"���<�O������RY�N�����TL�{ϸuw�j�~?'rsL��A�q�4=T�-S0֎�r���D�&*yD�������A䃙3�w,b�ϔ�J:��i\��t1���(�d`� c/�Z�Nq� cJ7�6�Z-V����iրm�;�%s�Ȝ0��ȱw������	ڏ����4Br�<���h��lDH7�i����7�-^�%�pU0Y� �ضg=x/���%o3�:��\�PW�T��X5�36�R
��MO9�Æ��������c9�h��@*-h^=���\��pi#U���
]�Z"�qk���I���R}Ġ��%�5';p���7)h��I��C�+G�7z��h;T��%e�I~S�햊��K�n���Pe^d �o�cI�ܟ��%O�ÛtP�����L�ʢ��iPhgLq���qٓ ���(і�|������M��H �����,ӑUy�6�[@�n�M�!D��
�~��b��>*��Z����wB�D(�4?���p̰��ݵ���=s����>錀\�`��f�r�U��{�[�'v���<�ߑL@-w�%OS���Q�{l����EB��� ����t,,��G,1��NY�
������I�_=��V<?�A⌱�5[���(#4;�|Zn>�/���{�V���s{"����d�ox�m�ŧ���(̡tş!�!���Szh�eO�
����U�,~P �'ڽNd��ŚpÔa[@j�t�m����=�������3z���8��?V��Y�"�m[>��N5����Ǹ6G�i�>@?��t�{�o�?)#�UU�ʄ��*� ]I
��� Fهf�R^�ߺ�@�O=�\b���HO�x��>	����1���@xw}Ѡt����Z��FE��j3N:JZ���|mz��!��	G�Q�'d��ĭIuL��:>�����+��ٜx����?t����"�F|.�i2�ϖ�`���Q`	c��Ց&�H}�=<g۝����{vP%}�]W�W2�Z��"_��9�U�������b1���L��	W?���i"��5Oٳ���=3����p"��҄�����n�:ps��*C�k%������B"5~��7�!���BBmі�"�3�**c�.:�v�LRp�ء�fׯ,��R��I�v�&U�|Rd�ͬ�oTA��Ixj�f:��u�/�,�v�֢�Ck���]W\KI�fW��GS
Ls^�H�( C	7H�n��r�$T�������ֽ�1���q!ξؼu:���{���(��H�����&,e�-�fg;0�4@I��q說 ��R#�%�V���#�W����U���ݛW�Z��8X�*JSA�������<�1cU����-���> e��<r���y�۩�&G�!T�Essɇl�K�兦�x��x��W��H�`[5�*���j�VK���N�S�Ͽ��|�zIs��� ����?p�<�>=68{f�a�?i���^��
���hv� cVlOemg���?�A�	�U�W��bnEryR�4��L0����pf��eY�'G�!߂�x����4bdM���]Ԣ1��g�>�-��55��`�N���Gљ��x������O�HW>h|p��jw֧N�a$�-9� ,j�� |�JB�Nuac��<�{&�����A��^�_l<��z(��Q��w`Y��=�6���x%�dY~��:%��B%zm���Oz�@�m��dH�
��EW��S)����,S ����`A��ei��B%����a�'�^Y6l�
��d���G�O4�ŋ��9���a��� t�����A H&��nt���k(���8O0��~W���K��c#��B@�f��6��/,���jJn�EF�Clb��0�{,�-�?%�I<uϻv��L����%���1����a2�C��nG�{��0-'?Y��l.�7� �T�M4i�E�e1���/��Fݹ�#o3B`ɬ��}�_�xA��1�`�OOR'I�������}(6� ܽ������NR�l�S!����'~��կ�.�k5U%��޾��ȓ�P� ��3�'E�hicx泇	
!N�u1��m��J�tZ�^����U�4#���ݞ�Ѻt2H�f�g�g�D��wO�������O��V����R-�[�ŋ�n{��"+�]?2?/���g��t7re?T�Ӭ@��~.�8�x�������A*A�Qd�oN��dJ���T�տj-��_H�-�Բ���{\�F��������g-�l��"3T\���̶;ΛO�{�F�����<�7^?]��O �T�k��2Y:�l
�Fxnzn8+���7'�c5�G�NS�(�%�>#e�UB��S�#.�3Wj�x���W\Y��͇ޠ�Xh���1�u���j�+�x���;&�c�!���.Nl�8ʯ]�[��˴�|Nz�p�(s�>tFC�b&��ֲ�,a��7��z�ў�� ���,�F�G_�V���LdV�"ԝ0@�}y�\�w(P/������%��{ܣ������(ﳵJ�w۰��^�,����	����Ck����% tH��Ǫ)��:�
Ù�%q3-:�od�1]��7 �?�a�=�R"�5�2���'E���u�@I�]ļ^�z]�R���&C�2��v�/y#�>�)��'
ioZ�&V�x[�lg.M��,��Qyv@̷U'|,�C��̠�Ux�\�3x'�O����1�IP@Qd�Im\�;7��;\����7[��w:����6Q���: �f%>oA�{Y���t'+=����!�z���(��
��;�Xҷm }�;�&di��h�vP8,��m�bt�V겆!k��������r��V.�ҼÑX\Ģ������<6gi�@��Se'6� �3��ީ�N�|�K#�zs�C��IԲ�1�ƣ
��anB��+!%p�@+���C�r�]Bqe���4�Y7%��I>�o8S�h�&�ò�1���?�4��a�q���}����r���Z��Z�&Cy�+�3��S��|��5�:r�c_�x~�S妶�_�^�s|T�4��w��0`�a�+�O�_,�V���FA���Cx!���q�F�c�4�v�l�Y�83	��8��t�J���x�(���Z%�ĵ�4 ���թ�ؚ�t����&�M�y�� F4B�fr�v/ǉ@