��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jåا{�\�u�?߷�dn@6�zf��r������;�O):�l��f_l�y�g�
�>-�5�67���&5���S���m��jڻ�f���:e�+�%ɔ�p��-�6M
� (HI�-,�p�;�A1]`��7�h���ٹټ�շsD"�$��A�K���A�t	ct���"��e����=v �-`_	CF��(�p�����^���1襸#�Dk����/]�䋹`��
92!�T�A� �gز��C�bm%�Em�Ap�v�� �J�ᇷ��N�RK'~i �>�i�r�h~A�=J�L��\�F]zMwO[mXl���3��q��1����1(/"�M>I��4R�cn�D}�~n_�Lh� ��6^�,M�xa�B��tr��c
T��G<Cۺ��$�ѕ�7�M�~k�4���ӕ�"E���BD4�̀hY�[��e�b�eXJEuֱ0����~�ǯ��[-�:��N��gr�������JP0�F斡H�-���{�%��Y��{���;��/� {c�?����H���S'�7����jP�sbu�����$Nj5+��'D�ȵ���[W�/��i�\Is�C��A%c;����ϣ��܍�\��є�9U��%ɴw��;��+W��{��Q�H��%�2��˼u�u4�g�֥��׍w���Z�H(���ly��s��9hDo��h`Z�o5�z�G�L �,������S`z{z��=l�[d�ʏ�U�8"=Z�n���8#Í��l����4n1X�fb��j���3ZH��#�M���3D��0�ȫLWp:���cK�ڟ��Α�}��܄���%�f�.p����d;�bǧТH���PN�������/��k
�ݥd̍�$�����U���<3����̪ȕ���ıo����M��x�t�i��c��`�S��c����g��F�9��1���,8g�.��� �ukȩr3��ȇ�G�Ʋ>�aù�(�t���}��p��GV��^N�ɖ�Y	=E/�0�������2K��몋χ�6|�`f�)[(�C���E�.��[���B�ē�˞bE�A�:�я/������"��pW�]?����sFvFJ�*��>�O��F�@Y�۵�a]1|�:�Q��hm'����&�c��M�UF
��ni�^��KhL�g��Շ�Q���}&F1��z��3�(�?���I���-*n*h�X��bɞ"�;	�Z��C��_���i�9�x����NJ�W*3�����\��r����%��cx8��]��P*a�[U���=�u���5�Dr;������GH2�t?ve��D�HdX����qX�0�H��z�=f�D�W^G02҃��eD�����d��:g����N#����7|��������6c���[V���Y�^�!Qz��	�i��s%�1X�K@��X��bLA����o"b�Ѳ0�Be�I�u�ʕa�an\�<� �:/�$S%^���k)�2}�1��Gf4\uC -eֽ������Y��g��\p�S`',���n�HG�#�jb3�'t�瑢��=�N�m����n��o�5[H�s/��t �WH	�*o}�8�I8�	|���>�>F�o7 �� ��j`�ݟ�����u
mp�N�}�����p;GhM[!��M�W5PJ�vt%�C���y��|��uY{�c��������jH�6t顩�qj�<��*ll��@����_��N!�q?5�!٬�����>6�����8SA�W����o4<wD�,DNn���͵6�\.�_�"|����YK:X8�y}�|eO�'�D�Zv�պ�0�'��D|�����Xji�Y���~
��|�Yp��"���I�Ш��Ȁ7]�pE���X�6,�����C������������N�s�[����䜠Z�˿������1�s�����D��eN�������i�$�p���<���kM{�Tb����e}���YM�S�L#1|^�I�ĭ���hu8�WiVY;�;���s�ŢL2+Y�,>6?v*ߠ������W�ZĿIj��%s������1t|�}�C"U��i��3�Zz�z�<ڃ�8\�#`nr�SDn8N���H0;�3J<��!��hЎ'�)��},oC����<�A�	%��OD�����>�;�̥]�B���IAfm�[�� ^�B�����s�{����z��o�Z��`�|��V���%�(;e�w�õ��TK�F`�S$% ��6h�]U�)�}V�(Ӭ��c/�o\�`��؞;cA��Aֻ��:#?ls�-��66�L���^R[4!]y�<�f�&���Z��#
u:T�@^C&�Q0�J�a⹶�$�o�0ɤ�]f���"#�Ȁ���c@V����"z�h<�O��˓-6M�=.���R�0��}V�6L׎�P�ì^�>��Z��I3�׮io=�-Y++y_���{�̚�����/�9z�-�B��T�#"LY�b��)T?��،��Z]�t�%,CR�������-��Z�;;�hq���4��uMǦ ��=��O*���z��P2g>4y��3z��RlS�DM��^�f9���*����)�~8��������;��9y��V0�?FL�i�c��ۭs������x���$VT����Y���^g�ԡ�&�|X�F���Źb���D��@���B��h���R���[�l�8n��M��m-er�j�Ώ�\�KѾwT/��
*aS^��~����!�5k1�}x�k<���"M���~y�k����r�G>a�h��<�TN�
�C9�&����"�u��->WH���7�),s��"YŹ��Qi��gƻ^:� C�Y4= +al }#��1^�ゃh
N�lEsIe$*��U��_��@ }GC���4U�V�o�Рu�t/�s�]�$�]a=�YC�	��.���@ ��yO����-���
8-�ᗮ������:>�<�ɕ8���)�	�����$-�E��(9�ӷ�H0�${:�&��*uD�ր�K���}<a�лQ�z��]��^H]حzL�9Ĩ|/y���&��-z�6ߴ��C���}1�zD����nG*���i������d����􄃖m�����3\��XFd���䞽���,��ǵ�_<f�G�qQ�
��ժ ����Ž?Ѥ�wi	�[��k�z������I|��_���2��=�y��5cR�̰$�a���+I�닽 u(���Z9�6L��PT���y����F	�������� ��^��/��#�Y�>g���s%2�{G�[<�$�!�Fh���Q.r��0w�UH�_Z�Ή�N��4����r���촱��ڨF����|�������C<th��nI�Z�m�r���@&C�3�d�'�G��Oc��Գ���M���u0[�����x����kd������.~�~a�UGՈ��Y̷$�_<}Q��lӠs���-U�Q�}�g3{-ʸ�$��3�E�� au��^��?M�Q�MbSi��Qz�Ƀ�F.&�5��;ȝE�؉��)�J��3�����Yz�!�4�b:��B��rZN��j����?��V��o�7����?/�j%#�v�s'0�yX�1:�~�[aS٥ȭ{�sO�ȍ����la��y��H]���Ԧ|ۀ>��\�����QL�4
7{�^s���]�!
���@�)3���	������^y��ŚTt�]0���Х���H��M�&4������bxY��T�u�����L:�z���E&�/fw:�}8|�O����x ��ğ/�E�J��t��R��`|�ۨ��"���,ϯ���.!E�*I^�B9W�y�#�����Ҷ��j��˽�Ȩ�~ʷ �r_k�5��:^�|B�G�<:�	������*�&ζX��ݪ��c�OV�.���^���>�뿫�J��j��+�݆%�kr���u����W~-D�m�і���3o}Zv;�1�vn�uj���r�D�_b�@Z8�8�Z���Q�(�c3^�}P�� 	X�S��K{�.rQR�Ҍ	[9$���ƨ����,��_z<m;���+��=�bN�W�V��]r��,��l`B��E���>I�P���A�.�i����#V�v?�`��5�a�}��E�����.�m�B86��o3��)�W�!��3wڲ��A��ё�ݭE��]^���B����(+&��^`��;C�ǯ�D!k\r? z�m�/��
�.Z!���c,�B/gqG&�G �P�>yq�<y�T�&J6����Q�ݸ���zG�.c��T��/z�l?���iœn-?V�%�	������_ΛW���&�O����ԗI!XY��wVq1�w���F M��0e\v4����pW݌�<�b�d�
ń\�^A1�f}�*�%��{U&�����g�T,̜0�R�߾��~�Y�ץT*K���D@��><�o��5�P.����a�Ӷ-�����Wm�1�A�9�xY[����H-c�*�ixs�� ����3mz��*�$p��J��-/3�>uL�i�YO�M3),���L��Հ��b��tF*�t{�$�?1J�>�=�1h�D�3�º/��1+г�ܘ{�:�B���Y�4\uۙv�'�A^��OV�Z|US�B�Z����1V#�vm���Q�۳:n:k�����t�+!^��嘇~c�;�Nd�5l����⁻E~@E(�Y�:�����Ћ[_P�6J%�_k�b��\'3g�����׽l�q����b���ޒ!ѓ"������z�2ޜ!�O�v%�#��Jf����� �a�c�a?D����F�ۛ�dD?�<iG�/�d�Ê-/�4l�(��9y�a���&����ri���Ew���W�ù{J��'T}�#a鶃vn��p�*cДm[�I�o�&�V����O�}�6aEԛ0)�#��o���q?�~�=�ڠL�ҫO씛�r��E]Gߒ�k��`�;ྦg�J�m}~��.������WW�r���xq.Хa6�v̻�BQ�}=�X}�%���6�s6\QնŹ��h�*A;��o��3�q�������i�a�J�7���`�l&��J?M��ȿO��VQ�R���H�CX���9��'�b*E�)w`Și|}e��W�u���?��f+}!{E��1�j_�!�?Gbtf��f,��M�)c��3Ӟ�,5��kZD�\%<ǂYYi/�Wp7NFv��~��9d�5W�]ji��G�1T�I^�B�|����Z������J� ����0���Y�z�T�=*>^��́������W�?^֢���ص�$���@�M�u֒w��]���.�33�|~p�M�H�0�f@�hJ�ʿbi̟/� <֐c�������q����&/�A��Ş*���H�Gr���[9`���H�Z{��C�q�ݻ1�F�v����z��O�Y!�Lq%}��������N'�������&��f��>�-4m�_�5��ԣ�t�g|�����9g��i��[���"4^�z^��x���@1����JG���G��c0�w�u�B��@62�f��+�q���/����ňu�p;B�GAiX ���MN���4$�� �jo��j���ʃU?���BL�7d�?�I��ʭ�cl��d>XB1�Է/�N�l)[���M��dx��zm���3,Ɵ�Y�+�>kR��[8CO�H(yf������5t[~$��G,�s���%��i������f�Uo/��_����k��A��!�E��{���sb{��ه�.`���{�*�)]��%.��� *4�C��Y�iOd��"8]��W�����%�gP�l ��� ��1=�p6.�G�������8�>#�PP� �qRVWb�."���VN)/�i��c��)����	Sw��R���wߠ55�1��ܓ(D^J_��{Z��V�Ҫ�-�?��\!H ��5SS��Jj]��4|z"�9�t�?�y�c��o�Ѧ��>�Q�@^���O�b��T���
��a��s�?�y��lۋ)~i�ns�㫘-�ޞ��v�[0���{5�}��)��,r�rz����/� Vr���ы<U}9�;�j�پ�_�s�ѥޥ$�1����_ȗmUl�UKY�;��(n���w�rs<UD�Kk��,N��4�� �z��n+�`gf`�G�noh�|�6��َA�"�\��5���f;,��Ě��a�^�:wn*:��	Б� $+D�p�Kѻ���]�ǌyb:�~�f h"*����f�Դ\�I��B��]�U��dq�v Dd��� ��I�܁C�	S��M�2�*�?�ya9��ː����������Ґ���ΠG��˄�H��oO�z9Hb�NF��.���9}Y(K�5�n-�f}m�?t���{�[�^�Zq(6�����"�*]��_��2�������6?�͆W��o�e��q�����Dz<��yo��$W��������:>��G�+	���Wf�i2Ww��0loZ�oL�bC1�όFj�l1R���T2/����)�uL��y��N~A�"��$*ř�NZ��ۤ&k�`�&ϰ�h��ʷSY�$��w&�o�侽;N�����Yt�u����R��ڿ�l5�Z�Op6��������-Y0�-�Y,=�����X�f����ˀ.[ڴ�4(��s�sk�e�*��GBZ6Z����~"���/M����M�WVY\��l���R�k�)��Y�p�+��j-q����U��l9L�T,��^u����1j�?:V�+�q�@<ipS12�8����,��k'L�:�c�1���+=�O M\���rM��A$|���t5C��I1�d������+(w(EX������]��ܚ�����O�y�'0��nm����i�]�KG\�LE��1��L���L�>aDz��I%�r�@�d�b0Ҍo�º��B��i*���Z��l�>u�D�F6�U)Y�����1�mB��نV�3�<6����"���+�c"_�/��3����s#��)h�U����j�
δ��������~-��V2�ޖ|��y���.Hd��R��a1@ce]Z�b��l�5���8EX��O�1���	��֢O�`��ŕZ�T�z������Dl����@?�R�Ү��.u��#=�G�qP�@bX�c��`�S>��ԧGp�H@��������O�,��z�X��d<��M���<�ӰC9#c@��ԓwi.^�LJ;��r�F�2ȴ�i��ܦ�A��J�b�Y�t�r��g��������X�B$J%լ�f����7��Jg��QV�j"3ŉ���GD�r���!�Y9��ql]��{3Ժ^�+���id��V��`��x�+O���.գWj��E$8��oO�ı�;��7S"c�4/�����^H}��h$
�Ӛ�����#����9�������9:���/��{m�B{������Ɣ2U�Vq5�q�����d%+��>����������aTo��E#���#��c�a��ވ��I�EB��� ��^*��i{'6=�k}��$�3��t�5�A�y��lT>�*��fm�a��/�!�����F��Kf�b�!)�"�Ŗ��ȼ �
PㄬC���%�G�x5�����fR$�����ߤ6fqm��g���P��D'^��;��P�C�*�)ȟ��T�����֜��>��V�4\thΘ���U65+8���q�GI�jv��$�@�9l�����%��m�ي@
�U�Rg�qxf8ص���ؑ���oSUn�B���?~�����K��/d�e�|'g�4�?&�f��W��Y���:��fNWs� D�P��d�>�D�3�������E��v�e��۲Gζv��e��)_�
f$dt�h�o����k�W7����1�2�)f��ɗ���h�\�N欀�8Zx'������*@����1�9d����pS�� ���3 P��G�Nb��*惺�T��v&��PVV!op�&��[����� v-�|�t݌ ��ʹ�g
�O0J�]�٦�&��T�Zћ���g�+��D��0�8�h��:
��{Gi(k��}��� �x#�b+�&c�M�ϵA�����p��>����Kp�΍�ަ���q��*�Eҿ�H�ŀ��z��x�\�<��P�g@	
���Z'����\����Ҫs�*TM���.}|ޞ�����,g�f}�gi�����$TT�죊Tj�~`�z%�Η��<褩��pd��F���{������.M
�򿾼��h~<�ܹ�@ǉ�ͥ�^�-�T�� �\�Gq<��B�&j�F<ġNO<z���0{z���8����8�P��Vϑ��[=���a>��u�K�0J�&�A]����XL����ɽi>Je�d=����lο!���*a�?h�ye�����rt�7���ܮ�A����;Ʒ���t�Y��A^y=�b��3'%����x�|�2�T]"�2��p�ҡh'�}�A;��կ/�Dnnt���P<9�Z����b�����|�$fX`S�vXOB�J��S�n�v��'& �3OSߐ��0��;Q�ؑ=;ƥ_����ً6�������/0l���q�߭��L �ݰ��G��J0{y�d��0���%���y��<	ҟ���S!Cȣ(�ykYz�ȢU6�*�	i���:�C���h��:X~��r�o���`.i���_�z�Yai���ݏy��H�ʚ����4��4ve��m��O�b���˝�/]�^L(G���o�趸[���ף��-k��r��Z�M3C]��D��Ǯ��V��K���y��:��t_�{m�&�K-yk&v��S�����p�`���uŦq�D�D��3Ґ��SFe�XܩF�Y0Nh�<� =Sg��}�oe��ܠP
�8�kK�!`��E(J�?��dz�C��XL��B9�����g�2%["6�����x)�j�����$��\���� ~����˸�t*1ȵ#����x�0�w|K���m�E
#+��`��nf�3��l��"�$֟����y^5�/���ݔdr'�56c2^��{�ِ�g(��U��=Neb���u'�k�#�����G�KH �I�is(mr��+����~>�܈'� �y������@�I�n1�C��z���[jqR�vgHt���NS:��h��.jcbq�������e����-�a*?��� \D��Vt����!��u5�`�û�T��V�A�ݬ������ԉ�g�������,�2���U)ǴC�w�B�*�b��{��,>�`W�������FY��:�UB�\."$L��}���F_��־�P���[!*�/��D��M���#���r������ش�j��8;�	o��=�Eo�:�n�Z"��֠�f�]՞�7����ÖN�NeY��X�	�Vh0ln��g:[H��0�6ó�2��j� ����x�nE�#��z�}�QV�*X�Z6����*`M�'O+̃�ik}N����%hK�|�sk^�����(�>���e�	�x����x�y�!�P�yP�P�̎�c��|$������w)�c]2�����\!`�^��)��K3L�?Ļ\|%Ld2�,���
-�}�I����6�k��9q�(��Η6=}b
��O�VuJ�M�(e�(���.Pp��3�=m���O��i�<��k+�	*X;���U�^�e!+%�{7��,6+�:^�Mi��������4wZ�J'pr;��H0[�2��lF;1�A�{��k&ү�G��1&Jb��i�_�\�x�I�1
�^g%5u+� i�f�h4��NQ�p���Px]R�/����0��I�"�I�$��RQf��R�}=-���ز%V��pSy��U?�MN�IԈ����|����w��ɯS�B֬����ڍ��?�I��o�j�3��ɟWjB���UW��=ͭ;'�'���Y��y���t��n\�����]�����w�g�}�\^�J\����z��Q�PY/|�̥4E��{|%Z�H@	��`�P7Wu�F��)�Ӡ��"�R>��@A�=ߜ:T��T\b���dJ�<�|��a�,�Lk�܈�Ows)�p�(]�h���ʮ���ˑ��;G�K�`z�|+yboA����@-=�Q�M�Hk2`|�<}�2����f��E~#�g����O�b�)*4��'5x�dQ��C���
b�0ZI�\�RM�����bZ�S�����E| HsS!D��Q�j�-������$	�A�g�w�?�{C���mZ�o₇��}�t���`<�:�4���6p��nb�A�KסQDR���#�����M� ���fIW#H�a�݊u�2�e\��usv�����%��� ���)��J��P�bܓ��u�C�n��?�фd�O�|���n��P[)[5�=k��gƮ=�urE�:CS���K1��x�T7�e�0��,���q��}�v1���x.�~'�qf�0�FZ� p����1���L�)B��q���Y��վ��u����;�X��ZF#�ܨs$�L!t;�CZ��Wg�,pQ�\?�}��aQ^O��� �u'��0���W�1=���\��Z�KܚG'l����;��KG�y�ϑ�j� �,�:y����J��3�*1���z�	\2��
V�o�U��?�qc���t�ۯ%~���(��=��0xӤY�"FK�P|x���Y2�KIf�q}xc���&:k���֙�3� �
�Jmą��a-�C�]xY0�Im�:=Hļ���'��M��7J�nTCL����kf}�k���P��C�OR�ěn���J?B��zʼ`刨��됷]D\������R��0�}�Ğ��o��v��p��U�uy��J���(�>=�dC�p�69�-���b��T�#�#�	;F/�!�
�����ߩ|�֟r����e����/��]�H���Ύף]���ZuZ�������t"x���쯚�%�	����`�#��d\']��~Ny{��8t&�z���nؔ�i.�N@��&��iP*��vY��{<�ӆ�xq�ς(���B��@�N����Z�d����^D�h�c��j�a�r=A:6��h@oV]k{W�W�
v꼅+6ScW��w�oR�?�	�w$%��H�w�Ws��'�9�ü����t�M~�D�-1U3B�;Vd��0�����֞�l3��330�_x(�;��dq:�&ݕ/�}|9��q�WY}��2:�9�[8}�~�Gq�U6o������>��q�%�@.��ۙ�$�i�z�9Wπ�{�ص�'�����bV��,����῾m%�(`^��`����E�Ҫ���хE�Q	�CR7�x*[��
�F9�=�������(�v.7��0{���6y�%���<ǰ�3F�K�X���ޗ����i�����?2.����H1�Ndp��e���R9��`��gq�:�\��z\g1��8=��
Ah�7+�P,U;�E��/��C|�J$C��V� ^�`8�m8-út��jf�$�+���-7�@f��r��G��EyIǪ⫅[)&��Odç�
�)�uen�d���~���)�հ��G�l+�?�}즘��W��x�$�&'�}��<���1��d.�{����^�ڌ�X�&Ȋ�[�4f�H�#���b�Gׅ���6|��F#�<�{�!6��H�B�9����C-]�eӊR�g���Wk��)��,��儋uW0i$�;�HgêPW��PĹD�!�$�4ː!��S3kq�����+�Z�S�������?��4�rn� 3�ʔZs�^>Q��HU�bc>#��L~82,E�Muq�6�k�`2Κf�o����:�e��e
��%��bh�Z.����q��l<?4��LW@�kдߒK'�k7c�m�$�9�bv�� U�8� ����2iA��i6Ѐ�����R�O�`0~�w�L�tj=ΪT�Y/
i�
���Z=+�6H�����G���m�m���M��\P�h�%A�iz���",�td_5�y��6�r����Sl�����U�n�7���_>̞w�i�6t�F�(�K]]�mIǀ�����mx��#�x����N�V��?�LLf1�J��`���¤�s[�c�=�0��)7�|r�n%�@֗�h[|��!lLz�M(�2�'��R����t���e���� 	,�JI���h�:rcT7�y����l*N�.�V�;�������ZU:uO�:\9���������%���ƃ�l��cǱ*7.��`D!�܀ɝ�����A��yFSG�(��'r ��I���;U�;��~��l���`=!���5�_s{� GP}�qn�)6��o�e(\��*2&�����3� �j{�ϣ2��)�o�����ŮwF��"�w�'B|�*�=J���ty@]�]Rb�ǧ$A7�2w޳'b���׮�x
�2��7��*�#�������Bk�#��G���]� �_W����G� T��Z?�ֱ�j�J(ю3>P�����y)9�fbξČ��R�k�n���lS�Ou���;/%���r-Yr�`R_�n�'q@f��?�*'*W��1��\�vTB�X8(��N�����S�V
���j�2��|@��ҚIM���P.u