��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjfm~���*���`Jk8�ݓ��
Ƽ�%I�A~\����I��3\s*�O��k9oi�=�ے(F��Nq/��㽠q���X�E˨{�bi{㏔�㰧a��m��}�����E�+����8��\���-2���L��ût���<��*Q6Ҋ~vl-� a��e��Io�"�$|�.1;B����;>�g��4�&��:t7�"zE��X���F�ft�PSq��^�F�X�d��6<�o+@��i���h����Џ�d��4\7���0G׼Ұ�mblO��hW�����G�๻�~?	�FP
	l�3+�JVH�n�6��:Ue<P�� �~$F��u2_'6�g�сQ9�2����Hb�bg�.��>`��s���U�w�����Ɩ\�ԁ�3������U &繫���R)�R�ʌ�Vc���k���i,�1o��C�����.��x14�����]�8�]b{q�� q��!�y��/flZ;����<��2s%��Z�)$�3�����=�MΊB|���m�GA��'Ȇ������]/_������zX�p�³�6�h5kI����ў]g?�,޻��y�s����WJ��B���P(^Nk#AE�!e����i�>��D����&W��n�Jޝ���������ɨ���ޓ��l�<�X��g��v2*��'��u��u$�b`re��y���o��3�SO�NGN�L��@+(�ݰ�W傪/ ����4�*i[Dp�0��4�Lm��7uf��𽷤�IQA��$@)��9��zf���HL5��&�����!$�������mvuшec��'�q��.���ڶ���y�Y���bu��%�<������]B:>���A��=��`�T�z�<b�0���>k��8;�^�u7�WQ*8�#�*��4;$��`=f��� F�kK���0.�Qߥ���h28�������H��."ݮНh)s�,�$�x��W�7����9��Qe�>4p7��z^M���y:��r�ᖝZ�����&��zCӑ���5:�p�;�U��2���_-�pj��@�N��nQޫy�{q��!���4��jm �_��!frϺ1Y���Ab�E�vE~�(�Ru�L�Oca/�,�������Q�����H�U��]�Ѥ����q�b.��?�|N�+�(������cf���I���=�A��D nSuS���0[:��ܟ������:�UH�xA��R�n5�+�=��j�S�ܝ/���h�	U�Q��-")��bU\�rF����-&#��y=�ox���i�C 0aY�x&��=����� ��:l�^�܅E�8�5}��P�p��Ry/�*�/. �FeG����k�]�Zk��X��Q��B^�|e& ��*OZV̣q�~F�v�㰻[�vUa��d-��ٝB���"�sY��M���CC�}�fP�'A��0�:�<6!��N��Y������Y��sT�2�>E�S*■��Q�;4K}��6&{���m�9E�ڙ�@���c�`�L���ܴh:��[��`���>A�5
+a���;8�Yu���Ğ�eQ��"D/kj`��!�QT0�g[p��xO`n'W�����*�%���z�"K�0
k���x绚�`)<7�
�)�8a1Hk�Ǵ�n �|T��q��Vrt}�j�[�n�z[}f��I�K�й�]�z�`�y�sV%ف���v�o��#W�?ΰ�8 ��-.L}�8Q���^hC�Ы���� ü�����E� i�p�ϯ�ζ��{�.�M��ʮN��L��#�d#�j�ł/�|�AK�g�i��{��A�" R��a]	Fc����Mr�La�2\}	��*?'�G��`Q{�tJ>D�
��}��_��9-�;>4����6�d�̾��A�	{�~�gfi,'C�O#��励��c�)w0&"-41�������jN��){�w�P�(X⭌�9��k�	>�0R���,_�{+���݊��W�f�9�>��� ����y��ǫg14�-���P�[���y��Cr0��K�^�&����+��)��~�Z�2��?Y����cUծ�|n'��"0�����|����L��a�pљ�}m��n���T���'���p��|����q�f]��xꬭ���qo#���c#�(ZJ�Ln�e���eh����b�ǚ�?"��s���de�Fm�����yT��4��´h�/�W�9%�A�.,�y��>�^����;�:N}ϭ�`t����chz�ţ͎Xu����yf"'ci�V�W��(��{J�v��ǧ��x���?�$��^�����}Ƚ��/U�K�⸋?+,�g�hW'ٜ�:�0��5L[T��a?iK{� ��ىu��N�����l	;zu���p�N4����='�����<�"�;Q����h����SM�!�i��&�c���b�w���C���k@���`���v1RH[���zoh:pN���xC���p�D/�� �F	�<�;v�3����kv*1��!F���)��e;�5;�X�N��Y����򔚥�m5��4�@]�b�,�v��Qn��yh_@��%Z��B(E��;���\�K5]����͏��6z5��m��| ����ذ��/�B4D��������.�n�!�<����D���r?�.]��&�L�����������>�����Td�kS&�=���%��r���<�e�{�=��Y?N�r�l���Z���.�?�8�G�b���)�
�����Q�%z%}�h�.� _c���L�����9r��FY<��]��H5j�DI��c:�-2�0'��PA���h�z9�L!�U��<�w-	�b�!F�T�)ן��bL�)�ʶ�E��]�ʏ%�(���s	��q����>Ly�S8f��H6�e���a�
_��.Sk}l���ҽO��,tg5$�󻜞�����fJQ��LH��_F��G�?�ߋ�Χ���
�cS�u���2#Į����dNʵN�dq�1Z��V%3�g��}Կhո��@ h�h!q�e>z�D9<�h��21�L�S%X��}��
�R�z-�}QX��7 ��P��ϺB����vO����㛮�0\E�/N���e�	S\+�8g�e\#�vo�8@�Nx��� �2l��_>�R��e^������#��b�D�b������y�L;*ZS֎��\��*�.����,<C�Ņ�������h`o�I���j��:�|Ks""��%�G����V0YL� ��#�s�L
��i��W�k<�T&����HPA%�$��B����K'}"Tf
p"�$���g�W�5,��o�(	���te]����z`ہZe��9�+NJ[ߨ����|c��X�AT>�m�9�@�0�������&LqLm �$v�;�E��'��5�/D���tq	��U�D��6>��/^IA����X]���>�l'=�!�	�]���dD)B��^�Jw=��S�EY4P�S�&d`uQх���94z�!ƺn��0�ǿK@�T�=����mnw~�V�؟�p�l��$~@���`/�	�Q�t!�Xu9U��!m�����l�IE��<����9��؂��)jV-���k�
�>r'��(��5��
�wŢnP`k�L��H�JޕI�v�,V*�L��KB9M��RW��u��r�3>1ac#2�b���������Y��k3��5*ʫ�	���87�ڕ�٘����k�D��`djv�ZV׻;��S�E"ߴq/�G�2~��4�Z�?�Jg���.����z�S��l����;'h��Ϯŀ� ��ܻԾ���`�����L��I���H����DGB���/�}��V^dǔ&lW�NUH�c�c;�N�ew���_��=D 8��k�*ݸ>�7�8��td$����ؙ�V�
�_�D��Ղ�E�6G��x{�q�Z@_L����B�)�z4X�L�= c-��G/p��������q��:�k
�-� k��v�hض�GQ�H̠@�iIK)�d��l>��t'��֘���u�f���)u:�(�Ͱ�n��f���"��RgF�)��1��D�4�B=E��Ƞt����GQ :u��2L���k9��	`��pE����fd���lfii,/��`��������j���u�&=W�4N2DP PR0�����w1��9I.�V��G����,�;8�.t���ռ��G�*�6PtSsF�*��ϡET�D!`ӈ����%�>j�A\j�I�"�LFC4'f�3��5�̞�G�!�)��� ��S�Ek�:�@��퀭 d�z��UG�͏m������v/�$
M��\(nT^X�Q�����m��O�[}D�\��>� U��gB;,3nj���[M0i$j:�p�cuX�C����i lJ߷G�V��73K����ƫ�
Zf��S��7z���3n?dI��ڞam�Q/0�9W\+q8���98@�!��.YS{T+Z:�:�����9��Nk�����׺��YQ��� s��}��S/-�������8༺N[M���Z�d�T�.x��R�m����q�<������t���6C��6���.e��=�h'4l�+'�(�9��!P����2�� n��$�a\E��⒔�M�uPO��-W[b�%BϟHuL����eUC���q#hm����t;IP��I&L≀�	�;>�R�)����$U�������{����;^���[��e]ߠo�<c��fI����R~q&��"ŦD"��Y�-u�Jc2$�������	��������G�xRx�'����z&���c��W,�TU%3?% �No��Q�@��U�.��0���8��%:/&[�×ř���c�R���i+�����"ld�ϴ5��� ��O���0o�q��;���1�`Gۼh�ez:������嶨�&�i��f���9K]ܨ�ψg5���6�b�D��6���˅��IԲ����0������?��7��&��> s�|������G�e���G�)n'�K���g4m�dL�d;��ن��sUz4�?7�H!/n��.;�z�4c_���\��#Lq���n9X�U�Y%^�չ͚^��fA<�'+��.%�pv���[�i�K���|{J�N��1�J9`�����^_|�P$��%�H{j����J�r�5��w6;lP��$�*i�%�A��"_>��y�6E�a�{9#ԧTP�ѯ��c���Zu�`m��N�P�	�S@[R��ˣ�\�@���l��B7�����2X���\�kU�]!z��$N}/7��񵸺��W�.���F<�������g�~C�ptdC���s����6�Ō�����C�`&Af�o�G����``n�Hy��a����߱��P壙���q���Q8O�5�Q􁑐=F�xB�̸�����vQ)n`�H�ɖA���:�����o���kd]'����|g}�����ܕ�y�-rY]���%���+��|���Wn�duV�z�;�G���ҭ�7��-Efp8����U����`���p�G���R�|���,ZUt�j��t>�^�ȴ)�V���O��z�(�{L0�Œd� ������Q�>�a���W*�����ۋҎ��+*��~&�o��{#��U|r}1�ϼ��4�p��o[��l��k��{H,����ǧ�: �~�sc,Z�<��a�����8�ﮒ����l	dϴ�n &�݀���<A�(����~`G������"b\���Ҟ�rAY���ͳ���fez��^s�?p�{���U�����l���Ϟ��o=���^��Ii�^��.���7����$6��	����¿GL���ToJfG��c,B�z�!!��7G�<�w��T03��ȱ�2�Z�W��N���vv����r��ڠ��̵,��ѽ��E�����you_GwD�<˦�J�7,�a� t�úøpAd�ƹh�?3�Q��	 ;�8N�B/Z��+Z��)9�*?��b��j��7'�jB�>�Z�Bo�y�=}~�>�#fD���~L�!��W��堥�C<bs��%|t���S�í���Cu��I9����$�ss S�J��1��(���,�Vt�Z^�YOTyO}��Ÿ�|�Q�ߦ��J'��}������zl�������ׂ������0��vbDg�>�؛Ӗ�1=A�vv����.I�>�(���_�D��7^�� Z��;O���
�(D�� ��i��v���I�ci�s�O]*h��uD8�|���U�� [( Z>#8������l���0(�u�K ��� �f���^^�n�Q�f�����Y7�5��ݳ�'��u�d`�e-Ρd_���zͤ&4�mLn�7��9&c�� n���R/��z`�:A�"����y�7��\�|�b�l\dMψu�c��A-z��}Ţ1,+���˳Ȁz��0��`�#�@�yK�_�]�>_l \\�`�yo�[�X���!C�@�Q����v�2ײ6��2�F|�AKx=,B���X>`.I����k�d���U�,SB���Ti`�p���6}{C]�K��@Ly\��d�uK,_��]���De�Ng��\����ʧ^ {s�}�|��|;��)(��"���>��P�[aq"�*��sj �2Im�F�B��`�\�ĉ���#����9N)��8��߱�盫.�:o�{d��_}�׋k��P��އurx��z܄��d;B=����,*�QxG��_uo�hR�!XY�:X2�l'����Z�X���یa��]xy<��틐���Q�*�K�W��K(nR��(�÷!�^�e4��R<��������G*��7̚h�����m�~���2U{+Cԡ"�tψ-���^���1)̋o)H��7ʡ"���>��n0'��q\�S��ZdutK�!L���OUjo/G�p�ܛ��>15v�Z)���'TG�a�mq Ĳ�t��Jr��4{4�ΆM)�lċۊ�w�pe����r��֌�͆f�ޠ�������/j���B�Ӎ����LY7��Ku�	�Y��ב0������5~]���ؿ�s�^nv�L�.��i��G!oR���LLR���7�W�A�)#�~i4!y�Li�,z���qScgg!ۜ2�����)�tF&��8��[�H���=rU����vW��ф<d�~
H�@�[m�� q�??�0$\��� Q�˷�ǅ�81	��+�Q8�ב땤k�jj�z���@L�X௭����c��B���$��)ű�Jg�~��پu���m��zDtz�F\�H/���`����D��1�4�~��<�EZ��느�[����ͯL���/N㯨�/�Y�a"ZlO~��
;���ۿ�r#?�k���'�CA��R:��]p0woۯv7#ވb}�C�"��@�Ĩ'�6w	ۚZ��(e�H"����I�1����]�b򛀇��o����W�V7�������	�T3ZX��XC���]�Q��ZЁw88o`�I�}���H��[���lxh���ZS5`%=�X�����íGz�+R��מ'P����C]�Ԭn�dH�C⮷{�$���V�4%�����	(��W(�rg��\D2�bW,�LT#�P�[}lY&�ߨ9s���{��ݪZ���S(���R,e�+p��Bx�@��b�L�j�.�ˑ�e�49㞚By�RK��CH/���Ͽy�z�/��2� *H�����D8���k�?�f>���9�G��iukk(�P@�\��6�ݔq�<�ѱ��+IU���pJ��rPL� 	ʃ�����a���n��7:�� d��#Q>C}d��@��O$KjO���ξy�ΆkH��'l�!P�N_�W��/8NV���G@]�3f.��9|�$ά$/�
:�W^R��9��cN����/��$���Ԯ�)�+7�bR⊖dFt{��r��(F�3W�C4�7�E�I6UܸӠ����d7�#V>�{aeo���pW<��Jhh�¼*7%F8^�6֑���z!7a�<�8�A��[�0�?υ�d1�ӫ��x⑫���]����9ԷB͇�o}k0S!�M��hw��
^I�F?S�}^�2�k
���O6	����gL��B�q��i^45���q����QJ���"�a�Q���g9m����2䬿�����X{�.�3!�d�?��'����SP��!��HpY2�	ɺN�X����E�k6���t�"<y�=!&2�=�N�B,�jg�V'Z��h=4Ȩ�PGL��⵮������|x"���~�>7`�>^�[���1�_�>�S����7>k�˼&�nN܏���z�W��,K�SS	��fwY��󯎈݇��%Ո�!*N�΃�!����1�c'��^���{@�Ow��6i�4�(7����/F���؞2�e*U�"��ezU�]����Q�����۽ ����8�<qT�T����U|x�K��}�ǛSA�)��g��{��,��C�1��!�YI�8b. d��W��I:��L���\+�A=+*}��k��i!��# �ޞ�_oL�;�ljq�}�6�>�'"_��Jzg�f�mx-�|�R���t����x����a�1��+��iv�B��Aā�ʐ��B�)"�K�;b^Q]�x;R�j��6%��&7����l�8%�Cp�۳0�+W�#6��
��fxF��Q;!�%�����f���y�[�/P����6�.�C��hOr���y26Q��d)�K��l�+���vQ��_�`t�e@j�H��E��О�ϴ�5�b��4]�eǮ@ G� O�n��8���|��a�E�\�W���܎Ğ��xwh�>���O/>{����-��SV���	�;j�GG��2 �-A����I�	x�����9-���1�:䵊��,��Ȏ�;@��_�Rl�R�]�e�������0Fƽ����.[3VP&�2�:�����"�C�d�f���PnBY�\/�Z�s��(�K�a�#��{HC58|��4� y&�k�<�8F�AY���]py�\�����J�C�D���ff@��Mxh�^d 2��O��Ű2�!f��3������?.��FL��y��xx(g��AB�ӷM�8��C��E��Y:Q�N,�~ H�}.!����*m{��	�pe2T�j�Y0<F��&`�d˖c�O��jۏF��+�t��p��9U�8yd�xfb�n��푠���0��y��z؅oC\�i@��4Dۃ��o!%lN.�����9 �s���do�=�!8b�[*�����xr�Jx�
cĔ��#�Ҩ[=?�ñ@C�R�a�B�f$m ��A��]z�t;��M�v��b&$L��|^�ZZ-�~��3*�1��p��Q���s궐�bq�Dq*���mf{�4��|���;�f����G�?��[�S���kp� !��8M�/����	&���lZ�j�ޙ!����a�l��=q��VU��w�,ά���YE�lS/N�����&4�2f�ty68�ʁ��}�0%'���-��������a
�l��Q�eO��H_�U�X�?�n�>֙���eSS�z��m0�.��Fxu�RK�i�rnA��8\�0���sξS� H8Y&4n������aKT�����i��`Ӗg�Kԃ��QY*�Ao��^5F�va߂�e� T�ȷy�Y<`$"�XD����7�*��s�#�MNK�u|E3U���2�t��-G.v7�q|�9Lﲭ��K�Y��P���
!�B��˹sl�i
9;���S�(�8b[®�h�����xDTW."�.|���a��wݑ%B�U�hY]��x�������d�;9V�S� ?���	���6����~i��u	|d���e����D���u���-yub��=�ԧ�C��;�v�Vz��	��ҸԞ/��n���oe�lrۤ+���1�/<��tj������<���uk��
�����O��ߠ���e���T�(V-	
4��o}5.�}����T�k�0�j����d
:8քnT�^��?Q䔷o�+�̵�<˰\�,V"����F��L��B��l��-@����֝����HY��2L��\�D.�r���M���E�,��.b��s�,ߑ�m��kr��	��w����dv� ��r��>ϥX1�~��1�^��r��<;���i�������d2�s�����"=�^3s�Tr.�xĬ�2c�S��,��!*[���8��N��W<�L�3Az�,vr�%��C���I�2H�Q}-(��B��rW�K�cEĨ|�~[b[�郎T�$��kK��*�W�0{(�B��^9!�2dm���JLcc͗F!�%�[�lQW� LRE�HRN\�����.L'&N�ߩ�}��s����,�<�Ϥ�;ӵ��x$#B|!h�@��v(�F �[Z��:��F	�I���1�22҃�L�3[�[�H�FV�eJ��3u�Li`���-�)m�ww�f�S�?�0�A]�/�;n�*��'=���^2ꊋ�Җ��:��::�s]��/I���01�_�����38��\x4��[���^�*z޳�����O� ֨�̶p@�n�3-�.�o 45���������}��MxX�)0:V�L 7/���=��?��H�.�f[�p ��r7��c��;#��%!�Sv�gJm��ڎ]ZM�pK���HH<���_���X����	�^�F/�-��TCf=�GR�ryۓ��O������U^U��m�l�"[rqeS/X�K&�sR�N{{��h�����-��Vo�N�`�Iſ�8x{��xA_D~x[��]:�z ��9?O䅴=	�� 4�;��jn�u0M�n[^D!��5�e3.)AY��%���Κ���ܘ�FZ�P�c�龄�p�s��ֶ1w(���:ۏ�<�z�$�ȳńtQ韧8Cb��������ļ���Wm�Zx��Ϣ��s�!/���[
Ӻ~)X�J�j��ٿ��Ŗ_a�^�p1�g$�Ď�K�	Ü<G���sN-����Nn�"S ��Z�����aZ�����i"��C7�l,���@A��}����In�p/��J��C��Fb?�y��cj�8�K�)N4�Q�Ί���h�n޽���gE*V�i��ϊ��M~���j��DK<`��Y߅-�d�qFn_w��UY�d��>O_�R��FU��
�w*�cx��U"�
$�6����ewV.#��M����!hیvr�1J�]}tnW(%^��H
��
�!��c"f����u@W�H)��b��,�+��j��h��iXj�����Đ���d�5ȀOr�Z�gFj��V���0������1�N�N+��ș�	�
�o�E�{b���Q�A�����$�_�_��0?�~An+h����o��>���-�,��Ƨ�J�;�����\��:Q���G�OF�Q�$]�y��VY*�Ϙ��+]����̺�1
>�;=�@J�a���s7"Zj��Y`�&��H���X�|�	%f�@�=��������h��3l����n��G�kXZ���H}-�]u;����H�{�spgF7�N�&'�b�}��Ɠ��}b��\j�>�S*����8Sz�t�����4F��l%�6�vy��Ԑ~�������/�3ֶ�_*���Oj&����N	��q��Ǿ@(�d5�U��8��|Sp<V�x�66U2�{emjn�$jE4���<d_�0�x�M���Qdp��J��`,%�*O����h*�n^��� HG�(�p����Rl�B��o�/�K�l|�r����\7�LĎ_�7;f����_�WL�h�;�&l��R�ĜN��\M���#7�XL/x\���-�A�nQ��2�9>�Yn���BS��V�q,$� ��M8�*�E#wwZ[�GF[�I��l)��8�]t��b}����!J|���8�-EG!}D-�%xY��Q��"�aLDS�(�	����etl����IU�
P��
F@֕T3l���T̜Ƅ��������	����]În�t�y&�۠
��u�6}�}���>.�q)1��6���AIX�۠�s����o�C/l��p�Q�i�"��0Ya��|Џ���FL�M���f�Nά�	p��5�����A��s�G!i
�o:erwP
�lH|E�5�_��v�Ҵ�n��3y6m┧��0��qmz�pa�}<z�ZPG6=ڲ��Q��=��������;݀Y�V:�J��$���	.!�H��
hLGK��7D�S�CM�G�W?z��Q6 ǹ\Ro{�.��ٞx����6<V�ۂ�,O�_|�;Az4�O�a|C�,
ٹ��-`�>!��s�2^�/Q�����I�G
Ĺ����h�k25XM$���Q���v~����(���(K�<z�oS��;/a6��
�#@��S $L�X��t��On��YCm��޹�NQB��qB��~Z��TAW���D5����Ru�3ݒ���N���RO�1�!5�eڣ��
����/�S�_������>k��"s�^@i�Z��7E8j�PO_�Ҏ�4Т�X.�V/�RR�oC���{-��Kq4�&�N�E8�SU��9Q>�h;c��o�!^��"�LF	v�@i�?�3�,;�����6�~�ܦ��h ��j=2�F��q��GH���U.�߽{����:H��^ѻ��а�]����o[�>"����;�*x����~Ƒ3�^��vωW��P��*4cb��gS3�S��t�)�3����
w{��s��?E�|>CT q���X�נ�޵^.�.N�Ap��Xފr��9l�I�k�Ctf��a�&a&�U#:�"����;�
磸*WmZ(cM%�X<J���lt����1G�+K7z+���=ʰ�Pk� �����p�̛-���&�#�N"X��pRS��k7������n�M�#�. n[>2Z=`͝����t��v��+S��]B���H��	k(O���E~g�$��W���"[�&�۪ІΣ��X2*���&dV>A�bs�a.˟�A��ִ'��x����~٪���)�3�G�jRO�U'rrH��lԠ��MH�DQ�`-�pN�S%3rPcM��d�Wk	��%��!��@� }��_�����g\����'޾�L�_�:-t4�P�8��|�'��@D�&o	ں�k���eH�C%G�՟²|�̟W8y	�Ќ �5��gk+�0��~ 8�t�4S&�>�����e�.KSR--:�A�����Q���v�9vmv&�ʟ��*�n��Z���#̈́��ԕ܁�:��I|_�b[	����a�����wA�|�(%���`�e d��Mh�:ã�=�'ǢB�D�4�=7�UPu�it���{�.��	��T^o���Ŏ~����B�,���H��KM���X�9�GYL�_� ���8�_�aFbG ~���R��,o��/r94F�V.LG$��c����ӿ1��&��]��D�ND�-�K���\�j�.a Չ�gR������1ُU��V���*�w`�q�w�5<��B,#�zS���㎡����vQ�n��HQ���_��,U�������=	�����"����s�&�ɒ�˥ �c7�)�D-n�t�x�����{L�L�N���v�����)�8������ڀh�q�%W��O�m5l����3�dܦ��i*�i#N���ž�.��`�V�v�ÌROr�6���T/;�FŎ8����M�2|D�,��9�^���%��G�do�S��?r����ȭf+��H1���TU�κَb�X7�(!u�J�c����-��O��1��D9�%��%�ad���m�C��b{#�s�˃�G�x"����0(�c=Q_"�N-�����J�@��pթ۹_� �C��Y���}��z����_lF�~'�Kl����YeF�O�:%5�4��0e�Nmm6�h�V�1�!�r��2@/z���[0l�!z�FGc�mc�KPt�G���z�A�\�+�4�R0����ig6�4�~�#��on|F��]�႟}u�>��dpO%jZ�ُo���:@�TU~
$��$QDv���}���˸��;U��x��;����:����-�-�ڏ���a{B�g̻�>H�r�nJ��aY8�,^�l��̃R5��.�d�nl��kd�e+��pZֵ�/���Ck���	eIT�K��/�Y-{�G��L)�%(k>�mM��>뷎q87�f#��@R9��$>�99�Y�[oR�6��c�U���n
x~���VU�x�6ND��;_q���0~CG�G�N�=輕�A�j��sv�
���)��)Mv(�~���|����%)�fJ��q�7�8ޖ��Y����ye��9m(�j3�r�rH9������簱O=ෲ�]+8x���^��H�cr��8bӼZ�x����$���g.pX
ɹT�<�^KlEİ�^��6�抓���Ǩg������3������!MX��Ҧg80�嫿kc��j�6t������y4X:�?3�$Ft��J��c;��zL:@�t8��xT`�=�����QQ���.�֧z�El�r���%#M�O���Ob`$u�dqh�$�/�+�x���<�o�.�70�����$ȿ��m:�f��W��z�@&gbP���U�FS��W�z�y�jRx;_E�M������-c�{�_
0�kc���7�(!h�S�W���D�z���z�"-�ϟu�����+��SR�����K�"�Kx{��T���I�����wҹ������Uݺ�\B�ԂK�3p���R��WY,lG�:�Ӆ'�[�DF��j������5�m1b�:kԔ�z`+��_;I��¦���S���\��y֬n��O<�0�He���ó1�
9tV��*������	����Ύ]��v>)�������;��M��s�c�i���	8�m݅��a�۞�!rRf<�+#�FQ�l�u�6�䯬��6\����K�#�^��5���?� e���LKv"�Z���-Jq�D���C�3̕^d]P���G	����&iF>o�s�M�
"�{�þ�I<ךN�aڶ�-�
��YgK���gm��h#)���9��K��~!u�O󼀆�م(�'^q��I'AyeX4U�gS�>��E�pA���mZ�W(�f]m1�j����sG�X��|ɲ�(ˬT��3����XE����T�V�]jm�/`x\|Ј*���8·��em�,~�؃�&?� ����Q��~���9��4ϸJ�CN�)��y#���J����Kh ���"S�%�'Ցd��͸��"�5a�'��/+�꽜.ƛh���E����?�W �u�6|�l�E��N�7��)n]X��RP��[�8�:�jR�P]Y5/x�a_d9���'T��m�y�Q����.}�΋�0�����EW7���3�~f a�i	�M��A��w��������^K ��o��3�Fp�A�Ru�2�>���gI/���m����d���^�O��<WB,����.�u�Ƒ��ôI������b4j�7�l��"�1�hO�nŬAG��P���$7�Uj;�X�Y78��JpHr5ݲ�`��9R��
���=��;#�� Z�{ص��NS��BfX���ȷ��a�~��!�3�O㵻���$�R�!.�����n�=6�}�����d���6٩PS^(x�s����Z(	9�t�d) \�A?�`���6��O�@{��k˞>�ʋ�B[��j�k�k赆�5�K�:���
L�P�Q�ά�kҧ7#� ���֙㱃�&�B��e2j}\!������W~M�XY��nb�i�#��i�0�n����S�=�ߏD{o�"�"�LX+�^���՛�s�&�SP6f(nĎ-�m�e-�kM�hJ((�~�`Q�q u!uۘ�&!��c����i���F#_�q�x�9aA����x�r� %�0y�ޖ*�SݿeN�:�j
X��f �K�����p'\Q�w���:�[g�W���t�Ud1��<zK&�B��{l��y�Z���	�@������?.R�8��.fUv#)[5ի�ـpey��jj���S��_��9����U燋�7!��p4����Rߞ.���͙#ؾ.��d��V�)HE��Jzϯ^e��A��(#/q�#Qg���@�6�a���5�}����TB�Ǡh\,c���J��I���J�)G���Yֽ;A�̩33�w�b��)�(C��5�Zn&����St��xZu_ؾLP>�}�_��{�?�k͌�p�11N4��M�u��X*�U�-���;˒��Yr�q_Cԑƃ@2xLLD�,,�j;��1.�i�5���h��^gb������%��L�w�dH�B���^�}R����?�_���`,ik�pߤ��] ��Ale�����>�����8�;\R��o.�o�A�6)�c 80��A��J;���Q�7�����8,-��*c@"��cQ)�Ǳ�?O��/�y8����r��]�pkT��Z*>�1ߗ�Yc��
�TѰ?��*�aW��%v�A�1�����0���S��9��ty��&T�%�<4S� q"p�KH�]U�Cπ%��w��?�$�y�Frڕ����(h7�k`ő��)��0�\6p���[�E�i�`��D$@���B����h��2���ם<�k�h�A=��	0q����_D
�2��:��ʅ���^����g[\�b�:a[)�D��ߐ �S�����_���jd�y
���V�V��=r6��3�Dz2J�K���F�Ou���<�R��w <ލ�����{�c�L�q[[CF����j<���DY��x��K���eFr��E�$�V��)�5I�k���q�m����:�H�������hV�=��)ϟ�	��uc�[�T0�'�'/���F+X��
�f�K'�8q�����4�72#�۹��]^����f�OBv�~�Շl��N� .�Gh-wK���t���(�w�*�iP/!)��w���hjQ�1ި�Ĵ�@Y4W�ۆU�-ݤ�:�����Ǒ�f���qNF�v�E����F��^C&�I��Y�h���8��P��&��@4��aj }��a�l�\�����4��'M��Q!���7@7 ~��yX;�qP��}����-0}�39��e���3�DG� ��j�Őa:�dP��@j(�-�Z�5/9b�����?���O��fLnII7�v��c�t�̜���f�Z�7�Lm9���܅�(�+wXWl��hRh\�M��uz��V���]�ho��+�[7�*��K���m2�d�Z5V�Sվ=W���9y��w��lw�(�3��G�s�����WsG�4�	A���D� O�h��\�Y/�Q�<��q��^�����ە&<����1����� w��K�U�ݦ�YR2v�4�~����e�A����n8
~a��j^�y��K��b�\ˣ�6s�fu�l�еXc����&�ɧ�4��7?��q3�j<v8dj��8�n/�l��ҿBT~Xh@Q
v��:�9��(v�	��^�˛���Vݠ��
XN��|�	���<�tk��*MڿH��y���J��\���J����X��Sa��~^z#T���9d=�h�ZW����o��v�D��=b&�Ո���{����l����x[OoAzķ>�юᅀ�tX����E����-�HRT���^4\�*z	3RQ�1�Ngw���矃t<!o�����Ehr��O�~GKC��i�� �����uv=%
����^FfdV��l@:̸�ơ!���u�8�Q�P�]��x��0��z���D���gD�ڹ�7� mQG�����,���O� ЮR���-���#D��>�X+���R8�[sb�X�S���\�M� m�B�Rgޞ�eE���:�7T���3A��73U5�	��c���R�M��U�I�6��M*�4�����O���0c+�1~��!9�g�f'9����IRg+Y=xU/SX���.�������2C:Ȕc�"��FN��Г�%����Vy{:����$����GaЁ2�4���w����+��~���㠥]~fL8��x�/��ΫW������߹."� UP>�(H�X6jH�o��V����I�v���9����.Z\M�r,��.�	֒���6!��t˦r��9����Y�"<P�ᴅ���P48Q���dq�fb�<Lk�m�C�g��i�X�u��ZdU��ĵ�&�L�[!�,�0���.��u;.�C_�]0�;Z���S�Xp�#�c}�9�}hrlJ��>/���++m'���I�̘4����:��2GIs�h�-�7�l�r���;n)Ԟn���z`�+��mJ��-�qN�!Hy���1A��L��A���R
Or��ú���[n����� !�o�;p�Ui|:z��3�o�����HC
��<�q�����r�{4���DMۘ"����y>6a��z �P�;h~`-��lBhy2�ʘ۹`���Z���)��,퇲>��i�a�t�E"*%���4�J	�� ��i8ᆊjjȁ@�L]�n	���f}�w��˙z]�r��ށB~ �G��{E�=3���Ķ�)2�}8�aЃ!Ȉ�vǠ7���&J��?�ĔZ]\��� �g{���0!�idR���9������?E����s�q�MIU{ *#��=Z�x��D���SK�L��>��e��E#�h��:���8�#ܠ�$j�I�����"y8��;��ʗL(+ngO�EЮ��_��o�K�9J�?(x�#�e���"��q(��S6���,_����FO��I��
�}a�J,Y:A���qZ �a�"��z�rs�uvv!:�𡆑���#D�h��Z��u��������r7����3�KU�x;ȃZ�Գ�u�f@�	����
���L9�!���s0�3�N�ޠ��k�D�c���r��q1�ݞ�^ ��������M�3`�U*7)>�� ;r�C�)S;7 V�B5�!����@@����t!نj�w��?}��k�@W���B$)۳���(��0?����g�X�w)1�x~^̊
E�ES03(ho�m��\��ǣ����L�%�}�_�S�&�0!��!�>�*��*s����4���������#��"���ۢ�d`���稨_^��&������|c0�NԢ,�5�Y��Ix����eJ����.e��1ԤfnI�����B���׾����f����@�	����`e�nw(T����X��(�-h��p	�Xf��i�ʍP�mD�ƿ2?]�(RBB~'���E2���f����&b�uq
PP�;d���0���qV^s��r��^��|���0�j4�i0��:��2:�M�|�=�}k9�/�=I->�k&PCB`���`�ر��nJ	ݲ~�7�T��0Y�6��R�$�l"��Un��0���Eû	����y�fnrqB���@���Pznp�gZ����w�����ۮX�b�V��
b�Ep���2�h��i:h��P�X���dU(cK� ,��B��+[��#�h.2+�h��-�������i�#������W�k�5$~��(����X	KE��s.��֜_���
�=���3�t�B|��$b�ˋ����X�ݔպ�.`���VG�� ��>~�'�D��>R"cCj�?h�^��8��P�6$N� -�jiV�2c��G)���%=��kҁg[�g܈��&w��:i��&I�m�{6V8b��;�Md�h���@q�:�R'=Q'�6���jd_9���EB�g��䶉�lk�˺��d����Mx4��;�o)]x���D�+���Y�Z�E�����Mꀄy
�.R9#C}9S�1W� �Vv=���kN�7~�����m�</D�*���}�@�t![����a�\晥�ٔo�7X������$�cW�V���c����&(]��I�΋��p95��`WI���6��?���%s9�����V%t��)�d���������� ��"�����|P���k��ƛxtMt`f�����P�2j��g��z�fb�GYŃ��PqV�Q��x�_M���+�$c�Ps�7 8P��Fqq�@D��^�h�����ތ�^�+��	���S/G;��_�z#^��UnT�(�Zn��hk�M����#�x�U-&\/%)�p����ߛl*���zu%@�*I\?t�lZ̍�J�`ׄ�4��"��'꠻N�&�F��8e���8�܀�P�z� C����wE���
���W�MF
��'C��0�n >�F�yK��	D}�M|�����q�B^xzK�*s���:���:���#�<v�r�~�S�[���M$�ϯ���fU[��7G��G��TNܦ�g�#��	.�O�w�T����`CO�2ʽ��S��Sة�����+�I��$��6 �:P��~������~����է_+�%���𮢽 �H[XY�����Ș[7ly�fQhgP�,!��Y�2Ό��gN�qj(F$H��j T�e�k�&q)�I�{��`�(|u��B�f;�?�9��vk��X޾e��,�
�y;�T%
Ҡg<k��El*�7�:�������b�םcХIݪ�9��La.�T���\0��[������t�vdޜ���/�)ҭ�`�at��\r�L j:��}�
��zJ��#<�u���°���>�e1�߱%	%������B���|���*I�+��Rk�#\���Ŀ�p/O�H(|U����YHlWU>����]��z�Z���lݚv	㠽@��w����8�PA���r�X]mk��W���B�&���i�!7u�>"�g��HI���,�P�a!nG�WG?��M��wEGL���.��ԣ���z�\�FG��z֥�N������}�鏹��f�v:�A���]�QB�kak��3�U���˿(p7h�Xm�v���U�c��P��zz�%�G���5�� �1�EQ0�������*�L�;��B�;�8��4d{�VnC�9\��Mg6̦J!�E^U�ևviek�T��x{큡C��|%Q��9��2���֭����t��֪�3d��]���o��X�[��!�0��J�F`����9�*-��!��'���t��p<а����\/}�=��Ȳ]k�H���9�yp<,̸�WR9)�(c��7�Y��S&3�m,zDdB�m�w�+Y�Y���wKDȁc6��dt�(A+�+����-�2��� lꀵ�.I{�c��������P25F��Q<�df"(ʴ���G�k���_{!(�u�81ݪ��Ri����ɔ�! H^��3�\��ғ/�s��c4њ�����˕9�1��1�4�\�Q`c�����%
Gf���[�A�?nC�s�.�!h�6o��#�������A��gс�*ZOJ����D�^��C���Ŭ�g��2���5�kW/d@�{_�_��vy���u��+,�A��<��+a.�d�pb˜X�H~1&Vf���I!z�c����(�b��۷�xU�$	b�ȵ�Ԯqm5��uF��xË{����v+���3�zC/Tl�B��b�j�1�� 9T��우��v�(������W�O����V����\������~�Da1��>�~���ǻc�F�v"ɠ31a��^S���%����R�W�b&{գs? f��N�p
��ZVY�F���Z�'�M��)��[Q��JW�ɍ9�V�K��g�]SC0)G��ɋ�5�Qy3�sW�*2�_� .5qb;a�DW��2��{�]�j_95�H�H�uU�y�dIKKb�Sp���:����e���S''4��	��iק��tR�T��<�6s��Y�=�ʓٝw�ơ[��`_��������e���`���	H��͜��Fi�9����r|��UG�)_���%��nd0�7�$WG��.��ڵo������V݁bY�j��7j���	���f��� ���2�	F�~Ї�Bt���~MҐ� _�Y��:�V���M�R��f�(���2(�Z����8-�������'g�H�c�q<�sX)nq���j}Yв_h��ܽ*Z�$��y��'�4�����\d-aϝ�6F�?�ޭ+�vi��*�a�q�ѥ6�څ(�*L�غ|�|���H�_V��k��O�`�4���~�\�3�T'L,TPs��o0�Tg8M��Oq�,��51ơ�)�����C�<I>�c�TЛ^5�k�pu���I�i�
�ZL�Z���#����;0`	Ra��%��~����;ۇK�P����J�p��l������]
h���[�2�����@ƀ�eȯyR{?�]A=yݰ��l�ŤO�hOg(
ͣ��0ц�ܛ�����g4�k|�p�tp��Q<�/	f��mU�t'��,�>��x�V���~ܚj��IN��K�' ��p%k۝��I���nT�1�L�72'K{������j�.7�����B��
kH}��fѨm��Og�n���w}� Ҭ�1#)W���00'Q�M����(����� kz4[H���8ֺ{?J��2�*~�?�D�NC�{,(���._PS���H�Ѷ#z��̾��E�?�Z��;n���Ǐp�`*派�cj��8{	�c}��!�����4��[D�î��jc�/�LLC�R��@^q�/"i��V��&���"�D>u��V�:F�/,X4�����["���hi���a�4�U���e��8�o�M-k�bg��s4�w���D�6]C~�N?9�s��x2�,c	�Y����T�[?��?��rm�bc�6rq�t-7���#����j-�M����y��P��k�ɑ�n�C|ą�L���a_�4f����u���#J���>��5�b»{v�e�Z�B1�^K-�)~�SĹo�E`�!�yk+��׏�;�/5�sFD�3x�2���eo>d]���lDHp��v�Z����B������~���=@W����F�Ly���M��F�H
U��26���\7 �a���g�y+߅>530�9s,�P�����w��<�\��r�^�5�47�#��-)%`�Y�	����,�qU<�B�=�|!�?�ᕨ��6�"M����$�#d�IH�j�+n��ԤJ���Km#"���ůS��R��VZQMMh��3���:�f�Ue@o�^}�y.:Z�4J�ԗ��ph��x$:tWv��r�b�1��X_��B1�0��Ysm��ԓ�ki�9�bƞ��`︓"B(�GYW����5�3o��N�3�k�n��m	J���,�g�������1�ǌ>t�T�HE�7 ��.�REH��]P!A�t,���_E`; )*JG���s��G�C��P��k&D� [�E�[���h�L!����::��1�)�y�!h����Q�.���ꤤ��E���J�>x^G
�"�L�O������B��̽X�)�j7�����\G�A�6Q�=��i;5��V�����v��<��j�ml�V��?�������%%!`�g�������7j��9*�Fjz�!�*�^A{��Yw��*�yh*"5��B�����6��䚄_��\�������� <�*�U�N��-<��U�"?�*]ʿ�Cz��m湘�Z,j��\y�#7t;B7�%b�`۷�����5p�&>�A"���� l��'@d����E��Ƒ���aam�I�j�����n~�P�/���m���(5�t�F�ޝ�h���
�dÚ�d
d�d�q�y}���n+�]�St����pH�3"��d��)[t�q@���� �|E�*���̥�v� w{�Kkk�@�:c1/0��R��^��װ��|�� ^�z|�`��gz ��HN]x��1o�k�)��>��'8<:��.�7Q�u�t�n��{f���0[e�ly{�R
SR��=��)�&��KP\�� p�;Z0�fF�M������/,a�]G*�7}�J #"
�V����d�� 0�� 0iM�jK��(nPN��2Ӓ��L1Kf9uA�%sߖ�p�\�y�d�ܤ�xA0����2QY��hgyN�U�gz�H�1O����ÿ�7n�M���\�Q\�q�<� WGl�X��-�v[�!��������Ϋ�Y,�*ZC�9
~#�J���2�ҳ��Ň�� ���E� ũ�!����|i��v8H��*fP=	.<ֻ�M,�Tcm���U����v���z�̦[Q* ���O=�_��J�D*��E��-���~&���Y�)9GU�ny�RU����갋�������;E#^b�@g��#�o�;�@��|v[ ����Q!H��]b�����,A�I��rә��ZQϲ�`}�H�D�.���"od�4�c(�5צ�*9�Ns�o��ث�i^��=�L2�D�7#�]E�M��½I�T�T��ܶE�ZV�t�\�Mљ�wT_�+���Up�gL�4�lv3Vf_~+�7���'����=\v�U �ZR����X���W	P1���hɪb�Q�.�-x��k��i{M���CV]�ʬ����a1dQ\1��Cir���n�W�h���r�j eí��,�޽2dN��R��>_�b�]2OzeU^��k�8~v�U@�����B�c���+�d���+�d�q�����^)*��Ys'Y�Q^�G]�*cU�]KP/ޙ���7��I���w_�t~K,���Ƃ�i�4�?�������Z�F��ե�N��j��Y�W
��	Sږ���	,�0��w�����z'��󄛺������D{���Ԉ�R4_��'�& 6L�5��E���t�"�-_,�=C��2���d�v;hu�~�_6���Y8 :yG�D��t�/�c��A��t؂ڦ�-Rݺ+��cbquNE�P�}���i�z�a>���I��OM�̢K��F��d�4Ex�apfo{��E�#�2�+e� ��WTx�2l�貇��ꇝ�n �����A�f�x5��['����D�n��\& ���[R���/K̢D��X����.e�Kz}P��I�D8$��vC�[,/�I�>�f-� ;řT\�����F�+Sk�4�z����f渏�y:˶�F)oK�o<�|O=A�4.�Cm(���/ݕ.���zC�FKعSW��*�C��#�}�!KP�ɏ�nW���5���Y���K�|�suFވ]9`�P\b�FFQuL˔�G��"�SI���x���`1(��:�Ph���N&lAՌ�S�����-yb]2�~H�DrML4P�²IJ؞8�ݦJ�:T���O�0A�cܱ�U/�dǖ��g�F�&�v;v������Hm��VA��aNT����.��4A#N���f�Zc�b�N�b�Q��ZAK������N��Q�\kΒ:����4wU�l���N,���]&�Y{K���Js�lHˠ(q�K�dBp1�-�_���������~ �%�7=�`������޷���e�p���W��A��4p��x�~ݵ��]�j5؃�zO��/.��A�f���ں�$�R�7��N�n|��y���>������6m��*l%��D�g�]�8V��gx;��P|+9^��c(�9~+"ۯ{u�".`�\����/g��0l]~��:�7s"�a��+��7j�������`�����)H��L'v��`g����O��A_,λ�).5�9=�T���b�O�"��s������bP�h2��Fp�t����~��m�=��`���b<��b�=��$�A��|�D�3�	�ob,%MI�V1?z�{q�a7%X��ȺD������ rv8���P�K~L/�,�z�
��?�ak�@�Bw��첣�'�ϕ�N�����k1s�'�݊d���˙����d?�򼎺	���,�~��)c��~�X���&�}!�R�;�s�w�_h��7W���D��_I~�r&*3G�@�2��{5+��xO���X����w����1F��V�xd_���s9�5�y}ł�}8�Ԭ�����b�V���Rq�B�g�E�K#���D�I�l z=ږ6]����7H��KAY.9}��[i�^7��z�}��<�{ �S	qf���C���"b��i6���ŋ˓bE�E��/ܽ}\W���g��3��z�}�},5}h��b�W����Z�GB��=3�e3C㘾	b/&�)�ue������z��B"ؘ�3 iq�<k���P2��c`�|�8Z�S� �X���iJk,�t��M�u����Y����P��)*@ �if��n8�4�x����e�ڈ�	�������`KBg&f����r,��(~��Y����(#Z �n�S�Ao�����ONL)R=�N�2AP���p�C4zn�t?3����A[r�s�)E`b�"�rmI~[sR���
ֈ��ZۏQ%�v)A���IW� ?�^��y=����Rq)��?5�Tnu����h2�"I���~�>��/D�UQo�G�_'�'p�*�xH���}���b��b�j�	\�Y�F�Ә�9��2BN��!��&����]T��&ʘ����Owƫ��zA����C���"x�B)�,�\AlD.+�%��s�� r)����l{�	�j3b�ۤU�WG}�}��KH�����H:��,�"c��1����I��%�t�uG�;��1ӎ�9.R#��ӻ���Jy&�ަ]�6�;n��z��b{���7S�h�q�^G��@6�l��u�����Ư�rȾ'����v&T���3�ֹ^���͈�)�Z�|�[���̓js�>�̠˧h���c���Q}�ЁO�6(Y��L[�Yx�Φ0(P��2p靿�����n��0��c�+�?���+E��/���>%����Ƶ���F���utXv/)?v��l��,?�ԁ���h��ȣ����&B]�]>I8��3?���ը�.�ğ@�*_�Z���B2��m��x��3��D���������9�@���։J(�;�0������U8���t���}�w-�7�M�)K�./��W��Dv��}n&\L��w�"OD�8�xՇ��(�J�����TZ&��Hc�l�U�*�rXs��V�o%�	
F�^��j9����k��|~��ρ31<�������@�>��SE������v�[X-<]+6�#��w�Hc�D��UŨ
L