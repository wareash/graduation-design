��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jåا{�\�u�?߷�dn@6�zf��r������;�O):�lG�31SX�����V��[�F�*�\�R(00Ǧj����]uɞ
�� :7Q�&�xaȅ��5��� � e�DO6d�A����sv.ck��U�O�ugl�A~�~�����2W�xOd~!�L���u?����\QE^��d$9�������� �lL(�����˛�շ�R�X����"��-M]����3}EQJ\O�
��a�WR��iMH,ơ�+ɨ�q�����Z�9�!�� ���`��nU���C뼐��i��B;>���,�>���2�[ƑI�pcZ��;�i��#���^������9��0�(>%�Y{�N��������<v�ڠ�����n&J-���Z�k��{_J����l`�F�oH����4��Zve0���� X�a%SVY�g��+Ya�G��ٌ8֩�����#���Q����q�R����E��hy�۩q#᾽_Pf�̭1__���JVo&�q1�{$���\��]��f��&������3���l!g:Rp}W4�.��I$q%��JUx�E�<��|``��lg}4����~����ը��O!��'*9������v=��lYx�D�e�h��6��Bb��4l!콑_�y�����s6	/�92�*{����;g������c�Γ�#��7~�ݤ�/`�q߱��Թ�)�zN�K������������X����m��+��V�pw��0rB��4iw5�F��O�~�T�.�:Dz���������3�����{�ƭ���֗l[��=�&+��-Ҝnp\�B�q��B����P�s9Dw�kF��ԎϬ2_>�#�VNĐ�n�H�~a�O㺖�j��R�r@��PD�-ڎ�G�hP!l����D���'��)UZNc�#�=����Mb��_?)	K$�C��e�Ԝf�K�*�\Nh!�H�> ~�E�j�Ȫ;^��t<a!qKrѷ��.'fn�{ 	"�mo�͢q$0U����[�ē�H��8��%��>u1�p��.��VGx��jLW�B:8��TQ���6���?�_��h<i"` Ew�I��4bi�^���Qn)���b�\o���"� �����g���[x��ƅo� 7Yi�ŏF!��g�Oۏ&��կ@��3�6�ds%?��͌;�j�_DQ[>�knF�+�>���,W)�+��hع�h�ml��?���8���YuY��SN�nH;���5�.� ~)}��}�E*7:%�Q�8��Y�d����z$����,M����f� L׼�7z�CDxT�ԍ���xhU�I�>�)�]�сhk£�>wW1e �B	أ�sU�|Gy}��ky��G 'Uf^�
�� �169ε�S�Yә�7k~/����t��c����Y�u^�ou̴ky�c����<}��n� s&SY����hA����_�'�ɏD�W����K�s��	�(��vj�`/Z�ɪq0��w�a@*������r����t��s�5�ȁb�t@��)�A�u����y ��/Y�ľ���T_�=�؂%��˪:ܓ�?��nxJ�}���\z�V`������i�J�W�"�T�2Ov���U�>��sn^Ԏ���"b�����0[`>��h��Ώ�f4�����w�]<	���h�k�T��΅�܁��PH�H	�z4�Q��e���(�^��F:��҅��\�٫��J?k2���_��G~�B��~�ztgL�-荫�n2�-d�����=<X��4��pV.}h��#���M�+=o|�E���t��b�-(`B�åBy0&�}��A��d8;��9,w���=�4��@�yaL�>�=��Oa^���%�s��[Q��g�#���e�Ķ1���ǀ�i$�$ql�jF�qV�T���x}�**u ��f�9FI|q��8�rr�}�E��&�='�����[4����;�
���{Q2�𾝝̮yj����k�V'џW�/�:����y� �����P�ZT*���A�����Ό3�񈣽���_2Q֘�����J=�E�e7?k,��X|B��Z���1���m�UD9��T]�v��>�cŲYq���Fo��ٚX
�\D�?N,��Y(DfIN���0�����Z��K>W�����!ĵ��Ȍ���)�D`�Q��~SM]�	�`��;A����"8����b�#�(����U��˓�t�y�S��4I�y��/��Cgԩ����ٛ��qM=�~��5'�P�r�w�N�"���t�� �kR�͘�/�־���QfY�m������~����UM0d�Kd��I�)I� k���:N���ګQY��z�ֶ.���6������"�nk�(Q�˸"ZO���`�F�L~,�&8\X�������I�������i埵(��7�����A��K�ڻ�:�[s<w��H{�Xe
�|9�����~��=d��<w�9e������/_�7t�-��@�n�W��cnvxKe�pԚh8f[��%��TXK��P}�,6M-�G8��,?Fw5�^�v���#���yE��Q����GtED�5�����ڭ�X"*s�)m�R��C�)Ѥ}�rRe?��9
\�����ݢ?�	�[����`6����2�轲��f2�~.�����!�z�r���X4�0j��JxU�2D̻$ H��`�G����mU��p�љ��Ik�z5U�Jt�:��4�#�|s���U��.L^�)��"�u3�\i7mH��F+*'��{t������2� �^��YK��8��0��p���v3�{ȉ��^����2g���H����Z�X~Dҁ��!V�41b�uŠ�!�c�LT ��hO]�6�O��.���#o��ΊJ'+���V)-�i�P���	}�\��É�����Ԓ��,V�v>�2����o�L��� ��j"�pd�Mu;d�.���Ac�X�X�˴�#un#��}������;y��NB���1�U�k *���R�"Ug���'B���𶿪*�$f�y���i����xQ��:��/�S�9�����5�׾��>zR�3�5�1��㽱�it�C��Ĺ,�������J�������X��I�:�54�?)i�7���	O�� @dÚ<�K�w0:V�ǐʉ�X}"#�4����C ���r#�����L�Әꃦ3�`��7 :���@u��1���s��&����#2���������%6�q�w%.m+39��VS� Jk�G��1C])*C�����u��X�ɔa��q]��5��db*I��噀�Ǥg���E�,��z�R	.|%��6���{'�-d]il�|�}$$o�\����e=&��_s�-��Q�'�r[�&bcsш:.)��i6�M�~ԡ�p=w��������5��uP�eF6���ܡ煋�}������&f�>�w��풎HQ@�Վ���2�Ak�i��V�xPA�hf���!�Dk��{�!'X�ډ��?z[�+�k�NR�`�NH+B�Hɿ�a��M��:������|���ό���\p�:>Q�g
r���C4�_һ?�}|��9K�	�4d�o�r�y�)�`���� C~�4]n
����b^�Oor8̰B�/�Pw1��S��=%�y�|�y�$;��}�o��m�Z0X�wğ����Cs���x������c��{���&Sd�܆ؤ��0�ї>�y�GS�_ F<Ba��{�8�g�'Cb&6�Q(|=�&s��P[ ������"4�.��S�����}p�-
S&��B�z$]�1����'K ��-7�.�Cs�U��c1��1���\|(X���)�t���4Ĕ��a�!w<B_��h
zv�:ڮ��ӆ��,'��.0��Z�+j��f&��12�t��Q������~��H�Ɋ��̸��uPz�J;.��d�;���wk{�P!=�D����~Q..r}���G�����e�4�p�3��q����v������2�L2ŋ��ͦ��TV0�bO6c��XR��*���\��ZY�p1F�<�2��88�%���O.� >d��\cB�x#�ȿ�I�?���4l3g�&)
�!7PcCd.�$�ɿ����.̻H��H��b�G����s��Z�[$��z#�e����R[d�Z���\�y�o8�Rl�L/fHҊO~6u�x����r� ���x��9�{KB�������$a�48��q4��ᕟF{%�C':d|��EnQ�ӡQ$i �ҟy�_�kk_��T:���$�9Z�E6}����~4��0�t-KkV�s�L���:�[�d�7��
��Y�wB�Q+Ve���m,9X��%�������/���𘃩0���H�
��qPa�r `�X����c�c9�EOJ�SF[N_���H\f��1��_�=W� ����ٲ����f��B. D���nHf� �1���S|>-����m�[wZ��=����ޏZ���y8R��L+j��!@��/G5�[��cyq�W��#��'ʰjP��K۟	���޷J1���	m�|{q�'�C�{�Կo>Z��g0Z�ɭ��6E_ԒX�t�����*�W8�
��'�!:����s���5�����v�ѐ�v"��4�:��VWA��)�%�_Q[��7i�{�Q��;���=ok�� 7_��G&����s��W���5�@\��̉ș7��>�h�<D�&�����>�K��d�'�Dw��'^~Ź����� 0��a�X�1���I����Qל�b"N�)���Jb9�4��"��+w}0-��$L�g�	�'���n�u��h�T�&y'���`��	K'M�y�6
���xu-
�w�vF�ڌSG�z�	���9B�\բ_���N���r�������":�$�����;l�S�\j>� ��Ω�4j̕�x-`�]ҹ�vW�{�-ޣ9^�=��tp��$�m�?]fT�}��R���lWX������(��Y���8��-��k�aH
FA��J���w�B~�Y� ��ν>n6��_�_[�Y��d5N(y�nk[�Z�5���Ծ8i�$N'���~���lBB)���	���u��ގ-O�! (��*Ō5֑�E�qPwP�V��#�Qi��0w��X��{���8w�����'ʴ̧V'D:���b��v,��|ZӼ�ʆ]����!=6�=�y���3��uF����Dhf���_�9Zl���Ɨ��t�7H3 �1�JR�쑋AMx��2�8�M^�@�.�Yְ1�.�U!*G���w�}�fg	�DN���`�}06���/�(y���,��I�"��k#?S��X+XV�N�.����(�� "4��T�oq�AMߵ��O|N?����ſX
Z��]q��,hkt�k�z�q^+k���/�I�X�=D&���t�)!�Yw��B����Ū�9�K�^�2�ŝ��!�Ciec�7�5h����Jw>���ӽB�|��NfP?�ؗ��А«��Cc��6ᘢ���nES0�/j��	#wHy��&�"ʤ�����)�4�	�7�9S�~��Кy��� ��ZY�{>���1˱,@:���`�vɘh���벶�HE�p���l7�:&q����|��
���c	��T$WARب���A�d�J��C���׌�]'��j���+��=
�Z�Ȋ��G[;&���TB;2�B����|T�x�Ş�|��b=)��A]m��~��h�n��m�wO�f54ck �
��ka����A�X�H~	׮a6��j�@ ��OB��	�"O���
2E�������iߦ�+}�ٜ�f�ݠ�4��OsG�E�;�zl���aF[(�x���'3�6<��<R'��*�������l�k�g�S��8�
����Q\��ܮ�h�r��Hמ�ɥ���p˰2�.0��<�T{j�g;\�E��:W>���l��>-�VD�!R�����"�hT�.?�9oc	`���+���V��Y�t@��nmq�]�G�D����@52%7)D�YD�(�2�ޅ�$\��/�-+<V�"m�!��F$W$�ls��p����*la��¥G38���$]o��Y`O��	{��������e)��� �9�_ow��묘�8#e�qq$NĀ7:d�d��W�b��m���p�TZ��4�Xh�T��&}{ne�<���.$ ���%�mH*����'��/�|ޯO�j/�w�;uk��>멓oQ�]�w;Q:�Lg���*�33R^ǭ��d�cuo�)7M�C�,�����J;Spxza��F`�I���3f\�e�������{�K�,�cF>�����DQ�=��D�T�?�p_�uC�Ḅ~�(׫%�Θ���E� ��Br�����1�8�1F�����'�X3��/��k��e#0�(�d�XS_��{N7|
�P88����#%�����ɓ��g�Ċ�\\6ؿ��GV�������"*R�L9J2��`%����
r5N<60?��� ���/���͐�ńE�>�)�ug��@����}�$ܬ�
�/�����j�^CJ��g��8ϴ86$��CG|�[l��y�k�9$�3j�1�Bv�4�\�;�^Gַ����I+�7���qus�~���� NpFH���-��C:~	��Ғ�X����>"��m���@�_��RD���k��}R�p>�#��'%�m��޼��:��/ik&��=�V׮1�����^z�c:3G���;)$I��y����
BL`�'��y�rȏtF�&�&������QȐ 1��=��uVC[M�L5��;���^c�	��Nlwʺ&�载��D�~�������E���S�<w¶W3&�_��(^�	F��y�aN	�\>,��#*��|��b��蜷�sy�tk�7W�A͎ʚ�?��.|�P�\���9��Q�B���uO�)Tc<%y'k�!h��}����ˌ��A�>��3����Z��|i�Mt�씠���l�R�����Z�u��.�����.Oϴ�4���BX��C�vՂ�P^�u�հ4��,�bK�v$�IL2�#O���<{g�d�@y
�0{	�U���!eޏi�J�r��O�]]r���U�A}�9�DP�ſպ�Weg��m*�k����a�']yg����F��F�6I�j�O�zC���n)�	����?��zQ��`���/���4�����-�w��4XS��ӻt0��UI;����ӯ�c^�WD/C�4Iِ�1��F�။�f(��$t�&o-F�����r5s>�2f�q���(���%L�|��'�	V������O�;��%%V~���:�_|�L�ILj�M B7x���eⷞ��yy�����'���e5�*�|����gֻ��Oe%3L������u��n�� �%"�y!y�P����}R%���?��!�p�+���r,��D�"�J'�e�8f�����ȣ��P�+{~l}r@�%Ũ�������vH(1H�������
h�H��\ScNv6�+h^]�єi���k����C�C#i�ը`Cx( %OzQ�|�d)�9�cݝE,�Z�u��YY�ݹ��L�$sp���c3��U���<�b'��=�gN�?�!���Bl���+���Y�o���a�K7���l���W���9\f��ʠ�����-�#�Rs��S½�)�(�ǔ�6Q��sǙ��A&��He�V�Z׏Xx�>�������{_ct� >���G �&�^9��Tg����r!�6��c��uL�ɚy��J� �G�x#�oQ�aӉ��T=F~�h�c��T��38��~o��>ʁ����_���+������qj�璡/Ĉ��I�W�z��"=:�7�A�R�3�����v��NO�3�N�hA���r\t��a$=�+ѱX�20�w��Kd�>U��紭���3+3���&��8�K���b�==V��q0ٵ�F�m_%���8�!*��7�כt|q5Nc��\�rN/�9��0����1��7�TƉ{���(KAV[���i\krfj8G���������F�b���T6ܢ6�p��͝��==Q	� z��$k�ݵ#- ���Q����j^��W��"pb�7����Z���v�� ��(�mF��i(��q҈}���ΐ��63d�D�~��^8L���*^ ��U��Oߣ��8���
	+�D]��UDT�����