��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�tڐ�!��Q�����xZ�H������
��(��B_K;bA|���.-ƍ�B)�wr�q�h1�oDu�j`�3|�?l�d�U�J��%��{�.Q~Ѻ:��E�)�֪�3��g��UvT���F���ћ�2�&�7}C{ ��e�9�W���Z0bnf�$!��k��F��B벭���49	vr'�`���H���rQ��'�/��<"Q4��N�i�ۣ����� B6h��_�M��'cN/nO���C�a���}R:����Ķ����Nka��q]�2�d�p#*�L4��'A�D��bU�u@D5P�T����?�w0C����PbI�i�$�8~sɣq4
��Ti���9�(��"3�|�ƻq��Y�#ǁx>�*��ꃨMdF���(��Vp�t��5Q0zZVDX��#�)h���+�ߐ�Q���#��lK�Gh�?�R2�C~6g��/'��>c�L����������O^�\
�T�㺚�@�A�u�WBׄo9u�+Zo�Shj����#CcqĞA ����]8&�@M8��s�U,�^���3����%�H��_����L��uR��#�[����٨f�_3��˂���F�d�̲�a����Lq��5�
�HfvU�������O5�0�������j������h�MFa������.��P�%�עq�J��M���F�ƀ�PsF��z�)4�mT#��\��ؑ�QX�T��Ǎ���O�k(+M��`3���nj=��Sd�+��P�b�Q�����ޖ[�� �l��BC_:E%n8�(�e��"/0/1pp����G�Z��~i{��o�4N�|�W9:s�f�6�xfg�ՠ=�#[M�̌�c���m��(�*h�x"���*�����OB�4��4qƼ>�vW}@����n��$>�I$�ʽlZ��aR1RN)�Z�"����~�^�p̵'B������x����Z ]�9�� �񹮇:�T3����	�R�dt��	�Ē|����
�fRYڑ�u;_�4�94`�CRB�_j(?�tK�?�q�$5O��PA�v� <XR���+��fDÓ@d'v_����C��Ӟ�-��<�E`2�d9)]�H\ �i��}�hy���5D��F�x�I%*!>J`/��iL1T�^�&"�;O��k� 0}q(p��Zތ>�!��WX����5� j(����5�_Hy��Ŀq#Z
1.��3�)cd�%ϓk�0w�py{�GdYs�2M���p�oc���,W�LY5Kr]��W�Eꭰ���k�=��TA(�-^޹��!�N�pL7f�S�D��Kq�d̔����Ik��������HD�,?7:ФCd�$��C��
 �Q�Zegh`���ҕwu���؃���C��Ӊ-���D`A�&V��q�w�v���PR^_���O��pq�6�vp0���X_uh
?Aq���>+<��f� fyXw@&���Q�h�C��o@�W���D���;�o�)&5����fT��N"�GW�b��b���}�"���+<�j%��� 0"�kHPD���bm�%�8$�� ��Rh *�lZ'ǧ��y�M�)=~V�
!�ͅI}��o��cUh��8�0���] 3�� *=!	-ƫ�-H��{)h�u��8FQ��x�i�ve���qS�.NԲ[V���?]���;��aPd2E7ɳ]���51(c����^
�B����o3���i� (UwI���s#��})��'C�W?Q 	Š�t+���+�a�O������Xa2�Q��oq� ���o77�G�
8;_C��1���޴"#.1�
Rh�b"˲k���ή$�v,����ST�.o�]���5iH�sQ"[j[�L�^�:�T��y�m|N[ԉAa��Tx\C	�9�	����G��Z>T���P�Ul7���Q�6��v\�eE�c�"�� pG�-�S��� lh<ƙ��
ky���(1�צ�~��`m	���H#��<%c���fpH�_�����"ِ�{j+"��7[��l�P!e���. X���zq�O|�/0h�����������?�4��
(/�9��X@�61|#�ß�R1l�G1��Pxf�o(33�F{�R��XCj����G���~���(GB��b�s�����''h�i�nY�vNb�&D�̳� !F�