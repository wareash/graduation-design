��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jåا{�\�u�?߷�dn@6�zf��r������;�&��0.�S�H�%Ѳ����C�C�����t&,����,p�23Wpݲ�/��8I��F�:��"ԳsnƲ#��4�n�
:����y�o{�K�y�*Tغ���{1��I�݊ҷ�DP�
����������f�>�w:�b;�b�0�$�V�W���o�6�}��ԛ>�M��s�����@�4�T��ɼ�^u�~��"E�.������`m���a�9�~��|'�;x��=�mV�`�D���"�\�YޯMr4��d������\�yS��f�x�#3��Q���0�i>��f�̣z���?�'K�T/ ��g�����Q���!�^����o�_7�>A��S�/�˰����POU��0�Y��s�dZ��A[V#5�u_�e���ac9�9�g�-ǭ[W�Z��>��0�|����ӆ�*D���yH2��~
i0���Z��jyHÔF`��z��m�8]	R�VA��T ��v�5�v�Ŀ��kEߡ-�@��0�PҚ,��1}[�Y!-5[�Ȇ��7�~a�c!X��i$���j��kI\U�h�� `��,��q4-���|/�`l�g7"k4��4��S�$��=n#����~������Y�b����ƭR0	��f^���/?U�2Z�Ѭ$�J��\z�$���������]��r�k�-m�p��-�����4B�IO]C֥�#l���l�][�My��Q�3�������{�YS�����)�#D�5�ߚ���=��M��R�[�j���)(��O���3������ʻ4|]���ʵ��<m���9K�.�f��U���A�+J�;���"Iehۣ�H|Ӻ��Z�Z#w ���^�]�r�dx};�	zP?�+xɓM^��u.�g�}}XPJ��lC�ae�讟�\N�=��<d��zs�,hF%K]��bS�}�����/g�l���[����_c
�L�s�����Hy��W�)pr���ٚµCMO�)�ۨfb'r�{X�M���%���g��b�3���b��r����3�#��tL���l˯��M|%�''89��+7��(ݽW��/ Қ�l���G�ɵsp��_�u2��R�*�p��Vo�V��,Mm�а�b�ץs-��D2&
�}���>f�D���	\+Nt�P�Bx��ͫHQW��Z�L�W�j�&܋s�� �oe��hحj���.�3��7��r b�GIW߮���l+i�<�v������ZU�P��j��9��o[�����:
��i�O�"+�ӱec���O��X��ıiE6��w��i�	��I�h�P)��O�mA����?n���R��k���Av;@L#�$��fj��% �e!<�?�@F�{���#�&��پB1�uYR�S��Nkfl��t�<���)���]�jY���e�	|��Z�_0�ܺ4�Z�?į}��kvr]�kM�8б�1><V��.=�h���ԯۜ��􌾟⒊�|�� .F��w�O�"M�`O���D��C��֜�Z�cA�ik��R�����>2�"�X�&r��`TnM>���\�q�j8}(�ӆeD���rT?cֲN����nF�5J�!Q�0e��V��`b�1��Ic�!XĠ݂��v�$M+h-�unAT����<�"�d%�#���	״��,/ͼ׃�����χ��Ӎt6����"K�e���~�B<.0���b��#k_&:�9�c��}�����d���	�)39�L4�\����S�� NA�k�/ٗ˰s36s@�i���L+�@I�5/xr���|:>@â2OQ��;�DQԓ �&G�����,"s��h�i�'���
XdkԳF��}�`rdw��ڇ�"���j�!�Sl_���-W�=�����^Q%0�D�k,z$��1G�,�3{�������[��:�E�ƴ��,M=w4���o�r١�(�om<��ʲ����z7�ܹ�6��=J%���"�Yqh�O�RM�E��|?��~���Q���
s� Z)A�Ŕ�+���	�%C�H�
�7�z"��]+6����*�raۗ�#��<�$v�M�A=׶r�}[����;����1KRSW(�C�cn����:Y���j[����v�:rS�l\;������8ca�"� �D��K�,��D����r��]���e �贳�<yJ�Z�5�,P!&@�w��/|�m 1d�~���(�?��^u���:A�^�B�x��TWG�q��"6��lh��f��S�/�ψK@&�o��V���B��{SK���7}h���r۴��
3�v&�@�`�f.%���=�dv����<��.��6�j	�ݱ-�toz�f#ƠDk�µ� $�1��|�
݉أ�� >� d� 9 >���j��r�$��yX�.,��!-�@�f�Wz��o�4u�j[�̸iNJ��z�;�@��{_lW��佔|�B����ˌ��iEC��[�S簻\]�ګ�C�N�+��wh����~�� �i�UY�����MUNo����ik��¦�K�#�C���r�}�
Gtt���m�� ZR�ͽ���i�7,|����QV�e�.F9�D����u��]"�f��N���<��`�mEj�s��4�x��\�NE�$�u�D��P� ���p!�+ZK}����1��W��"�(F��w uXi��Eg8\�*j�����0��`�(��`��IO�K��#QR�"Kύ�[R�U=�,D�i,qPHT��m-�8~p�|ķ�4�f�9����kQDEЇ�fq��vb�}��E˳�焮 Z����!�G!bp����N:T�����v�}@��+ٷ6�?e}%�U�Ǳ�z�F�)�dA?����'楼2%�WF��H��M����9�2(2`��#*8�!��,]ƭ��
�jː���"�#Q,��59�jp��n�ZQP�׶f<2u��xn�$�gfD{C�T�HI~:TQ�[�X訰t_>��������%,F��b�D�'�մ�ɬߕ�����!�N�:<��W�	��d��"���}NsXL<�<�{�<t��2�����<�/Z�-���K����C���3�'۟ D|�C��,P�Ew�=��`��W�r����dw5���y�&k=��vLNooYb����7����z�Sr�-�Z(����Q��Lz/*�8�֍p���щ~�z��h�ʓ!qޓ��M8.��g3�M�S�ٸzO#v�\֢��Ϻ��f~XĈ|��,].��.d=���/�i�&0*þ�/�&u���~�Q5~�n�ӝ2ۓ�h{䬪>����u�b���I�������&o�Mox[��a'����q�;��ӯP�y|ն�PG��B4/�k�=X2$ښ��}*ep)VIA�oCS�1����Wȳ�I�ōd��E	Kwg��Y�?�hq�/�3�c�.\5S��8����o��K�?�SN&ԏ�i kO��u�H��`qʹ/1�!�hw��Җ'Gp��A����T�[�%���QA���w\ǫ����k�E�?P�l&����w�����-R�Hґ���̑��<�kl�]7�ط�@�\̢$I;{x���B�e�.K�=����.Zb��eU��o�W�؃��G�m� ����QS�+�Cg����H�s�Z:-s����5@���NZ�ZiU�"aYay�9�̜ �d̑l�������Z���]iK%�����[���քs$*`�.���p���
�^]M �'3���3c�9�|���>ULPȾ��&����]��Mͨ��}��1-m5l����>;��\7h�����ƺ�XU����D0¦<������ny��! `���N���6� r�/-U��dE�m4*n�X�:�y�|��^& a�p��i�[[\�I��"��߈3(z���{*��V�[��J�.0��d�����a��3���Rw �Z��h��\�>��ά��L�4���dȐ JİSZ肽����~�u$�l��m�ABr4�F���8�\(�n�d��$6������͡�3�~�@�w���V��~��1�I����t6-50�mK����4�y����E�d�ٲ�Il�ч��7K%����E�1c���ݚ�B�'.�������o�!W�ҥu!�4T�+A�Ŕ�8��ǨGR㸱�%��A�S�`�!��|��}�ȣ�`(w�/&4Q~J�?�+%�Va0��+�!�Lk�e*W��q{�S��_L/���+��i�=J�X�"���:z��aX%&��_se�a�S ��,���(e]���ъ�Ƚ�6��
�.:�`��ze��A���}�ru{��UY�[�'��M��=��|\}ȟO��xtAv*� Sp�J(���ܵN��������P�@�U���\��4#��=�hr��mq�m�Ζ,c��6.Ƅ��/ʯO���נ(�_��nI���:"�?��t�6E0��2�����!펔������Z�R����		0�=��ڽ��7�}��ԛ7>h� ,���������)��_��^�!W��o{TN���%��EoY;N"o�͌�����SM��Te������a����m:,����xf�)�sss��|��:��C��>�6��MFY���=}V��C����i�zE�B:4��CƖ���]7O�c�j�|�a�7tz����H��$ȣ۔�)�r��o̒��{al?�E�R�{ ���&�݌�Lg�����m�m+�u#���������q������bd�@��7��y.���:���+)�˭�YM�81g�� ���s�n���z�pS)f��F�wQ�5%v�*�,|\�i��p�]��3JV5���rS��8�q��d�o��p16�o����8��+����w�z�ފC�!W9ͯ�h��Z@%Sf��~P�eC�[��B�0�`�x�C-�n
 ����nt,�:�K>���E�Ҍ���>��OK���ZS�cp`��6G*�A9�.̮���!�d�m�W��*;��m�F3�b���Y�������~�%ĉ+S����	m56I��ow�Z�σ;�q��:u�<��*�3'	���^����� �o�GX����Y��rLy���J��<���2FZ�Yӕ��b����P����j��}6Al��y|��<ɥ���;����-��ݷ�̙bJ���ܘ���g���zb��gHm�	��)�;�^ƙ��@�_�&}����O'���bM�V�af��w8�C�vX,��O͉�����>��T��G��h�<�����l� ݃���� 
��S>�	bDgSB^b����OU��4ѿO;n%Z�uqr����ո�E��p8hN5_s��zʳ��p���H,2�M8g�#s<Q3Zp���J%�%f��Z`�҆/Edm%!n1�A?���/��w
�@���䕇k�hX�Y�H�!���9~Z�{�b�i�$��y�z�ϒw�$�i�I�u%�o=�Y���0�ec�c˕����'��r����_�'�5������	]�]��0C�����f	�)H����������>ÔWO��Q�4���N�"�0���O�xay{'~���h$�Eͣx=�(�����o�q1�uY�~;�>lB+���E�@���A���[�r��r�=�!��Z���!�o9B��:�{�]we���U�h����^@FN����	�R�������յ���m㺑3g����k��$`�ʙI�3�8:���'>~��˴F�]�y�[�����A)S��̟�ͪ3�/Ϊ�x!cX�$u��1]�t8E+�k�	�����[����U�{)��\���b�U�3�CVY1Ա��FjI ͒�=����c��<����V�t��\����]Ac]D +[�g�M9U^���L��:L<|D�($�O���L^|���s��)�qp�.���Uަ��[t�2kcB)f��ъ���Z�S�\Մe�]�����Z��K��#�8o���u4��3�]2�G���lG%��P{Y;�d{�P�]���nP��#zC�j4o�/����!_5����p�@F!�}0��Kc���d��º�)��{3��V�� ���F��	�H��*=>�W�-|#��n��}:e�/���;2��'�r���-��dvm�s�ݽt;��� �Q�5bgx&�+�� ��ۨ_a3��=oOn��1H*8(�|)%�Mk��� ^`�4�5Fl0���\-�������Br���p��G[���Si��\3�N�6U*5�K*�^�*�k�	�2b,��_��GM�W�����ׂ�v.DrJU�+D��*hA��~9���v�![�UBQznP\�G"�S��?�טO��	�Z�].��_�z/dBl�
���S�l�9F���Ey�W�	�f���2��ֆ��|�e�d��b�7�r����!�A0�3�3}aQ��>��v��j
�V� �"*�<0�)ތ��b�<�ؠ���e�47k
RE)n�3��[����ړCA?5�W��N�Ѭ|u�u�=`��W~ݔLy��]=�'��z�bJ�֞���NI��Vq	`��
����Z}DqY^���Dyj׬��dd#@vE;���0�����褜�<'�(�NR�R_�X��)eQ�p�<���;��3�Y�J�O�O�����Hn(�%{H�0���r�ZI::&m��ޏ��I�	�J�&h�F�A|*��U)�-��N�u�y���N�6�j���p�-`�΁�,�W���k�	�.���;�&@AR�)/�ϼ�l�{�w�+�����RT�de�C���Ī�
j�i��������GC�>F� k"/ޤ�-R���N#;��T�,Y�{-$[?��ἂn�]Y�{�NJ#^}��[j��q�����F��1WM�zepUX�;e��m8���������ʂW�2�R၈5,�JFZ8�K� +����a蕃4]�A
>�ȵ+�O7M٭y!v	�"�UzpxDǠr���S��Ԇ��~>73�B�����%%��Z�떔�D{u�Q
��Nsh��3��4rsw��MG}�Vxyer�I
�&lG0 ^�}�|i���O߁��^��qB�\Y�J�8�ۤ��l�fodiL��&��#�����P�Z��w��m�eJ�O��:�R��!�u�������a�~-�$_�'�o�2������{�Bx�Ƕ��p9R���$�%@�	K�II��i���TuF�d�2C��w���+�ٹ��\��_���{M-~r�=�11�=�x�i ��Vۧ8�RN8�H�Ư`�Ѫ�R���^Y�:��n���i�*@��^DX���'v4�u�u�=CE_�.�(��`�}z��"���d�9|A��]��R&u� i��1GI����'�K-e�s�rjUf#c��^Ҷ݊���K��-h\��wF�s`��3VA�� <���'!P�R��H|��
�L\�}9����5�p�./�H&��8
e_`��̏� �� ���*5Ħ����w\ǌڙJ�ʔ��7�<��n�������%<.�s��.�����J u��r@"ݖ�Q���k��Jk�v�'c�!�~9�D�`-� �fP
��d��(�'���
n����]6=�&j~��v-��26����<I��S)��z����T2��bȿN��0�[��6n�N�' �u�8���S:�/���~��Q���
�e�sA�Q�p�X��Ei]2@��r0��W�Tk� ��;Jr��f����g��d�qW8��&͘��Dc��������A
����$��:�i��+?]�~�Ox�S�=�B^�\�$oW)S!�OH,r�r퉺ġF޶ f�f��-1���mR��M�28Tu��)y��%P�� V'���{��˛Qw�@d�y�ɤ��Q��}G�
;Nx�zw_�'��u� u��a��='iz턚��O1:�D΅�H�3tI��Y8�k���� 5�l@*���m�  dB�N
��l��Q��B�Ћ~dºK�t�V�Uf"+Z�N���:��hٕse�N�{&Bv��z�|ξZ�ru|���T�
-v��(p��0H ���M�zC�}���d�6A�������Q��>�YȠ��+�<O���e5�Y��qgl!�>Cޭ4�e� �%("�_�T���w���EMg��"��<����nLo3Gzm0(\)@0��~��#��Q7|��!H�ONy
�����+�1�EDQN�uھ��	��H��'�z�.jN�_F��ʛ*t�m�M�Ȯ��|��@b�H�A��+]4���Mr��}���5\z�ꃨ�lSE>�Z�̦��:��>\����+�8�b��&i9��4�bm��nx���z?�P�+��h:�kG�9�o2U���J�@kO+��[�st��"�6-�A`�{��}����zN�5��x��u��)�68�t���D�~~<�z�He�+#G�Ɉ����)l��4�,3P-�tҽ'/F�t�
�F�=�5�����¸��!gS��y���B6��J�m��A\$OQ�Ȉ�� %�Y�+�;Ӯ]���6��(�K�A�'��_���@�y��;�lԛM�/�%��h�$0��Q-U���g�G��5L�Ϥ�R�a^��kQJ3�h������8p�N�����&j�ʹ�/�+5 8��Q(�JtѰ�L�-�kq��܍�y��#�Hb��_GH�爚��C�,W�:�Z��yo��;p������;R1�\&�j�O^����	�(k�/nEq�[�"��Q,���S"/�P~Z�[���J�z*���]��wPё&Y��AW������fL(}��&��j���h����WPrb\���Z�6����os\�ߖ�ML]�m>�I�Q9Ӌe�W������cb�����R�eu�A����i���D`
c݈�J0��O�u�B#¦3����u���5R���ӷ�S��q��*X���!�Y@J_��{�5xb���ӭs�Σ��*<P�/����=��4�B{��L7��&���"G�2�4V��f���#Z1LB �ڎ��4�w.�Y]A��ʮ�@�(Sy�0c�t���h�`G������Iw���Z�Xi��G �gD����׹���rw�p1kU�v��,�}��i�w�u%��mK[��W��<���a*��Ӈ(���/w��
�� ���ZB�HԲ���%1e�aꁯ�`ʿ����o��^'�ҼK�\�n���Z̩q�wAq���c�.�"*�q����E�E�Q����;~��9* Cз��_Ȫ�RPz+qbY�s��y,��������,��e�(�����G�����;��V�>)P��Fn	+��V�E��a�aHKq�.���u�>��1��@54i'r_p��.m����a{8B8bu�t�����R��v������ٶ���lX0Qz��g��.���:�g�l���F���o/�k8����OC����p����e�R'?-]�&�(�b�׏ȧ��|����(�~w>�-����t�A�&��cr�A�?�v	����ܯoJaI#<w�b^�7�5(4g'�a�T\�Ub�{zb{���������|���	��@N�,��'��W_{ߝN���"flv(Jp�(]I��ݮk؎o��C��}�����n},��0V?y��VmfNv]�7����ly�[���2^[o$?/;@�ض�X>��m9Ѭv���*n�5����s_�� [{�9�qזЎ����?�Ȗ�c�B��̯C��ڻN�b�t��ٯ�=�5��k,(�&?ŠhP
V֎�\��n�k	aA��O�w3�c��Q�K��h ���0@�{��݋T�򤌏�"c��+�e?��.u|�e������D`��-�<���5�v �"��U����^nq��kIs���ą�ﾀ���������<�Rҡ3JE��[x��p��a���_�@l!�e�	b�v	}���h�EKϵ�HL��k&&�[���$�;��.�.�#��&k���K�Ĕ�_j�8���Ҏ[�,�VD��#\0�ɔ;�t�ނ��%j�{Ѹ� �!&^r�d%|+���/�J~"�Wi����b�9�[�ح���Y����o!���B4��NP�!�v\�D��i�C[��P��/{��%
�����
d���+8)��;�WTn�����r��L9��g3�
���s�;�1�lݘ�ڧ��4�o7�[zl��i�_�}Gh�XBF��TDFO�O���{����8y�.as�_(�⇥�m�pl�����(Y�1�@�x�֘�(��x��{��?���\���ﻢ���#ϭU�kl�P�kX���b��!P.��]b�pJ�S�^���k���긱A�ǆ���7�k�fZ��蚰��`�ɾ�ҥ�3&^ y��ߪ�DɿQ6�>g �Sr��.a����-�ԅ�՘�n"��y�㊱������K�ːD�0GBœ�3_]�Z>k��M��Vo�ڽD��W��˫����̣�5���괁Ϝ]Ӥ�o�:����&�(�U5���h ��'{:�$a���ᬠ?�p���.8u��*��N��B�j���4�ެ��/�b�R�J[�>�y���W��8+qK����)�o�W����*��"{M��Ή�]���Ǆ^:����o��Iג�]}�� +g���ĦL��^q��߱�PJ9V\+����~�UbP����	����*�,k�\�+j�YRb��O*P�Bpd�iA�p��P������;���Mo������].:p�_�J�<�W۠4o�<38���ـ�Ŏ@/XQ�ɝ���H��bBO���I�/a���*�`���P�t�KD���FR��.�$��o3>E�	"��	�ܮ
=~�ƌ:s�����
��c�M�>�d�<�_�Z���6��8k��!^9���w��;�����	,��z-�N�II���S��C����5�e���]o������ѸYI��Q]<s�qZЏ�&�<ܮE�sA7�.?g�_��Ո���0��lG�+��pn|�۝�9��a��n��ei�+����מsܾj��L	=�_���q���i��%���I4�
F(�Dy�KA3���e?�.�4:�,��I~JZd�@Z%�|�x����}��L��br�>��[坖��A�|�����-�j��Hp�F4q>wz�7ۯ1 ��ҫF�Oȧ��vu&�}%Ait�O��u��(��@+T.;=RL�E\�� ��u�G�[�8�n�<��[Pb-2����>�9�O}tz��+�Ml_)�ض�u�DZ�E�I�c�8F7X3@��?��-W&��U}�A��⇹}Kp�=�}a��KSē����B��3��Wb���޵�A��䌗yf�H߬�f��P:YljM�W�����:�c�_�9�%f�T"�K<����a��i|'��ԽKu�[v����k`������c������Jjz�?Z�%#���|��cOr�u,���X6�Kr�]����D����"GQ5v�c������*r��TI�v��ɧ���圸��fjFgd�Ru�� j���������-	�7'0mX�6{a˓/|q뛗�t�%PE8�IWGu��8�^ _h��Lk�۳�o}:R����R�\�(}@x[�!��Z��m��V�p�Z��P���a��9�ǈ���D�680k�i�AǗ:
)��f�@�ݙ�����H)Q#+)�'Q����������b���.�ǙP,R���r�Ū�@�b'D*�K�5ט�e����@����i�Cdnf:D�4��B�5%�?I�y6)�!L���ɋ���L�þ�~x�;��b�3,j���+4������m�G[��i����FV��7溩p?h��@�g����L���"<s{^c�$�(�(*����0����v<+RTyW��i{xH4���?��~��1���������f�c1o��}�Q�U�ɩ3���L�<�`%ݨ",�����"��������.��T	S�0��J4�{�y��gd��0�*�,��r�hs��q�����{F�m_��ٹ��]4	�=�r�<��#�ʆ$2�7o �;��ߦ����ip����P������4>;�A[�>�n�]�]�ݴ�592/�9��)X�,9��[@Ta4�r���m�ʏ�ѐ�(VЊ�� ���M�&�a
6���8�M ���٪*�`��=n��[ic�
"Ļ��4���z}%#��J,�_��ų�lL%0�(�|�Bq��-�{gaU�fѥ\"O�qո�.ʟ���o�NfC�`��"��S�A�� �*�w}*v{QE�g�f��O~]��T��I��I̧�;����TN��+�"0fh����K	g�7f�0�b\ܗ!p�U^#��7��6�xs�$b_�V߀�=W"Q��P���P*k�{䟽��i_�LpQ���:�g��0|PT��Mc�q*�U��t�2����yH��Pܑsķ��@��7V����J%��^��0�q��3��^�!�����5G��$�p/�q۩d��ݷE�kXl�~�����݆p�Z��̦��4�pkd��nr,}��&6�>X�Q�vC��&�r�C��)�]��7C^OxA%���)G�������_���8G�C3�ƏR�� ��4�s]#֛0���ۧ+�]P�ߟ�����~oM�P2�TaJ����؀�X���F���y���&���i�4�%:�+l }����
m��?"�k	�V�g7��rP���o"G<lT�.̑��l�:L��>����w��B���R8C��|U����Hr��ƻnB��3�P�N�{gx?�_]h��h"�cA��ŢD���OU���E(Z�G��d��6���O�H��[s��-��wI�~ګ�����X���;:��-0s]O��� 0c*[óˮ�k7~"��%�
a���ͣ�y��W��yƨ�`6��_�	/q
�k��ڷ��!m��N�17<J����Z�C��Y��a�����S7�ص�u϶�(���
��$��R��m�
%R��r�|\u�Y���QƬ�����(�IH� ��*�a ����p|��*h���gZ��G��������Tt�{ ���m��X�����J�My[Iײ�}D\�ɇ�t�b!�����B�y�� ���Kf?ڧ��J�Q��a�\�9C䗶�o{(��/>�"`O�P}ȯ�2#�N�+x����7�ְ<E���}����z��\"���Y�B�$ϱ�<#(�~�VMڝ�J�P䕅��TA�9�	D�]�~�1�A�}L�Y5�����v��K���Е�U!���t�\m���m��d��ch���O{[���#�x٘�/!�n�����Q�O�⭢�<�������^�C�G� �3�j��^6i^E��:+��������w��g�P�L�7 7���/}P���^�������;gWz�P�T��ϟc�Ƙ�X3xYk��0�4*+�H>כ�n�Y>�����ʂ��q�*�%�A�/�Rv,JY� �t.	�4�� 8�Yu�d�ډ^p#�u�a�m�Y��%񑃄 N�7�.�Xz��h߱�ǫQ۹�[�H��hI���+��M��M]]М8_"x�E�V")����
�Iw�;�¬���2NL�;���(��[�0%���v亃���M���UQ�rܧ�`��r!AP-Zgľ*(���o7<�B���G�{�)O� U�;��çR�ς_R8���ٺ1$�-*ɹ�jM#[��]�a9��臶^ZF�;���{
d�1��P�4����Tܾ�h��t�9@���, }
"�![���42�1�8^�\�����Ԋ��|�V�bJ6����q	��-�|P�4��2]"Uf��IK�#�,6q�_��[�����k�m8��,�p����s�� �/�<W�/�C�ك«���In_e��w�U5{_�$u&��Y���ƿB5(Y���,߉�3a&Z�
u���Oh�E#O��4�D ��c?�ؐsٶ⇗�C	>�_�H��D�%Y�7x�e�Z��{�O�������i�q�z�@zb����h�x��
\�̱�Ze�_S��L�I�O�S�����s)�����qS�&>o��<Cm�{�{��Dl���{��!���x`���XIC����#n
�A	�_�}���PZE��f�\��8�߄����Jr�A٘x%���FR4�QGj�>�z��T�q�yL���p��2>��L�w,-�h0�J���3��A��`��ҁ�̲�.�*�.��0��@cd6�)��Ya�_Q�޺|�����{T��/��XI�k]����C�K��R�����;��Gdd��.-|r�L�V潇�y#;k�v�ӐuD2K��ҽkڇhĦ������N���� E~�ޓ�ƣ��K�@�#\�~��)��e��EG����F��������������?T�y��V��F9�} H�{�L���}9�ar��oŉ�*���� (=v[�����
��\V��>Bd�P���v:���ch(�'��CNͯ�����˪�����$�lD���ɺ��'v�L�c�c��PXA,ݤЋ�VD�k5{���"N^���
��l��U�i��7ރ�,sm���Ow��.8Ss�?��u%8֯g0���7���ff��c��0/(8״��#�� '�?J�� �����,�p;�V@r�ɶ^s�G�z�TZJR��!oJ{4ռ	�Q�+���6R�?$���L^G-췤Jh��ic��5鋔�oAn�h�MOE2?X��<�����G�K��j	�|'�(���������FV��l��E�!�2��kMtV��}9�bЫFG���>�\�ǲ�'�?��+P�='�U=��p ޖ�h���V	�I����Do���p,���z�Ei�:m��'��ׂ��Gk�&ʹ�C���d�S,A�!aKpڔZC�b-���@�l�[Ĉh���4���L�R�`�T�i#R��%�{ST�5��q�=�r�����ݝ��93�t%wbvQ;Mg��yj#X�O5W�.��E�@<�퐌�i=:1�ܶ�����z=�[�2�f[x2�$E�s8�j���n|��:��Z��3X%��_$�l�� !q��^���M{�Ç�@�*q`F`w��XD��;8f ��t;�_�5ʜK�"F�7���Ҿz���l��F���p/Ӿ�R���� ~��Εx���$`" D���ҙ��H��wً�f����F}}�Z��[l&����0����� �`;_W�_4oKYc4�e���	s�s�$q��*�R�m�w�[�z�
����kt������,ڌ9�\�6��g�R.�P]�0���� v=��j%���ܐw?L�1m����C��@H����G����Ĕ��_����ա��~~<|��![�m�ZuE`g���J,C��I4����`V8v��pn�������z��|m0�L�c����s
�k4a��~tj�ߓ�5����B��O��֋��>5�d�&.��d�?<�%g�����a��yݻ�9�V����wg�v+^@t�|\��j&Xf�C��ɥ��TyuߙZ �+�����]����Q`r��Y��Mnq��͡a��Ñ&�����u=���$�,��������xU���ʖ��YBڼ֬�9�x���-��9�FYfbb���`2�7+;e�@�~�_�� �:�sb�3��J�?[j�ت�'$s*�t�CyfW�ns!���5�=�c�i�E����,�������Y��¾�a�&/��O�K4��[�p�����]�: Ȗ]�h�H��hl��ke0�^]>�KOݣ�	��7w���Skb�c���V���D.(�i�=��+��%�rdњ`�W���`�Mle�H�ۘ����F%[�4ݲ#.6?�X})�⩂1�e.SPN@ʫ�X���oB��߂������k�:��B+����c�W�E���!��7Au1�d5}�Z1��Q
���:\�/�y�D&������4�?��P���	�r� /�4�f�V��Q'M��8	߻�e�����>?>&擊~xG�`���m��x���s���Yl�Z�Փ�b3"�¬@�Eg!���X��������kYl^���}���$W&��迨�Ｐ)��H_�6%���0&髢0qU������+7+�K}[+���c�#�]��f̾��qȝ�ʥ����)<�!wO3d�]�ӓ}j�Ա�\�ܖ��y��}��߁t��A�@k�Y5��cU\L]>�����X��hr��sԋ�p؎[L^�iÂV(Iܾ��Dψ��$�|��*
�u�FS��ޫ�����R�9��r]c���*�l�v���bbٳ k��~x0����b`uH�H���FWD6�,�ee�!�z�?C�Pr�u%�̱�e��ڋ�~�@`F�Нkۛ�_���y�p����&ˬַ����Q쯱����!LX�����Ԯ�����<_�T���v��
�#�s�iV�R��uE��К]� 4�Ҋ�c�8l���#
�V�Ab�o�������0���*������Sȵ��� �xՃr#z\�7��1)���S)ѫ"�jԐB3F/��1��@���vŝ��{!,/k��͌|i}�P�� o2�w���~J��7O�ڛ�(L��j$��| n̩~���++�xt�8�ʿ�Vd���˚C�0����'k=�
���gq���gv�H0I��_ årɹ���|�?���y��}�x˷�;8�� �����(䏅ZɬR�\��!Y���+��k1]�W�T�[�Qp��?db��d�d]U����`����E�
w���� #0�?�<�sPe��W��p@3k_��0�$�hZ���حP.���?'�)^��#WOM݀��J�	9�h��R�c�:CMu(��&�z��|�
ˮ���I:ޙf�ǣ�&�ٛgV;�r!V��!$�p"kd���]$�Xk�wj����B�㢫q�zQ:�j\�ome�&ueMT8��5�[��i��ŵgo�Eg%;��$�k��Q�T��]�'UK�{���&�sT7M��i_`x�	�cu�;+X�%�;/���( ����tDoTeL����ڃͪb�
��t�L��6r�bf� �"���^K֜���.6��&����t"O�$ϥ�f�p���kVb@�n��}��YjÖ}\�ݏ��0�*�� %���u���-�B�!6�&��}?;؍��fG`W􄸰���%"�tx�=z攮ň�nS�Jڔ�i�&����{ǧO5O^)� �ì�@eGX1����J��۝�p��i���Dw����7V��"��ܭ=��|���ށ~�+P[�̚>w�aH�#(�f-�sE�sEm@^����J�YN�L����|%�����[�8��\2wV�� VK�QB�f�8x<v (�Tq��vHd��K{G2B����c�\\�?��=#cB�I� pC,��g�<�a�D��u�8�����G=i�NǓS���`��ێ��t3)ޡg�m�͢����}�Ȏ��O���#2H6{#�9B�G�O'�O��3���@O���j_�Y*��1���	�[�<_Js����Fʉ�F�s�u����N��@�&yı�3����id��;������D�]뷇����v��e��!�T	��>B ��Y���9�M��zh��!ϡ�G�AY?L8��x�����[��>AFǚ�a�:�˛;��%��ļ��f���$�� y^uT@E��#oo�$2���χ!�P��A}f[�эg��Vo"H!w����
[��4M�m�AP��j��@���ƨ瀉홙�',.b�\��N�I�8|[Լ!�%|�Y:�6�[�p�����:�=��~����-�q8B۰�XJ;��1�S��{;�;��PEB�(�.85��7P��L�n��i"u�� te;:7�dz#)<6=�82^�
�F�Z�vf�������ǓϿq��4�E��};ώ�����S���u��� @�@�����}Qt�R!�?�*������P[BF�'��7����À��z�R��.<��.��C���x�J�<�Z~a��? t�L8b4^AEe�d����9���e޼�?$�Bw3u�J�-�c�wUx��蟙)���gt©���P�ד~����{�ڐ2y����|l�����g�Sc�VUzr!�yY���z���k����)NiK�u,��?�����>q��H&R��U����7a�fB��ob��D`A� j�8	�N�/��&�n�����ī|�}͈��� u�8m���$�/���?���ΐ���v�,�fP0�����8�X������y}��)�ԪCT^�>������/�V/҄����;)4�3Lo7�'�,<�=Q�R�� �=kL�I�H���B!(Y�A����~��)I�����X~����80?lKt�U=�v==�g<���J}J0]B��LۭY7���e�p������{��x5�)8��X?��4sg���xz�}:3�'��ef�R3=�Ӄ�S�Z��0�����ݟ���uQ=��|oD����c(�'�cԭw���D��r�����ic
���5�Q�R��ıj���z�6��r�ta2�nB(�ے✝�j&R�'�AN�I*� YI���T���.�+N?\���Yo�cq˱�b#A�����m��4qݏi�/M��x�u���o^����ba v�Y#0/���h*�"�2Z��e��s(F<t[~��ɚ�e��Wx9{��|b��y�/�.C�߸=SJO>�s��lob������Z��w�5V*DͰ����"���s�b�X�nz�Ѝ͡��_�!�!@���&�5��9��y"ٳ%������_��ɴ@�FT]���"Ԩb�_���l�����*�
r�rew����ەH]$ň��*������: g���pC��a�`Q���9s���4��&�\t�����;�Љ�:J��61��� ��k��Dj���
tq�0I����v�v��K�-���8������w(5_��291����F}e���˟���V�te�|'�{$���K�G0�N ��¢=1�X�/�:vW=��=K'.�L��K��*�ǃ˂�R��<f��Hq��֋.eY	p���Sl�[$\��y������h$Y���3�e4��t�˃�� VT�q;I!�/ry%��|Ĝc�k� �zSX\ki�����d��Z�?u?������+r�b幀~���4k�3f���>fRqUiZ�!�IW��xJ�d��6�mG��s�au*�h�Ԏ;�z��ԫ�ގ>p%MY�;��+�=#C����~H��ߠ�~unE���y�ؐY,��(F�����Q����OQ��y�E
�x��aU��G1M�n3�*�]t�]W��2N����\�3y��M�>\��.�ne?������T�,���G���I����%	d*�9n�d	c�)�{L��i��W����	�����`��~nD�A`_��>� �\F����������տ�0��M��n-j�U�H̐N��q�~(�D�q��|�,b�˧�A�t�Ne7I���':����)�~dD�K���9���^	�?b��M�<��p��ȇ4-��-q>h��`k��X�Ω��h�ᘩ:�ؐ^3I �A���o}e��0d:ۧ�e� �<02��9�5����B��dx��5:?����M���h�<3m��şT4���Sʓ���'Pq���ƹ�&I����3�O��34O���לm��0 j�B�����K���(g솕
eK t:_S��够)�3�^��G��e�L9p--��R��Ř�B�TY�v��iZݤ�VDWj7��TVC!��N��y��q�V0}O�j�t���������
"��5�J�v���fn�)��P�	�C�S�L��"�W��wU����c�㿆)����.a�C�m��%���<�z�_��r�ڗ�tZr߂,
�#�L�aJdx[���[��J�+	lG��M����Q�o����.K*d-}�P�{�0��Z�7q���S��#^[��!��~]���X�݀�����O+�B:�Յ.�+uXe�ulZ�`���+����n,���m��[���G��1Wtrd��Vw2�}� l9:��t�ZPe��x�_�J���Y=ќZ���ǭ^�z��q���.���p]�)M�&T�&��ip�?s������c�����2��)�Z���{�X�H��S��G��:N,��̋�({N��ӓ��U��A��Z`�C���JR��s��PrA4�"�����@�Z<��,�?��k�P�c�<��f�%'��%��;�OS����OZJ�3��L���}k��v��ж5�_�ؙ���-�H�?����bE}�<�a'a���vB��`�͊
@�����a����kJI �{HZ�'�~��4H;��q���X��_/F�S�%�g���j�hH8��5�0ʃ������b�3�^<��B=�C,�EG�5�׿���3���s;tE��(����wD��A}W�1χ�}@t����d�#�>��ԍszc&�nY%!�{��� )�Y_��-�$b7�PB!���Ğ������[H(����_Oh����l��:�]r[�ci��:ڊO1*u���M](��c��8݊�zBi��~r�<��Q|{n��V�3�VQ�~!�&�o�d�^j-d���j������
 �2�8���i��VU̫J�&�=k���UT��ތu����[�y��~�X"'i�YPx8�}@��{7��S�Dl�?�g�����׫����W\ڕ ^����@�8L�=ۦeX���km�����UN�Hp:���>	!�c�b�{B;��GD�"��۠�[5�V�Vv�T�%.-P�x�O��(�y;�l�4�ks���ѰIG|#�<-_](��g/������7�?D!:�/LD������E�����,�V��s�lw�hc�6Cξ�|���`���F�ucm;���Ȝ���q����}mr~~G_5�Tĸs�.uw�������5w��3I�	��[_P�>o!6
;cgV�&��YoQ�yU@&�������$+E��?x�G]�<�w�ۻ�$L�q��ny�M���<�^W�luK��_M�ѹ�,�������:`w�W,Q�E]�S[��f~)��&:����ד����?���<�7�1������`�i�fo��X
4&'�`Se���S����^���Ze��(w��Nȑ�3��FD]�}����ψs��ұ0�S&5�����
�lL���/r0��K{0H	�=�����
��T(�\`�Y\a��7����EHÀ��튝X<t��<�؋*y���Ч�����<�Q���ÿ2ax�Sh�#@t�x��:�����.޲8�f�U���&]�5��@�M	���U+f<���*�
$e'�m���n�Tŏ����'��Q����zȵ���*�	�&��by����0:��9?�wQ���lK�ZJ���(/���XN��.~��s���b�P	���VZ�@m:f  ��7��A�	�~Qk�ܫ�G�rFk�P��UB
J�J�A{�Sq`ԙۄ��*��Zyw���~�ei��l:�@�ٮ�A�:�3�@��"牞���6?2"�l�j���S���_S:�werؕ�f�D{�\�L��Z�a9��5��Z����%8��J�*� ��\h �w����,�ǰ&���{�}QO���dN�h[d�C{[CUg�')�������<�b��`�V��Btv~����$rlt�����[w��"�W�^E�I=�bD��Q"�����B���ǽ����Ű޴Kc���VH��6����ɺ_��G�T(HM���YU�*ĴUM��)M�7�PDBign�}�]w����՜�LC7'�u%_���s�~���9��*i��'ss��������B�eή������JR�+��n/�����$6��{�T$���\p��o&��U�E7�v���4`,�����؞�����R�=�H�a�<�̏��  ��wU{�ǎ���c%X��B�/{������#XZ��LK	�������͆9Zt�v���[f�����鲇M����ݡB+��DԊO��=��7��R���@��c��U�\c4tKu�8�oy�o��7~?��*���[c��jC�j�����s�$/e�`��R?�B�7A�#W�\��`��%ar�fn��3x2�Z�R�d����3����S�w�5̇I�d������'zՍ�پ��r�M������8!Pp��S�?k3�εG享�μ�$�:1�T��������T����]\���$lQ\��*��2��Fo�$�՞��Qr�m5Iˎ[#���G�Q�2����1�n�R�{�l(	��^	�?i꒓䳃�V^�ګ#?~ت�k	�#�m�����n�\H�O5b6�Ƚ��e�q/��\4�~����_�Z;�t���~Y���)�inG�)4�k89�0EH
\]����"��;
�/�E���>�ꏎlV�p���ާ+�|��*-7��鞽iu0�p��:���,L4wu���*�ތ/�q~����%�B�;`���d���^E:H}^@`3j��K��q�m��YJ`���z@��"X��ڣW��x)�TQ�e�=��s�8����O���3�����9�X~B���X�P
47L��%���!�&�f�����x�Ȣ���Z���! 2�\�-V���鷪�y(<I@��^C��g�;O�˷û]<��:Mٳc�c2h;q2�d
V-F� �lK4�N��8S[�q���ã�R�,����v�����^�w�w|'�y'1�����+C�A9:OC��e�V5V�JzIV�<ƥ��NJr���E����4n�H��?�R���"
nE���6�$6�
�ji�x����sQi��:��̠�ׂ xJh�}��.��%������"���fˎ�`W�K���v9�����H���v�A��;aL���N�Y&�`&�u@X���nH��5ȄH_e*O�3�?iW@�|`7q-ͫ����2�P�N>1�9y���(B��?�b��Uw����<[�K%%�d31.�&�}�
�;���<���'��������6j�`��@yo��y*�<2^��В�l�G�>N�Y7*Q�����������"8��!� �ݐ���n�or�
��}<��H�W^�շ�*���&�����%��,X�j���0b�*짱��F�5c������,���ʭu�<��Sg^���f�(� X)���p ��jr`����?�$4*MW]����-x�%H�
�5LW�O�2�a|D�,i�[����\�EjB�����]4`�������[��bW��a�-��o",9��R^�͞������]/�δ�d���4��e���!�WbBIk���)ɿ�v�[_�=�߭Y��� �)8��/�j����A�-]��o9�J�7A膰�/��3��9�N$Q�[�j�|{T!��g��t���$��O9��[�ׂ�ű��?��xزO�PD��\�.xn[��V6��9�R>w&�`^A���+�)��y��r3k��w�SE��Lp9[�*�������(F�ivĎ�Xp�<�vR�!T�#���cMԒƳ_q��A��A��dMFS��Ot��0i��B@�/L�Ev����)�@��X�W�<�QqX���Ƀ�s��S��B:��-��n�$�[�	������î�B�l@�|��˶/�&���Dˢ�"lb�E+�?UK;�i����s�X��'��oi��f���F�E���0�=a������� ӕ��+a��1UGѡ؝�H�C|L;��3�(c�30f,0M�WP�f^�t�q_��$�i�iЬ�B�& ����lP�w[)��~�wlz~������Ep��2V��x�G�k�L�h�m�y�kپv-�yQ]'��D���������ٿ�nu�yлn9�-�|�r�f<Hkh�o�O��=m��tO6�� tg�]p|Y�X���S�����ٛ�Z4�0�9�*���!ɗȥ0�c�H]����'����-Y_iڻ��呅MD-�ZA/-[f�04���~e�1q�P��oG{J�X5Y�w73���;.�N}�QE_��|n�L/j7'��ұD5������ZW������1ԾLPo�<#?�����hUҜNe}.�\3�`�?Λ�F�T��Rg���h�W:?&Z�"�c�CG��h�m"c 8���3������uڪ.R���}�9bp%�7s̝ŕcFI�4��.Jd��|!��L��y\N�M��z,T��a��\|��Sяs(a4c!��O��Ԉ���-�P)����K�&�{)9>�"/��k�Ȉtng":���/^#����Jx��h���&L!��9f���Mi�+?Zӿ�=�Pj��Q�$j�7��`��~𸀡�%�j?�b�Ö�/��~M��l1�'k�HgG¨�j��3��"}6����痘 ��D���R5ws_�clpll^SJ��Jէ��%����PHz��u��Z�J�H�/^-�:��2giH��z�c<OZ� �<n!1X
Z�_��J�T�*	�w���^�L*Zh^C��_�'4�fW;j����Ia�>��s�[
O'y����v����c�X�6����y��b�WS��i?��-!-ٗ�M�Nt���=�j���l`~7!���xݺ�u��&EW�P|Lb���R��S�4������ap�"�*�������� =;�j87�g���A������JI���μ&�9'�^l![z��X���!i~L���4.�d�mH��]T�U�7S���0�VU���4�oMJ��P?�BT�z��^Y-�G��n���mM�����*�XO	������K[����|�^���+��1�k@@d�d���n��afR�)�{�7SM�@�wL!��hP���M��g�֓�n�N�3��_�1�W���a{S�pt�� VR���#�9�>b*��>.y5�?n� �@6������Qx,Zt<A�J���A�
���W|�5��2el�?�E/C�=-nLз��b'��D|�G���|7ʑ���R�3�v���$
�v%�Y|�_<����m�6|;|�мs��sQU���O�C��3NJqsu�b�c�:�ZJ����?E���w�|��ha��4�ȟ�{�W�����B@A��.ȶ�>��N�Ӟ>e=vXnʈ$�Y�+�����i��v�@�M�h����e{L4�*E��$�D^f��*,n~����1���$o	B`�9����Шkm�R5�����f�������Ԧ��O*����

,�k����*�Ut��_���N>N.����*���@QY�[(@����"Z=����}��X���#G�����m!�l�
��}9�h�V�ED��S
���	}XIƩ98�;|h>��E��Gk�L2��-��[dxԋS�ޯ)W�k9_Py��W���u�1� ���⳿-Mo�.m�߇�e��t�!��Ao���.㮯�g<[A� �p�9�5$���A|Q�شĂ�L+�͡nz���~'�@��ɼ���a���Z��|�2�����G�2���"Rѐ�b�\�3��#P���f[�X^�u�����<���F&&�~���C��� �*47�xE���Όh�Οb#��ss�D�0�a���5��-`ß��D.u	�Җz��f���/���/�P���'m_�z{;�ތ��D�a�H���l����yg(pן��������b��x��m��,ęX��0˕;&��.�g���_���\ёD.�*�=���'���V�)l/�+=��ӗ�����4��mJ�<���_]��[$�>�?G������?�q�x+��Vj����2��a,�/��A�G����9l�/��4����}�l�Q��3�J�l]��̽�`�4z�c}+���* ��<�<�
v`Ĳ�c{�b��L��é4��T��ѡl�ҥ\�_��y���r�	-�6Zf;aj��B�ɕn��lm�H�pA���@���Bֲ�b�c4�;#�ѴT:΀*c�o�[�\UPl�������EPz�$+��G��E�2���<��y�:��*���q�M��T0f};A�u ��\��5j s��>���M��=m�1�c�Y���xR'�����0E��3?���7%��e�V��v܁Q������3W�P��x�5�r�J3 ��q�*>�K�=1q�d���M�� @݅����9�[>_��g�*^A������}6ċ1��
��tP�H�b��O�C�Ek;��p�XX��Ⴖ��PQa�"��v����}�ά�ō`,����KNZ[�
�}h��5�$�免�U&#�?8EU��?�d� 2ls1h�n���u�.��~�K��)��+�g7kQM�ӯN�[����K@�0&�0)ui.��;HCn�N����QK��߄g�/��*R8U���Z�R ��u���6��,r�� hN�h�I�S�v��b�k��'�?*oǜ��aO���̭/f3��G_��=�m>!��Yof��'�%��t��x{0�_l���S�:��'��k%GSXG,��1�6�h7gL��ݸ�3�g�8ӻ���gWpb��b� �����h���k��o� ��&�LA�vy+��#�V7��3������������3Fϛ���P�W}�r��'`�8~46��[��ƪ)<"�cu�ps��)3��L}�p�ݮ��'2��$Y_ě^�*�������i�u�1e�� �D�=��x�y��Mui�������Q���r�D���6�l�R����m@~l�qwG�&mo����1�V������L�i1/cC@o�CI��V�ӈE�v�"�������	G�������Ƽ���Qt渜J��ΗPc�����ɛ���,���σ_`�*�#�E�[5�. ��ƣ2����l�Y�sM �U�E8�R�V��)��|��2{dh�n�)Nr�W��.@C�D�>|��xm�\C�7���rz���.��O]��M�rp�+�H�-5xjK nd��h���<k$Y`x����XP,1|�%��c��k�����3�S��?��8`�5�Z1�F"�ve��� ��r��pF��;뢐���;	=�#�ƅh�c�r9"4�J?v�������Fߥzo��$�F�o:j�u�#������Acű4I�r����	�:�>�vU�v���P���=_�t�O/�ޕS|Ff�G��ϟ]�g�L.��b�{M��6O`9Ɗ�u�)���@������0m/�̀�<��g�]��0�;z���P�Q�:���(��8�X���!<�"=IXպ�$�R���B������X�v��`O�..�!م��+p�h^�S��(��u������_�c`t3�7S_�����/��Bd5�\��f"Zh���Oe