��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jåا{�\�u�?߷�dn@6�zf��r������;��r)]��<��ih���p����*���U�t��c�Ύ�M��E7�f´���@wֶ��Ɖ���f��b}ί����Ŝ{�s��(�WFr��̘���9c���?˨�@�:^P��*�
��Jn!W����$��,u�B�7!LN�rQ�(D�-��"xP�-��]���3%�׈Q����;1�DSd���ߧ�6�),j��;���0+>I -P6,��hj�&�A�z���J[���4�$?�����By/b�
���Ш��ۃ-���=i+9<q�����Q�73�����x���=����څ!V���T�}^��`ĎFp(�H�U;����rR�M���=t[�Ą˿��w3pZ���l�l �%�y��ChH;�.�I��./�=����Y����=�X��>
@.`,�#��~�+o0q���\���6�b��t+���c���ܯk���K��d(�X��)\^©u!��gbM9�3qR`�LJZj�7Ds���f�K^�":�����Z�:���"�/j���`�����aɞW��{���C�]Z|��>j]"%W��(�'kY�?mn=�}-:�:t_ �������ם	�7N�O��vu��l9.�nuv�]L8�.�����踸��W.i(:�~�;	B7�O�9T)H^����oC����1M�o|�B�9��}ds�<�������[,�´A~R���|4 �9q �"��,w1���e4���YƤ�6��\QWN���n/D�q89�"Z]�7>�<��F)3=㙞)��`or��۞�ye&��
�(t���b��Vl��i,��ud�l0A�$H��3��Mq�]�~�Gs!g���|I,q����^���[+����G� �S����őX�s��W�M��|!њq`���sC»YX|�F��X.�JN�cN:^M F�3&��4�A�BzHА��]��M�y~6Ra��f��J��Z -Y�P8q�燴$ޱ�&�mya�<��f�Z��>���g�hI�2��+MY��~���Q�Q��6 �m�f
�P�	q6���N����`�O㫁qJ#w������ˈ?L�L�#��	�J��I8�d�VC��'�Cv��T�FB���HM�фr�;��K�,Lkl��*����F0�A���ɖ�l0�7��(��oL����)5�X�a6s�e��z�MLv�y�o���.��p�Ml��\���Y�Zxյ2\�X���v���P5PD����jW�)X7���%���4��vY$_}�f�uL�~�/��"��5�0��F�U	"\�̡YK��I����d�[�ZP����uߴ�V%�ǘ!oP,�CzC���~u�~���F*!��lP&�L�åF�׮}�a�_:�C�P}��Vx>�
��>��2�'�A?�t�Ʋ ���������:�/&�^�<��j���w+�:���@��^#�<P�ن��~6q����nて"����\M�� ��3�����a�;�k5� �C"��qߔa�㪺:��Z����Mu`�1��s�m<�;����꩷���[��K���Cx��c�����^�t
b�"Z�]�׀*��(����nr�%�Z�bYrQ	V����j#vX�!�ä�@����̭A��"�o�VWq���P����e|#0�[�"%Mz���f��"3e?�N	�<� ,���\v�gUW�e��{M���u�����gk��(�pQ1�����u�]�L�ui[r�;Ss��m:M�3A��Pֵ�SPA1Ô
�g�B�æ4�q��TG*N�2��d@(��=պ�J���j�����ޗXC>�~�H�pPSǕK�?���ߖ S�c�|�����9�Ir��A�lS�Y��	�rD!�o<�<��(���
��Kd�hE���|�_�`ئ��c�Wc~SP�W���GR�Ϻc�0�����t~4I��CA�-u� w��7�
����C
%:��؟5X�3�أ '!VF������7@�g2)?�z�_���Bme���|�3�[H|!2gϰ���<<�4�j���]tՈ-�	Q����Yz���������+S��}9�S��r
F�+��>�A�u�`wv��E
���f�KF�T��xuEs���[��� ;�B0��B7�=�9FI-��oU���%�m��##)ѿ⠘���M���L�
@4a�,G��$bI��õZ2(���(<tùS	>���g��\"�<X��\�sW��M��KW"h��o���B�c����G��Q�v��_��1��w\��k����x��C��3�ߟ��R�(G@���X6#�ڽ�{ÈJ\��e�Ƌz��J?�v��}LQ�G4�:���"���?���_54ER!����	V��9BV�Z�=U\��{ڟ�/)�kI*��_94���`7(+;���d����X�T?/&eFU��QW�iB�0R��R��r6�HAx��^�8���ͽ��g"�YWk�9�Bg[\�Yx	�uʔL�8 C�����H�c���b����!4AF��E�%��:�PN��������Ëޮ�V:�?�A��;�]�=\�v��=	�?\�u���e�yGC5%pG��
��ҴF�4^^�<߲~28-_�PH�^g�)��C��c�P"��2�AQ�!���0&+3}��
~#�j�I����H~o"�j��"���-ꋇ��Pԫ5�f��[,��Υ���"���w|�xiH��z�Y'� @��?dV28�J��	�������?:�\KGqf>e\A!y �K!���^7Qa�1!�);N�n���o¿v�0t��a�9��`%Q@l�{_�������mj|*`Uf����xf�`o�t�֎[ �ڋ�4KNjp^����Ս<����*���F���M =cU9�0����p�"�|���˷���rI~*�D��SR�otՃ#A�Ѹ:�20r�3a����}���;g���8��b�<��!,����
w�J�I-q�"Wn��[��]���X
�ʈg���4�4���m�Fϵ�^B�Q�R7���^k������֯�����"�Z�a�|�k̤�)k�X!�Cn��ӵC�U����d]�c2n�r"@d�D�Ӝm6����?�h!��*G�Jy2K�
�_�Ub�,��5Qb�&�-lö����t&}S������'@�9:���!��6y-p8��:u.Ǹ�3w'���jD���|�V�L1��W�	`c�Ͽ�Ni=]���x<��KT!�|��9><�b��m1*��}��G���j:�l[ޣW?V�[yt}^����r���L�������W�ϧ�E�eƊ"F���a���3V��НW� ΄�f� �Z���u���(=o��6|Ὕibx��
��q�)i���Hߚ� �դ������޻p�Z��˄�#���,�q9��� �r�ʚ�V-�p�ytq��C1����ӑ�Ub�%͜�K/ED�ц��ȑ4, �q�������9�js�������(�G6{�Sr��
	��W�p�b,�ۡ9��J�2�0]�FG9����~�q���T��q��.��+R�F��l���`��Q�$[�B�Lj��ќ�<��ٽ��u�iS��r�J`['(y!�^��oț��'�@��?�s��݅i���7���V<
��!ܫ#�}L���)���);��+%�>q�N��*��;͕��NP��PF����tMn��3;y ǵz	�����B
&�^Xmp��k� F2�es=����&5^���`皛���h�����	K:���*��F�x�����/״�5�qҸ�"�s:��s+ 9)�Iq��"[���5��la}ػֆ���j�^���m��D)C\��Pev-�Dqخ�����6��Z�]/Ǡ��>�_D@3�ty�XM,��T&?�2Ʉ��v��*��h�`Zr��N	��
��Z�;5�H�"�Y���|=ud�Ʉ��ig�p+�B.�V8F�y/e���h����gY��S����a ��������MS��E��!��7�V�n[��jK[ fܛW�	l ��}1�$Z�Y�U�xpFԏ����C3��7�~�>���lh�z��2X6*ĪG�S\v���d7}n�]Q������"
�㖢�
��ꩄ`�1P�����E�.l1���� w��e�٤oθ��i�u�	m��#!.�bx�_��KT.,w�v���$
@Ϧ�5.�*MD��dS�`+E�[g���ο[?11�wf�ؤ�Zl7�g-�v]�EŤ��eXυ��7�z��瓫���]6,/d�����4WL������?p5`C���	���LG�[D?в?�[�Y�u�ه8�5>���w�ь�W����S��2�1́�"�?tDva��Bgs��n�g��g�Q��q(�/�����c!�$������@�?���xD��,	j�>_��x1�f�:�Y��RJ��4}�O�֒��sm7��P �h��c���#Z��v@� G�kL��nT�0X���o�dG~�Dtu�X�MDlv5��י�i��� ���p��y��\�7y�M��6� �$�R6 8�7d��︯��cW�O��S_w6Yz����2A �����b�ǂ%�e,_C�0���q8h���k���k ���E��ˍ�㎥�N���]�ȧ�yO9�e�Ew���� �W�_1�FV�|^��zF��H��7�,�ص,�'&��pw �yl�%'hﮝj+���j�����}v��s�>�_Q'M���w��� ������Pp�0���蝯��ks������<�е3�~G��c�Gam����粣G��C���$�2��T�*0O�ihq�0��gjL��n���W�8 � �f���ZZ(V?�`G�ę�n!8�@�	T'�N�&�	\�t� q��s��TlX-�X���R���*��	�~��YV��p��v��i8A�-�)`�55A�������7x��zM�����{�T�J�NRVTu�+g5��r�@k�l�N�S�۟w����� 8�iK\ ��I6N6	���)�*ޮ��߷7��A>�ߩ۰,���;�j�⪳&��	�"i�q�C�/l�<k����7�Fg�>��	�Ͳ#$P��h�q�R���&�H��;ɃA{н`^:wA��[V�����{�A�+��a�9<�xj�w ?�]o��i_���"g-�e���~�98�G�D{���&�Џ*��_�:m�����r�芒��Q��������U���J K?��ʨ�� ��֒����E�ok�Ha�D?��#I����{��=n���[<�t� ��u�Jԇs���+�y�9%3�(�f�ش|t����1�n�|o�>z��y�)7i���>��㷠��u�h+ASr�p����,�>�w�_>` n��}}�'�ڡ�^����<9oC�s)��&�g���M�cA»��`��2Y`�$Օ�B�P�t@N�m�?Y>r((-���][!:P7�j�o:e���y��	{ 6/�eh9�����׆������on���8�t���g�:�V���J �����<������H�.�*�xV�i��8��{E��!�ރT�yb^߹�˝F���m���	��^!r��U�1��z�\r�5����b(L��A�����7*<���f�5Q�4�ޠ1JV�ޢ��_�N�Ōbʍ>̄熤��N@�|7YG��@A��ioJ�[?�=f�9K�#�}��JA��)�(w��Q���-k]2�=�5����
�����\oq�������í?E>�OH����(D�f�>��`i;M������?��� �i:�`e
ŽD�u�x����d�sթ-W�ֳ�����$?\B4A���#����~�W�m=�&�1��}��#<ua/y΂��͘����%�󲤞�x�7'�xZ�>_�Uh��@�����X-�«i�"��%@�y���_��i)!�1�9��i�]8rY�k���:��ф%JMbZ�tu�E��&VER[�H��+�<*ml�UϹ|]@T�`�ȱ��z�7I���} �˔�)P�wL�]	������捗Ùk�=�\���
�p�$�� �n7��y�E��^A��𞶘D5��L��k���x�_�6����͒�f�ܛ��㕰7��	��*-��n�|�z���.�%f^z�﩮��l�~�Gվ=��% ��^��M��)1 �f�WK�#��a��Fr s�"��5��x�f|�(�d^EMY�^h��ֶ�nƃ�����I7�Na8@sH��㞉�~F
p����J3�'�z$��
�Wkb_1>��i÷Bl���b��/�$�����l��ltyH�����0��h��+p�-�6�p=W�x�0)�Í{G 1�� �o��	����0���՘郺9a<F��ZMhw��lv�`%L���|�����Y�y����9sq���8�f�\H�z�/b;4�K���9�_�$��%В�����f���}�8�'����Ύ`b���RP�V��Lq���Ƒ�&;��u1k-�pWӗ@֣^���t��v��Q�A�U��p;���%�W<�&�Um�*f�[��Ӌ��qkޛ����D���r]���>,�gZA��a̷В@�j�e<��:�v��zd |���!�ut�ψg�	db�V_�Z"*._�1���?�u=�W%�pմB6��MB.ºI2p0�<C�H&� �\,����_E�F�(�8��b��IZ|���Xi 'T�����^�B�ތ�%�3���(�8]&7w��A�6�|>�Y}K��Yw'a\ɐ�3�7��F���"�6��x��_9P�9�	��	_��w[��8$����]�����E^}<d�c�������!:�eF�z���z�x���x���a3y��vȸ�}8�񀨄�Ռnڇ��N#���<���h��d������ g-�~�]?��۞w�T��< �PR�����&��<���x��g˲���eA�ܢ����_�4b%�X,P������hB��ޭ��^�c��(\;����T�W�u)���H̟b/S9���+��	T��G�m�e�׶�>����1I�l2�뺕#��Ծ��l��vc�Q����:�4��Ec��p�w��	���G_��LZF���N��-3��W1��|�X��ؐA}x�ot���d7���-� 0^`ͷ*�r�[Q�}����H�����⤉TC	E �̡f"A\:{^����3cjj���?~_U���P(`�$�ax*qΦu���&> "�ό�8=�X����@C5g´���OQu���!x�.�.�G ���t�L���./�2���^LT4�{�b�%`�����Kb��D�*z�00��R�6݉C�X|:O�:�
P�_�~�P�A*�j�&d�&*J����
婥t,�t�?W�R1����{���K����<�CMR��E]����6m?^�m�&����l�r\��!$�-w��cH�r��?����q�M�- �Q&�m�J��H�>�h��+��r�,Z��ј�Tp�3�C��ἐ*���c�;(����5�\ߧ��_
Q��oو٧��:qD�!k������6�ݛˮJ�t�N9K",1 �8���9����0����+Ү�f
��B�[��������2�M��a��ߧ�Oq�(��X���~ꯗ�#_���^, �G*�~�}�]�`3���m���]0p��XVC�2�����7Z�h�v�2:X���;4�+�0�^`�VW����lr)N/A�J�5s�P��sy�����G��R:5\�+N�ӆsz���<�?N}'��@��C�Λ4V7Q@ƃe*9\��S�p��"�9}#7Xsx ��S03Ne^rcLҠ�e�K%~��U�7������?�k�~B���3]�&q�t��PNa'�}���1+��ʣ�-��I9��	8�J*��~뱓��i51&ɰT?�k�µ�^�WE��:n4e�+�&=7}�b�x��_��1�Y����{��ΰ�2����\��1q�����^��8����`�lԖW<\)�[��9 V�_@��b�nT˯�VG���h�O���	�/��j	E� �L�Ֆ�3��Ѧ�--�m������;���:�f�_һQ0ObLFP�X$�pJb���%�����i�8�j�GpA/J��J����=��m�MD^Z�3N4�Ҋ�̤T�2����Y�ҁS��e~�=�wR��|lg��*)?%��!�`hJw�*��J�@��\V����^�	�4)v��Q�N�G�]޷�n���
�w��P�u��4�z&�)J�pw4*?
�#_M��Q�z��Fc�A��$M/:��cռ��G�P���,C�A�ܟ�XX�]�����]��BN��?)lO/ !�
��|~��z�X}�_b7UBp��͈@�g��q��mL *�6�;�ʨ3�':��u;�5֊��|���J��;y��G�"`F�99+�}-Hț\��9��o��$|���)����K&�e���D��8�_�j��Hq�{���tNa���<�>/9Ψ �2�&�+��3�g<���.$x���)S'T��]����6��A\��C[2��G�PڲcF�I�G��R��� �N�c�����4A�?\�3ʜ��v��;�m�-��J$���<ۦh�5�"Ȉ�ZS�����eʻ<=�E�pG=$�@����S��W��<n��hxc��<J�	?A�2[(p��Y�f�9�W��֍)�A;��(�,�r�� �;�4Ps���)ZD>Pj}ϯ� !��*m��t֏���<f��u���ca;����\v��$�^ֹ+�D^:��`��3r����D��EDi��e�