��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� f
���O�Q��Y.#�d'���J�"����4���d�"�Ŝ9͜����
�~�a�rN�����o]y����1���nJ�]s 3L!��,���zَaw�{,���{�b�[;ҙ�u�\��������.7���}����H��ΰ�&���ے9��y��y����͍2��ё(��7q|U9��1���i��$>�[�G���^#fU����S�"_a[7B��7~ez�#�5��-������>[{Љ�v��G]��Ew4��5`�|x}��4�y�z�f�|#�դ�e��5p���1��L��d=�㺔��y���h����V���Q���t�̿�rբ��6�j�mcP�iT
���c�j��5�j�KL��tlV��d��x�Z��"ks�kCK�|�i(�;�����6��12�XTeP��[��'�0u ����r/X�<��/�]Gȥ���%N��]84����Uwp)
���un(c�Åf��J��f`9Fqv]���+�<�w �N��fѧ�h ˞�C;4��#�i��T6n�Q�T�����ڸ}�rS3�*�x�٨�j���y�~E�s�~+s�G��'��%`+�w+.}��(Jľ�$SL�2-�M�M�W5~���/%��t%���0;��3��G�rq�Ħ@];
!}ˬ � C_3ZjT5�ъ���29L��>ԡ��I�#iDn=*oB'R�؍����v��< 2<���oc�M Yx�R5��ܡ�����2=ړU��oLW9oq��4S�um줂f�X+��t)�a��� R��M�Ć8��,=���LIQ^�H	�	�Z�K�M�I�)
�8c45Y���[�*�]�ƭx�ZT��>�~�K�gFq���J����ù�s��5���W�'_�w�yn�]�Zf�(�o�[�%�̏�m��lAZ�ˁ�`�q�ܳlAhϳ��Χ2��L�Sf�`U�z>`��(����΢`��0=U���,��L�m1l'R�Q.��|��u8ª�טU�.~[藣��6q���+˃�1�(�mN~�r�D�lp�R�ّ�3��xIm>�͎�CB���,o"И�n	 AѵP�ަ�c���u�R/YU����F��Yk'�핾����Tv��^�)�c@�ǎa�Uf[sz-J�V{݄�!M���,��P��1��Wb���Ց@�����2U�	���^x�tJhOO���>�iR7����	���b^�/�7��T����T&��ф-T��~w�>�1���9���*����HI�r�e�E�����Q\�K;�*��2�	;j�)o���eW��/l
��%�kÖ�5O��[���EG�|͘F~ay�?��Z�޻Ƹ��y�l�FO���Vu
�<�W���Eȶa�a�i��m�?�b��+RP�Ն91��*�s�m(z�624]rC�?XB�D���T̐@#�IhG٫Ɔ�y�T���$c�)�έ}�w;�]���+���"GɳO�S��~�~3)�;Zl-g���:�v(d��y���R�d�Nbด5���'�D�%��qR���?g��e�Ns�c�̖~NJX2�R�6-���k���/i�%SmtvBi�5G��Udj��8�O#,�S�oC� �|�Hۄ�B�w��h����q���2s֘A��?���{�+�Q�O���w�֗9/-�Ǌ*�s=Wqt�hX�_h
�o/Q���ˇ`��'FE�*��[s�f�^��q����E_Ю�Kqď�,�\-U�
4z�n�¥1���8��J8qM�>|��u������L�%J�쇱2��ߛh����ϴ=t
:��>q������۰X�Bg=r�L�KHv�^=���JZ��_F�������m�s��^;���v�}�r`V���<�D��u�f<�-�����-��1��
�N����wx���T*PX2cx���2�A��p?�k'���쒔���:	�''۸~[���*��(��d/jŐ�D���w��@	�;�5*�>����q��欸	I�~ڼ���&�Q�9�e5ER��F��/ ���xF|�V��&g�2Л��=��C@-��ЮF�:Ά�η��B��(����H�-�bQs����FT�
�0��Q��[�xv�E�����L�����dn��#��tu8�j*�|��vNcd\@������CQ���o��Ih��R	�0�����؟���`�'Ӣ0�[�	لe�6�M��������D����ߠ�B��Bu�Uczq�'N�������D%�l�ccB�cǻ�v�&��@�;�,�;ZBO�Ѕ!(�ad�6
�*Pe�nKq�Ǟ����3����x��
��%BK��κ�`4	�l�H�!G�&�݋��3�KP� SĞ 1 �N�v�;=��G��>�4����ffPw2Z�l���A=vm���4�T��2��A'���i�c��V�Z�'3nt�󶳻�1�[R��y^�UsW��r�et�ǼL���+-� c�%��H����_��r��M_����&�@����6�>^���L�V���6�<0��%]�K!ܘU-�i ܁���] �d�gE���n�A��deG�o4����e$+��H��� k��@ 8��!����Qp��a�+�~J*n�㑛V(�7`u��z���/��.�;'���V�����S�*4PJ�6�2���j�`�i��܍9�]�D ;�=W����Ÿ���=K��M�\����:.�88�a�l%��dWP�%Dݎ�ǿ�m��^'�E��t|��)e���3[�4jI�
�^!o��fP�gg�9a�x*�F)�	ш�X�?�W��kE�5���z7��$pZ�Yt?��׆�a���*"͗GPPJj��t6�"�����WG�" Uzl?g�Ŭ��Hq�}��$dO(*~TQ����Ø�I��)9�=�y��F��i�v���?v�$�@��j&���똢W�W���� @=!O�ko�r�?S$*����#X�b�=����dk:�)�ϐtу�!!��ɘ�}D��;��͟(mo������b���C��,e�k�f�	�W/�#��B8�Íl�ӥ+[*����=�����iF���	3