��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ��nͳ�R[�ظ�_����Qq���G�]~��\�^�W.Z��ke��X�?�I\�zA@���Y"���a`MBl��$���X���/~%�cg��OU#,��;o�w�F�~�wy�0�Sa��qC�$�_됲��ݗ� ���D��.����v��C��k���<�$J��3��I
����<[�P�}&ʁ_m3�P{�
A���-X'�H4Eml�}-���i���[�f�c�:p�D��8}X($7F�!�C�ﭩz3�s��d�A!r��6��
ek��C��RH����T������C4�Z����G�+�	�y�`�[`?�QG�;^�S�r��s濈&�����*�flq����)kD�G,i;eLWy������?��ع���%������.�l.�(��uE�}�ˋX5qkw�JL{J�վs\FӔ���sM���YIM�s۳ƒB�A���uC{�֖6}�~.sܚ��'�q�U7s'XL�V��-��KЗF,<�:O���Q[������u"E6�i̳nx�M��p�d��N��%��C&�Q���O�N�Ď�T�S
��4,�ʪR�Y��]kYne:�L z�4�Ӎ"�e��'w`{��D+�Z�~g��N���R���t��l{e�����jK��v�e���*�HIo��fd�du�@_�uɻz �[~W.�L����GI�����
~�����i�^����xd�1���BbF��Z9) ��W�B`|�n�i�i��0f٪ ��7Wʍ�=Ү�!�T�`�p�8t��o����8��zT�u.�Ԙ)s�8p��{0a7
���q���;<u�͝^�!AC
M��{�2�w���E�2��ΣbV������;��'��PGZ&�����fQ̯�S��sR����"��nA/�4�EMsi�b�j��'��B��BS��Q�i�V? 6�������P�R��$�yG��rDM��2�����,�oS�+����ַs��{`Q��WP�G#�����6?�a3"X��Ԕa!��ύ�
��#�0�#|Dҫ����Uo�\��~N�;��ow���U���(�2��s�>��m��#��88�m��O��3N�Un$��wa4�k� ��<mCA�u=�s'�د��2���"k��R1�@��icgC�uB�a�x�\�u2aD�/Iz.�vǇ(�e7�ʑ��Ș�p�4*]�#D V�����v�����7f)	vRw��FSȶ���!k���P&6%��t����ì`ӛ8������*?�j��6��p��7���7�V	0�ˀ-���!�*�r6y�C&���thS��R�S��C��a�^rŊ?�0�-t����^L>"�$N�o���7�1'��Z���fɔ�c���<G��i�T_<�8Ժ�A��k������ن����x��i�Ⱥ��Q�����5�*&�֦>P��[�S��=Ă}�����ef�Ae�ݯQ��?�I���.D�?�xRQl���e���X &�W��b���`�>���F��nwkcg�O�"��%M;��cY؞����2D�r9H�*$�m�eS�� v*'��>��׭����M�9�?#4e�����P��N�A����'U�|�u�|��_�/�}��Ȃs='A��iD�bFs�?*`K��":�=��/Q�8/|�N�	�g�2�����㳼vJ�C +�Ȗ�G*��h.�]JT����[<�H�qJb�;��Ʋ�
'�	$ꋼB�^�;\4���X�L�|� ���pԺ�<o(������2D
6�2�+"T�Z��&�PS�h��c~�f�Ex���q�f�=A����\�\�n��̹��׍�<[Ʀ�Rxt��ӡM��6{�����lw.1����fl("�>�J��f}��S��k�x:����CC�0�R�6�)\�o �^�,��@`�P��"���\�I
p±	؛��-��,��٫ʉI��\br�����b����%=�q>9@D�xk���k�Q�J�V���R}���w/�J��u�����B#9�pf��/�7	���L�c�b���;\��!iRP@kX(���?��y��+F6��r"��}[r�ם=Q�C��x7	�&��~BA/�8Rր27�,l}xth+�pJ�*f����"�qP�H���6��6������3�h�EB-Yt�B�
z6l_��b(���u?ֳSQ�k��[h[�ɯ��q��4A��ڝ�Z��}������geh���s헹r�LYH]a�.�5�
%��E�7i��!h����Ȍx��z�R��#�b7�V�:/���/�����|�Kչk���Ӕ��"��.2��b����c.��ZF9��	�'n��i�4�΍0��v�v~�
��30��`{o�z0J����]�Fg�۷��#�q��=>a� ��
P�1��e=oB�2��8�KiG�1�37��Y4����$������Y&��h�#�).^�z_3���]�3�jz��|�5czlW
�at2�3N���V��m�PwI�0oҊ"���akF�<����T�ӈu�o�D'��?��"�����]���*vU%h}�J�L��j�7x�
aЮ6�8�,Z'�6KupI���(��w���n� ���=�X^�/��͇/� �D���X.��pM�`aGäԦ�X�����y�?[:���8��IKA��Zݪ6��(�J�͕�,*Օ	��GQ����d\2�C�Gȶ�43�u���2m��$���r��]��U�}�(�j1I*�l��*�w|��m��|D�Z�'�\��k��?�Pl
Zp���Ju_�q6^�!��Q�	�1ź��9��x&�K���c/c���u6}�;��z�YN�����s��N�b�lŲ��d�D��e�g݆͏"�R8�^�������@�c�G�L�&�
jJc+�}�m6��6u�41��)EpCa9�+��p� ��k���B��,��&fz�S�V�mh�����֮0�p������P�RϺ�z��9/A��-1i'!]�3�����pWxm-,u������
L�\���q}����8���g�(�h� ?+x�5�[�ISj�q;mD,B�ĥ�izR�Ͳ�C�y�=)q�U'8$@����w� �A*G?d��e�������:Ӡ�[
$�R�wO(~P�B��`�/��"F�$�����1h;�%���`��,�L��x�e���EՋ�B���\�z$�\Pv�1�ɪkb���P3$N]ͽ@*T�ͥj;^��=?-��}���_7�wl0���?t�oWB�c��:��{y,��M��]@�$C:NQT�(f��}��L��7F�w�XjW�LE>��Z��l�Fϐ�"�i!�`�{8PU��D؃�#Nv���ӭ#����K#�[�@*�t����T�#���~�Q��;�c�p%���@�fbdrslq`�
ªFg�A*�򘬾�0#��短��[GfF(��ӗ����x'0��,8-�D��|���fW��s���j��7P�U�䐥���!HI�
�X,bog�s}7��?���n�l63����|ms�@�y\���N�U��Fz�II��v����&�{HB��.P���E�Ư�>���#�:�n]�7�5txq����:?5�^?C��k�2��tN1L:f��a��?�:k�8��]��`�"g ���W��<�.J�ʆ0<'M��d2�tֳw�eR��|�����Ie@s��)�(� d�~ÅK�z�s�2�I����۰�j�8Q߳�jEX�o-���i-���YX�ꢣZ�2�`�hVu�������Z}E���ٟJ�2�V�j]�Gυ�Q��4i���p���C��vQbN֛���0@
��È��`���6`:�n���*Lf�>ݝ��-�f������Ѵ��k~n�M�=3��#I�k�}��B
��Yu�\���Qk��f��_�;��q�a}��"��g��H�"x�	��Z1�I���Y8L�Mmc�n���}�R���y̵>Җ�4�b��)=��f(MU����/����?���y[�U7?U;�|(⣷�l�lߙk�P�x���\XR�2�YE_Ew?��7�m
�Iq<=Zj��D�Zۣ��d��!i-��ώ�C�������j�����;��U�Rh\��[t�o�����on�A��4'�3&�-�~�<XV�[ʹ�`��q�שׂ��/Ys��%ˬ&�v鶗)���AĻو��E���
