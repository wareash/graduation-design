��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e����d���f{��@����S��>���4{��ת�AO�Q{����-��TZ�X���LZqu��	;��7�c��0���\:aN2ϡ)"��t�F��ڨUAu��$��5T��u,A�~M�El��CC:É�+R��k���j���,�)+��`|�|}����)��[cb���\ziT{��QE?ш0����ɳ�|�L8=�Z��
ly�õz�d?�Y�o� �h��`V�߼EE�&F4�{]W�!��D�4w��@���7C��C9ӃL����
<^�}�������ۋ�5���T]������V
f0@����B'�����v�<�V%Պ~N�j�ǈ��㵒q�_�hz���,�wF�F�4������Ϳ�g���'Ș�y��V�LL��=�#q�ufҾa<4��6Ef�~��vs�c�`91��X~�@/�
��)�8�0�J�q�7�Dw>� _�>YϙxX"hsĢg��OH7��T̍���x�4�UgЬU�6�n���͡�\�6X�}���.yS�d\z\XQ��Z��*jW�ĭ*���m������K��q���nh��g�����\�] �v�߻/��[+�ݤ���"���-k��T��kf*���-B	� g�tm����%TT:.�D�2E��^8p��Mޠ��勒���̮�3	��~����L[�u�CK ��$��.������\�D�N����qSč?�W�QB��H��Va�==0'gn�n��gX�"m��/h�Id.��h�:wo1:jب��V����+�=cߩ[	BB����xłt�[|�h{z[{�cvAȟ����^�h9�����(�k�b�z@��� 1 ��?H�,<�UvKV� �X�T��6�A!BeZ��l�% S�P���jSWwH�A��C��@*#��^��������P�d���<�2�u �\$�h*x�ow�1�0C�抦͊���B�%���1|*G-��aŷ;�gǚ��@����+	[���L�E��V�^q�G$t}��f�[���V�ӛ���4)춯}"��}M(g�]�K�����+C����gP&:�g �h���ͻy��u�X�\�G�e�?�]��˨ �rb����Tvpu�7ަ|xIUw�W�A��� I���jb�N]W��^/P��5^���_MQ��K�_�z!z�YMH�g�����z2�,�^1%�a]T2��� �}��i;�=�+�-`��p�Z�`�i��}#�ބ���gf�zj7v$C�-�YoE;\P�z�oQ��v#\D�.8�L����u��k&�G�:"�tk����T��k�����<��ܦ���W�ܬ������/�P���.a�Zj��d����������1{�m�Pi���\=�c�R���7�� �Jh[����;	V�4�B�3\�qM�,]ѣ|7�A���l�� �2��ya�z!O$̸��k˂��ٮasp�P�81B��Bh�0�|�LvC���O�v�|��
7$����]R��� |>|���N��υ�\����he���A#ܚ8��v���OI�ƪ�\*L�E)?ל�r�:b�"�%��>7�W���I ��K�xsa|P��_q�-dO'_��Q|y����3sy��J5���8��cm��m!9
��`�:&C��#C�\�%я�����ޫ|��b�!@!<��H�%������"�k|_i�A^�r��-h��Hx��U=.K.��/EQB���.Y�K�8�]��R��b}&]�J����i�s/q׵�����d��=���T��}���<N^��<�WO�&���P�4�~��Я���u����]�C�S�Z~<�F����S��6�U��Zvq�57�B��@��C@��ݑ<��lm���ξR6ЦG݌_6��B�5A}Ok�ݲ�m�*�vL{}�������A�m/�[�+�����_� ʔe��oE���i�xx� �Ҡ��1]��z����ֲ����=�+c̫l��=����K!*qM�h�!cp9��\����}���]	vPæ���:���� 4�u���P���T2���4y���1��xz^Q&�<w�]�����>��p�\��ԩu��C��ޥ!@z�<� �ȗj`�(Alt�"��rkv�El�wU(*thVXtV�#�H�W��v���i� u���z�Z�Ij)RP!�i��*|	�J8�1+�K(���mEܥOT�DW��M
ɬ$�d�%o]̄�v% g�h>�����y���Ƿ~d2�oR#wQԬC=E~By�����A���+�'�
I:��3�G�.jHٕ(�wz;V�L?�:��;��
v�ݢ�=81�矌+ڢ��l��%�.Ժ�j�i���z<�0��Zm(ɽ�0|O��7�)"2�Q�D��������"�|\2�
���zL Z�Q��{�M�G�����,9!+d��cf��h����+�D���i~@W&�O�W:L��U��!Eg����B>�����h�[����ן1�o����΍�m�R8췾��(��B!1�f0�z-׬����cڟ�9m��(�`t�ζ�"j�6�o���*�P���s�l&`���Qc Ō�6�Y9\���Y��A` f����<\��Qp�����閠˓Z���!�3{B�
��`e��74�pjj;sH�e�U\|��3U�e�!�)��	�Gzρ�;i�c�+y �v�F��*#�r�����w�3��D�4�$y�����(����Y����e�4�y�k=wy�T��kZ���Ud��eog�Թ"#!c��Ib�,SZ�,��pg�z�t*���F��d'�
֚NS��g�-9E.�����,���n0=�Q<8Pk&�sQa�<W�U���	��X��9�K��E�Z��㣄e��b�g�\���z,6@[\�n�Ǥנ�����/�Z麁�<.��?�����o�B g�M��Ĥ��*
��J�a��9,Ų����U��wkU5��!5����=��|@>��X�?i�,Ʉ7F�A�܊��q{m��"������o��������