��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf\�|Vv �|�
�����W+i\�d����;o�o�[��e@[ġ�%�#`�G6D��v.s2s�
���Ϗ����1����ŰOy���f�˜��G\�'N��)�b��؇�>�j:�~��@W�/����*����)��T�vw�,��)¶��s�;)2�"��v����v/���1�qX�T���.��!��Y+��.:1&~x�:Dy����mƹ��Mz��1�V���B��n���t�l��q�����\2���=._c"Dك�X��?��N�7X!wI�e��^�-02�<T�۟ۨF�Uucn�{�KNe�x5�!���\UŢ%�hk�G�|�D`�� �%O(���]����Sq�h���1�	YR�Pt�ґ�?~)���'!QkW¾�z(�4xY���t�.T����r�G�G�qC�3���<�;_���Ah�3|���@�lG�ʎhf�J��g�3R�(���Nu� ����8�ږ�*z��+����pjw�׺��f�(@��Y	��=��I	V(�Óh�2�JKeB���.�&%
�Ѱ窮ɗ�vg��x�����֛�հ�`��h��&L���^�b�A-�����xh#�3R_����F��G�ݭ�fS�	�(j�`����?�M�2�;�<'~��Sn��*L�,@g��o��T���^^IE�v0�T��!4.�פ��盞�`��X: T�> e���4�vꩌ1
�����,چ���siO��M�΀"�q(������\}O �( �22����r�#��M�Bf"
W�"6Z�Z�wC���-u�+������;#����?H���~҄uW����Ɨ�a�[+v@��E�?�>b�xA��������\�=x�����NF<Eb�ڕ��c)n�v�5�����a��%���P�x&�M�P��(�r��Q����u5���_���+��@���r���ꗤ���¾>0�!i
lZ���{KQpP���nXF�rx=�=��m���K>����r-���-�h��˴�N���$��/�1��iEe���2��I#�SM��3����W���0k�� Ҙ_���������aØ؆	ct\�z�'@��Pc�'�ӧ�T�1���z����t�C���cbyM.'��o�����W�o�N�OA,V�[��v4���������.����F9Ce6��d�_�Y���w���\!�O4?��h-4s¡��?W�PY�c����e��#�0���5U��y`�K��D�r� ,���I�	����bs�����6�\�+����X���Sĸ�,�^s"�Y=�AT1G'��L�Xح���r��P�UL1Q�)�f����th�`%�E5t��(��+�j$�ǌ�)f�����A�w+��Ĭ��C�8�$����%t�j�7�kjRx���Ig<Ԙ�s}x����A�'廙���QQm�e;�q;r�Oך��ϯi��z��i}��`��Y|��y���b ����Jq�=�����o�~�ss�:�q@�n�"4�E�%N�[����{ZK�`n�/1�)BC�۽���s�2��"��=�A�5��e��<i(�V)��l����䗎�J�>���#�-Us�5�_��6����Fz2����o5�i\*�3� ,�A������LK減�
�3�p.�1�/�VI�)��YQK�h[����������Q�"�����J���ieQ0oU���>��ׇ�YsG۾��v$���Ҹ�ոw�+=HP��Rm���n�d��:����TD��B�p������rY�V��Ku���F(D�!��v�U��w���[6_�����qp�Ui9-uc���d^���
AӍ5�c�Cr9�/~b�f*��E�m��#(8�k��`��t��sQ3�ž��,oi����?�Fݟ��A��t-C�)2,��-t�U:f7���Ä��)�~N������o�%	�"�|�Rh>�<���RvZs�X�SI=�1�p!+/8���.)�3�uw-�JPIU[�W����^�p�}���㱊}���a9�6vIP�?f���ܾ3�[f{P_Eo�2B��_�m�冔�Щ��-�]ᤨ��6F�6�NX<_ŕ{4�+�5$����[��4��ʹ�#0�j�r|Z�D#5�0�ow�| �;�E�7�>D�O����#�����-��dJ&��zYMf�	숺��6�{	0�d6$�&~���OfWװzڝ�1bL˝���T����U�V�*v05ri�v\p��D���u?���tF�)��n���[1wW����${0�ﴏ�]a�9ޢ��p��.�i�c��`og� ��٥�\��j��$��In��V��}���4�� Ω�ڑ�Ѫ�N�W�|5P]�6mc� ]"E[x�چS��O�N®���i�."�m��Z���KdD1w�2��I1�o�G��n�� B�VC�v
�g�K��a�Δ,���
%!g�+���ЈY���>>O�\.F�d0�3^�b�j�E�:fFJ���݉�ȹA���"�y�����{!�����;�
�^;3�]jCRZ��<�M�ǐ�7ȶp�i�8_qxm�o<�悒�sr+#vJ�u���_^ych�i�,/�؅���4N��h%	e�3V�/VU��^�w�j\�Q���p�4;�G��$Bx����H|���u��Kg������I+X��Ԅ�+�ͳN�����
F	C���|�V�k�^�{���n�d��etGy��������##si���upi���Jr�A��Ha�"�$���Z�0tw���kt8'ðh��� ����__5zɐ3μ��5�y��36�_����a'Ɠc7n���2�U�P$��e���`�G�9iE�pB��s��J	q̉�fޛ������!т{J�th3W�h�4��'��l�-�L�XhYP���j�t��o�nycs�IUЁ"�:�#�4R�q
{z����@	$�n��~����Y\Տ�Uí'����n�����!�"��΃'SG1��$~w}��Q�;��˲�����/&9IH�j�!蓔K�2�[��Y��>n1��|ߟ5J�xj} ;G{���`bP�^�F�00�W#����5H��V�'�֕�;L��UP|��W��8fK��ض��x��-#�-��*���1����\i?��M@����?��.��!�Oɝ>Ȇ�D�zhm�3����"!lu.�?�k٪ݳԿ�ש'�<� ��c|�	ԡّ��Z���1�&�Ы�fOV{�;�b�W�������)�4K_@��6-i�9�Kã��9N��1��C�t5k�/ae#&X�j�c�ڿ��ߊ�K1m��y�w&ˎ����/��tf��2�'���Cl�]�nN�_L�I���,Jpn�]_����?�=>F{~Oua�̫X�S		��S�����U�8��D��1�W�"B�����:"2��s���� ((��ۥ��ʑ��m�'�]<�iE!>�R��K��)��a��8��-Ҫ/ ��,F�Ȥ)Mg�I8�
�"^Kwg�o�Q��,���uSq�ι�Ϯ�Fi"��C��q�����kbG�@Y��g����"��	�1�R���}#+���J?�u~�+��}?�zs,
�5�4�O��az�>ᡨ�i�d؍�ۧ�$(݁��0c�AN�h��U����,!ײ�qD{���q�����|���ʰŰzi�SeFhK�3D[±��
�
��N��'$�(�O���fE�_��b�¯�������/2a[l���C�WaOd�
�J�*A��p�b�b���Q?�A���]ѯ0����	���i'p�]�"�V�{hd,V`�Q��%�3<׿�s�1�bE�xTZ�W+�Yv�q�u�<<ڤVi���s�+��Fm�i&���+|�9y&���F����HнCLZIV���(|�kad��hYň畳�-Z�m����XG�̤Rr!в�%�%UhI�	;��Xi_���ڳѯ2�K���`i?8.����̯��3JV��}q-�2Qb�Z�I��{�.��Ȥi\�s��(�r�� F5�q��������ͥ$TҌ����G0K���ss�L���V��7T����&)���S����N�(�*s]���Z�bR!�-3�0U>�5#�3�2R��UiO�l������ɹ� ���w)ni�A��N(i�k�'�6��E`���屦�[�"�;Q;F��>��e���Ƞ��EX6����/�$�2^��S����,��F7����'�R����~��(����\l�U�g�[R��K�h�pz-�c�p"LQ2����y�Pg\���2W���͊u	/��gr�.��G��f7�]'��ʐ����j���E���fG�ʩo8�(Z����X���(���_��%�t���Td��f��,��4��E�a�7��o�u��]=�q~/����\�cqs���o�S�����S����8߭=�.+2��z��F,�GQ�?HZ������B�٧�Sًb� ���(WN5~W�n� .9���S��G�S����ב�/"���ɩB<x���_h{I{��>�e�a���-���X��8��H�s�cO�t&p`ނ���];�� �!���¾X�SO��7=3������Z�G�R�_R6�`�W�D�,�A9�zp!��:���N�o�V��Kg�IWP_s,at5U��@f90�Y	S6�}u�H��?L)���|W?��nr�U�h���J�+��]	{x:s��S���r�w>Ě�����ڛ�(���x�l�f����@��T���ɋ���p(��W

 (T;��Φ`f}��u�Oê�՛��,>�pm~�:-�c�Q�25�2\*z��'�a,�K�,r�K_#�k3s?M}v���7X6}�
��g���V�j��ٶ��a�����y^��ҩ��t�s���aG�آ��~5�N]�&��s�H�Ǳ��=cHwZ#2Ț$iW&�>��e���z�<����ٶ� ��!� 
����/��u��{<���|�)n�}���̣4�c��I���� ��0��lG^<w	�gbp Cd�>���nL5�Ӽ�w�ܑ�����Q�wK�Ⱥ$�D�>n����:sa�쁃J��a�c�8Xj��z��|�mx��,�����3�����'�A�1xW��^G�n�1BKP���x,2[��UNUZ�=�zgF�����V���kO������Pp�h:֙�'����W:06���+�B�ζrP��*��(�.��Z�>���ׅ���2��B�`KT�j���X^�z.�� �X�:�*�0ܠ�m\�����9��Taӄ��O+g-�@��w�<ehX��3�����K�ȏ��Zd�J8�_� �VA�O�f5�ͬ_-�HӤ����Lp�aw�Gp%�zy3���Y�B��[�>����p����o�Ӗh*oT�����S)����Q��U�2^z�|�Đ�^}B�e7���)O����Hu�f��X��<�͞zf�,ֈv@�ĵ������'���ٰ)�:�˔�y���>�<g�x���k���RE�ڐ�%�K �.��m�v���I���Q]{���ʳ�.�;N��pja��aCDB{��7Τޅw�tQӦ���^��`�3�)�,;��++��ʲ���T�\��ֈ���G�8f�08�N;�v��Ѫ�(T:�����L79����M�ʛ���v� ���K�j{P���k�;��������l�Јl�/�|�@�A!ka�$=;X�5~�l?��1>u���i%o����4�%�������_��W�G[��OӰ_%s�)��K_�g	}�WE~;}�5[7NJ�~������S�k�+-1�����^\W�`|ǆ.e6�j���4�JGa���CO�ñMA�(,ɰ]9xg�������<����ࢎ�,d�f9?Q���6�����2�wP 	m8q��Q��9��e����2ƦO����]=.Mm	yl8"菆���� �F�lk
�fP��#Xy�sYd��tΏG4��+Es��~i��כ�_ۛ;�"�Hd>���no��{���3!� ����d��z^�b����ww;��˸I$}8��y���H�����WN��d�-
�� �B� 3 ����W�۫�dNrm�5���1��|���q����
e�ݻ�_�/F��1e}}�14������ɺ*�Rx
	��zc�0���K�G�Ȉ"���a�o���S�� ��x�-�������p���
56�k���Om����xt(e̢��:���]:}��R��	f�ʒ�ÙI�W����|`����O�$�o d�s�v�Ɯ����ڠ$������ئ�Y-�xE)�֬c� �V����Q���D�˥��v��.�~_�5���v3y�����ؘ�V&�Ȩ���u&|��zc��(*�[��u�)�	nI�S��0k�՞LO`p�L���ո���F焧�.n膖M�_b�{��oJi�)�}Nf���r�bMʪI�[���g7�R�t�miT�(���աn%������b��D�Z��9�@+=m�U���Q!�ߢ�H�"�'��u3N�ͯ�B˪?��;��@Ͱ�u�ذ�A ~��󤭶T�J���7��cp!�x}>U!��i�c���I�L�"���M���j��6EY��M�������H01��{�|�0�ixj����e�Rg�H��Gy�5��s2�q*ʏ� ��N]����W��[�Gy�nv��F*"��K�bf��	�w�?:/�x�i�g�	�Q���@6.�S�������.����2�dc��y�D�uD��	wxC��s;��CxD��G�������������1OMbPFYQ=� �0�S�CX���u��c=��r������j*ȝ����]�_JKS�`$A´v�����k���;�}4{(T4�3�ci�9 �x���2�s��%EY�@���'�6vOn�Y����6Qߣ��V�)�0
���_Ƭ;hv@�2���QS�D�6k'��{4p�4�r��r%��}HQ7A�a���pE��6�Y��/J��v�Z2cn"%�w(�e6$� 4]�w���_��MK�A�f�=}��)A�;.�(��rr�%	��D_z8\�j�c;$�W
�֑�u9L��mne�(��r�g��B�KW@�pb<�w��tRŕ�I�͠���R<�=!��N����D4�2�Ph���%�plaeؑ+��c���|T��;G1b�S��9��5h����j ��U���ml�.�%��A�_�"l��@3�S�ҽ�Z� l�C|h`tC���X����];xθ 8��7 ��U���N���\!�u��H��rˇ/�@2��z �.!g�)����0۹�6��j�+ǰ$�3��Ku��M�!�{�j0�Qnl��I��w(���fD0��H��O�u�#�� ��fv��e��	㸖��u�W��*�f�Ed��+� V�\wr�L��>]�����J`3�6Q�߇[E����؆�������b�V����a�E�	��CA���bz�*GB���5��i�^�OĽ����*��F�� #��z��Bc�Eh@��}1�������!�t��I��_�������-�7e��I������]��\�0�>��cE}ya���!++�ł1���*!|��=�g�X\2���f
j.�N�|0���Gi�U�iҍ�;u����;ǊL_��*�{=��Q`Z��1�J�-�Ѿ�G�ա��%Z�|�c�% �)�y&9 �P�4l3е��
iӊsI�2A{z����~"Ds��e,!�`R��d�D})�T�9Ҽ���@[�4Ѓ�죯�g�rl�׺�G��G3��o%,��E�a4lK�z�g�g?ն� ,lydf�P?ga!W�ߍn x0	�E^%ǋa��£��3�(���9ژ(k���V����铉�C��2U��7P�0S��32yb�W��)��0WMx�a]�՟����`�A�j�^:����l(��_�E�X�]���2 �\���-�2]W�u���;�n�d�	\�5:PB�B���N�=���x���@�Y��x`<���oCV������ld&(�[��`�w���
5�sϏ�"���vX�Dvuv�v��t��7�J,=���qIW[e�+�e�A%�C��=�V�{ϓ��6K���ل���� o������h�?�bce�(3�w��9����|�V>�]�e_tL�atE #럋m-�ۥ���-qb�>Y���w�nP��9Xޣd؉�\(��p=Bg��{Dq'��ޮ��oۋ3AZ=mNx�ϳ/�&�
*��>��h��0���@�͐�:�i�������뿇o�c0�����<����v�U+����O�S��0�u)��kx,��g�Ő�S���� W���j4v� ���W+2C����ꞑ�W�
63P(�ëơAp-P�h`d������_��T���x���Z���֬���6��V8�6{rp
L�
d���[�Z�����i	�c<��aq�*Y1��������� ��is���������t�$�]3C@�u
M�t]�oS�V̋�75urt�LwOq�(F%�f�`m�n�}�z��[Rc@��m�R4^��0�����e8��D�\8��꣯�ix�O*z�K������ٰ�0�,�7�� $�������S4�eve\m$��a��[g��ie���_����<��\;F+㍅L���<a3O�N�R� J�;w�s�����Bk/e��L�9?�bno�`O�g�0�/��q�/q���W2�Qg(VK�"'M�ex$�p�}$D�K^�yD$�1f�ɜ��`�@���eiR Z� RR�� ݡ��w^g�K�.w1\���P!rf	�Vѻ�N�U�j�-�u����.)Ѕ,@�N�B
Ҝ6��/�(�o;�}��T�n��0S�+�4K�h؍&���~˟���ʓJ����%6ľ�춄��N��r�b��["a�9Bp���>k�R����ք���X�e����5��t�d\��H��#�*k$�O�'��@%��+�51By�uxTQ�IO~��
�YC�},p���������ó��K�M���GZYe�Tɿ��hfLu�{��C��[$�Q��J�X�Y�lf|[D�`����Z[������p��}� Z9�����ҩ/-�/�8a�2��y/>��6I1&��{UV��7�c����-tbq�v�YxO=�J�E����y���߬��(�{>���{A_,^؛����p�ũ+#��T���x5��
h�E�c�x��q�YZt
6҈�k�E�MFq�њI�<蔶WW���"Z�4_k%eܑ攞L ��a���*̲4�=uu]P�hl�Mr���F���K��W4�Rrݱ��x��)4���C�u�e\�J����3�����D��b�>�ƒ���OhQ�n,��td"h�	A���-�u��\�|������[&c�5�l���-����P&�i�7��ؕ��H�ЀtEƪ�����BV�ȡ�8ilE�JV�êͻs����s������8Xfxb˾��wZn2�����,���uS��F��}B�:Iq����7gK�ݨ5[ ��Rz0B���81�7���� ���j�3��ΞC�������-����4�T,����C���0��w��~�;����_wz�/���^7�1�f�e�G2�k�i�����3�ef�'�Չ�2p�˥���<����p#�Y���Ҕ� ��嗧��	�{��U�EP%�ح;�P��-Û	�����-�-��뭲G�i�O��u�&�����`t=�}٢������:��_1'���Q+\�څ�LF(ep�#�L'��`�:��_��U�IN����� h�E����{�����IՑ`x�O�����d��|�׆�>����:�*��!�kVF�}��c�5l�g�\�ΐ�� �PBhu8�a#��*@L��N2@�e߸ԝ9��3+c������/��D���x<�o�\R��=�|���hKH��2�:U�qL�����2G�i=�{��͈�[�}�p�8�4�FI݊	����,�H���	�U�^2E�ߵ�:5j�Հ���n�G���i~�}�*{ps%��<pFV�'E�Sz��Ika� ��3`�tNQ���n�6�Gsp5�?1.]`��4i�������ϔ?� �����?u:���s�|�ȹyvO�y����@ѽ����c�4I���п[���n������� �_���!�.��ھ�w��愶z˟W�v��,�>��.H�x�l�ݝ�)	�o���6sܠ���
O���Q�RB���(f9�=�졓`u�7S`�Z�s0�҈IA���k"fÓ����s��� �4[��%A9�\e2�V�:-�?���GH6��+��S._"�J�� �SdD?�e�����f��׌� :)�E�~~�B����\a�8���\sFu�%(������IWyg� l���ʤ�����&=|�/|�-���o�ރ�7�F��E��L����F����B9�ZI�A�H�����V