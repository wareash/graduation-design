��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jåا{�\�u�?߷�dn@6�zf��r������; mt�M}Fq) +����O�e�16����0���+e	�Ѯ�6����M��>}����A�jK� ��ǧG����K�f'�a������P�_C�~���1lK�u�g�F�L%��St��	�����wY�*�Gy8e�p[=��ΟZ��f_tߝ���G��4-���+N]��9�9R�
�q�/��Z{��s;�	���
�O�2�ޱ,D����_�K����-,��q5P`��9���/g�z���B�h@d�+�zY��j���>Ú*�O�F�s��>��L��q'i܆�]�@H~H�s�*.s����BU���� �j���,@��+�N�͝�?�C�r�ɏ�K"�>S�ۢ$� 69T�c���A^�q�WoEe�E޺�+i<PB1x:j����Bp��E[�����}����Uz%�DY'�����b�_�`���׳�\������v��N0�d�~�0!�3nf��bY�ʣ���|����d�a��x:*E�]r�\�9��&KS���U����A��R�^� AB��"��
��;���򦑳��}<x$�`�g�&�.��O�sxk�_-���4�����Æ+L�ʠ�2Sclq�AU��L�rwL�7�n�}FF;,��R��Փ�����ц .K �t���Ҙ���#i3�aO�7&=�D���,��F�SI��`0l�9na�����h(�UĸG�=X憍�D�{WIh�'dp (�!���]�YF��{=F0���ӆЖ;�X�0I���+����6J/ܿZƖ^$9zU��p�Kc�~�����OrK~�����De�����N�4�Ϝ�Y�tZq��
tfa�9���[�2�֙����P��2�R�k!w�*sUnW�3��P�m��L���1���}4ݿ�ĞE���&o����5�]f�-�����ʯ�p��L�X�NCS����ē�Yi��-�v5�'P�<O�X-!4T�i���Q�������kV3M[ʛ!S��}�3�D1�?�;��R�]ۄ2j��pZ& v����lmV%�<��aX��6�+��P(�+��䣠a Ț���y��1�D�}�:�aޞ��J���줓��ks
�)L)�p��KH	j�/��F,P��H�����ׁ�>?OiBgf���r�������_�ۓ|2u�!)��>��s�B�.�Q��[�-�Q�Bp�{��3)3�jBs/ Xy��g?tC<��Ҩ��O�Xh'O��&^tZ�8�؁��>[�e)�s<�`娉]���#O��C��ȯ����DS���yt�%����/6���O0��f��H�*ے�����޷ɒ�^d:�C(g*���+���!�l��Uɣ�,���(Po}]�y:�:$x`�q'�^ֽ���9�C&���}�CD�}����y�sD�_\?�īJ������:�+{�Ҽ7�b��Y��n�G8q�����|�が|�ңY(��+�3��
�YEnH�ߜ��:助Q���'_-<�k��DMi���{Ԡ��a/�GɊ�؟�l����>�B+�n*}A|BƬ��?�n�����]u9q����5m�᩶Ī���v�h�����;U>�d�=�p5T�+�y4�����Ɠ����\���^7���_��r��u}�خ?��w�%�MzO}m��~C��m���!2W�8���!�k��9�zQ�s�_���k4���(Z��t3�Lf��N��}�D�NA�>mm������hA�/fgۙ�o��mF&��w������g6ߟ�9�a��KZ-�(Z���}\<�+k��m��.�#L|���V�y҆(�]�~Ïs#&����U0�"���5U��F���"Q�K.��54e*�h��\��g�:��]@�#�ع���\/���t�e��ha@ҁ9U���:����f#t��=�tӓ���}�7�\̑���(T�_W����r�A
�N���VS���?�Or��B2Ap}%^1�fsE��_�-�<��@�bn���@�D[Q�ƍt�e�7C-
c-g�K����u�"�${A
�KN[�/xJ/�Ļ��33s q�s�?x�����qȓjt}�1G��2��?δq��`�nu�р:�I>3��{N���QvF�f�X+W�Y���$��YKI���j�A�:4e���4x<�y���{�L�>�[��o��Z��{B(sS�v�\�:t��� �ki�k�G|6�_�v�*T�*�i�Q2��n�T�薜�~��d�����s��J]�
��N@J�x�m�F$k��c�N�:�]�����h�T��x<�<���#1Bt�����!ĂE���s��]�[,��w������/�{��K�n�i���[kF%����-oPӚy��� h�竰��6�c\����*�� �r�
�_��9��)�/����uol=Hn�N�G�|�\�<���dx'?ֈk��VG�;�6�ǫ��,�ߡ��B�o�F��}:�Q��|>5^��v|�#y}�/�A����C^>P�D��e6� L����h�i���:�D%W%�Fƕ�k+��Qǿ����o�djޗ�U�U
��bgȡV�xԮQxl�W�kr����?,�щق���t���!�f�C6���x�@(�[W��3'�Fz���7�}��D��Ë�~����4��=C0"�-İ�~��c~̀��C�������8+���� ~w����<�&n�Ӭ��}��_��f�y���:g��w�i�1����������T�*4���*J��&Y-9ޟ��(��|׹�n�yK�|g�;o|�)ȱ��e�oy@e>~�.OTZ�q���l��z�p�J��䯻�(=���Jw{�I'O{�eN��tW��4��t��0y?U����I9���s��9UKU�x��+���m��]��Hɿ҈P��7�:����y�,P4]��֋mV�(�R7�"'))JD�F��
�݄����/HI.�V��M#�t����$26hb�ȊH���xq���-ע�M�r2��F,0��~�*C�9���.�1���)�!�q1���^&�i?�yb��]��P����WVd�%Iv4l�,�Lln�]�s[����VO��Gg�@ �c���rl]Q9y�D�u�� �;��-a-�Eu�-��oĠ'�H���3Cݲ3+�w'���cn5��k�T��� �~|\w鴕Ws�2��z�c�>	:��fD?2���oD�g�ɶ���:d�4w�8��<��(.�E���I�N�|H��㥺������PN��t\�Ղ��^Q]��6���zZ�q��Ɲ��V�&��VHL�.��򣴐B5́�C��:M�bV=_8LP�Z(u����b��G%�?�T�"�-���O�>♣�T#���,{9g?��� #!<�������/�
y��r[��0�P
|_1�X���yf��Ugĉ�ށͯ����a	�O���*nT�L0�O��p��D�;"D�P�Քn^��b���X�/(D"�su�z��"��j�y��N��\~�2��ϸ���n�&}�nVN��] �_��������tE�D�a{٧�S�UVg#�	��j���'���#����k^���{0�;($��Lz|ڊ�5tf �����L{�l�d�G��&�<n�|՞,U��u�<-ȳ�-�.� =��:x��[��Hی�*��n����oG�6�A��"_�J�v���0y/���x��A�K6��p0����ڕ����I��f���T��Y�E�osx�d�<���FO�p4�:�z{L�{��L�)"��R�\�F9����}���h�p�6)�O���eƊ����Q%���
��GLE�%ɽ�N�a�.`gK`���q���ݓ����ce���Qz$�r�c�0�SmB/��%@��Qv��	� �M���X�	�*|��@�2���R��k_��c���EYW 3�I#@�Q�fP�r@�ii*���B�v �%u�羅,�д^ve���)�� +X���M4$5�x��5�œ>F����f�λ�m�3hv���(�*�+5�T��:/t`��s�-���|�=�x�#^��_,�\`��W�ec��� �D��+���87�B�*�F4.���M9�����4�%Rr�R?m����%PYy��b1{ІӞ��~!~5S"w���V@@vn��T>��ɘ��$3�m7\]���e�i ˉaG�#�[�$v��>�"�ɻ~Ç�Q88yn,�����%T�n�߷���Rvv_aCX��/����X��=R��}�7��	�][�/�+Q�=qc����u�K�2*�	�&��]�5ua{�2,���a|�z�apQNI�O�A�𗷄��W�J�ZN�{hk#�\�/���mI8@K�컐t^ѩ
�����N���83t1����s#+���g���v���$ˊ�~��WSmYB䚄� ø�*J
U����Q���h�{ʧ{������ޢ�1��Ws��e�v����.���l���Vɧ֙���}Շe��UyXfq��	�TQw�d��'ic��㴿MzǍ�k{��Q|�l�_5F�]�sӍ��C@���@�r�S�bm<�[}�P:)K�2�l�����ϫa�7�-�ǒ.��3а.vV�����\$Rġ�֜�!ׂ��T��Z� ��xz������,І����ݘ��\����$���ıl�@N�� �q�Vk'�az9]F"EA$����"		��ɇ�dYV-�]
&��r�*��ޢ,��N9NS{](�H��n]Y���4�ݔev����/��wJ�&�q���~�j�*�����	���舐�f�</l���1\�"�=0���z�&O������t-�p-�&�}a1�R�ؼ�����q�-��X�+�(0r�i<�\ձ]?�����*����#��a���mP%^���[��R1#��+��b������	�6m����TAd����wX2�|�q���'M���o����ʭp6��喲	���0~�ֲ0�G����E�>�}
����:�����u�n+7/�lF	��~��$*��˶�~�o��u��q|��E��г�kBl1&��J2{_��	�8��:��(h�	�w���c���eE��O:���1m���5"F��v��w�L����+��t�>�߻�\3y��"�j���n�⸁&p.��m0z|Jm;'�~9�#��@��-J���&cV_�R�*?|a�2��D#3�瓊hSfϧ��'�ky~}p��0��x%K13���,�����A۩/.dCC�(����ǹ�g|-��!�dmVukǒg-%*��NO]��+:4*B�ۡ�,dJl�ioK0b�m�g1=/R������Z5B;oK��2*��1���A���{�P�aCy���ǡ��#+�>�فQS^N���^����f_�/'����Ŝ�̞�ٓ��b�y&����Y��q֩�5j�՞Z����=���&��c�1 ���(��n��Ò�bf�`��9w��%�v_�����sy�8��HnrY���t�.�ԁ*	��Sc�L<B/����z8���)Va�v���@T,Ԇ8s�o�Č�v>�VyY���'G���^�{1bPc���(3��U�~ ��Ɲr�a�)t/�bJa�`ه�Lִ&���"�I�] ���&�1 �cE7��Ϛ��3:�}8n�b@�5��jWw�@^�1��<��Պ�6 ��P�!�����>��D�.�B涃F�r$�Lm��6J���eo�6}yA���:*Pd�1J)��
6�`��3����؃�N����Ȣ;,�l��H���1fR�|�a��7�1�/�p��~�ӡdj��B.�F�~K�����Mpjk�Y����D��F*ܱ+����� ���{�>L0�I�Z>�ܯ>�Z�xX�݂v���z���D��t��IF��9�=E����L�q����Id=���1ר���\@E#�Y���0�_���xZn��1N�(Zi�
6k�vB����T�a\�!j
�}L{q�ԡ\,3f{C�rWYꢑ�)����u��R�ahߧ3���g�%݆��[k�8#��s���])�͜/�7�%���-͚�p���MM�u�܁>Lr������F������[���~k�2r<�f�p֘�G�7C�;�E�j�;i��2��L���`^�s_(;��Í
�YR���?Z�pA}o����Z�޺7rD/�@��~3��,�(�Մ;��	�Ǩ����w�emn_�u��0�f͇�����Z�����wcl�ul3�6�fmF�+�ߣ��A�3`bB���?��}(�]P����G��<S���<"�[5��*+�=�;ݣҁv�8q�Hǁx4
I�=�7�B��ԓ:Ɋ��{ɺޚe[_�LH�3�$^78�h~A��6�\-�>P�?����7�������~dw2����ch��>9�;*C��h	�G���Z�L �����<RX��R���	�Ī�
���-	H�ޱ��۸ ��a�H1;��Z�*}�!��U%Ө��JA��H+}w��Mn$GA��'���X>J$��\�	;��ӂ$�B�!f�S9�)��Q�(�_M��?^�S{`Ó���V�_�s�;�B u��jY�tb/G\,�����l�/�� #��	�u��,�����(B��5�a	yΛ@��/�$K���KK�G՜iw>]k�X���d?`�\s؂��)����nVn�d7��I�����	��9���@��T��m��ӵ珄�f�+&���É�� ��G�m�����2ѹ$�ǟ�jh�H��9O/��#2%X仲|��g�l�:Q�c��Vw�O��f{(�2].%���l�C�W��=%Y������	�i�-�Ŷ_�����;��OPݣ�P�VM�R�\��R�8Aĺl�H&��%k�M�2���^m��Vi�c��Iy1bɗ���SZt�K`��>%���V���ܫ]Q�`!Ɣ���!�D�>��h1�3�@����YLזݑ�=�Ihc�?4�l�"�6J�)� T�]ַǗ��ANؖ�${6�ۍhc'��Ʉ}�>��Ib��ǃT��aL�|[dT�'2�Hc$��/�Q?�_�r�{�Kevf�b�l,i /gf��S�ќg'���޴(+�,�?�M]�)��޳Pkh�N����qe�}N%�o`�+����������}�0��K�r�#u��S�p���<��ˠ�6����j�n�13�2a���ߣ`�^"�O<�&�NQ���Z]e3�2'9L�����,���ʬ��uZ2hF�H�twS7�e-��E����濆���1��"�'y�a�$t�ː���rzI�F� 
��Q zN��WK*�3���Ph�-`�4�ѝ'�l;6 `W���Nr�?]�ʺ@m��m#�Ok5/o���.�)�sZ��P�F�-gC��W�l������]��u��Q	|���ǘ���U6�PD�+�B3����Dae���΄2$�bFĂ)��N��7��Y;P��i;���F��u�R�V����n�J�`���L*\�(��g���5xv��ќ�j�%?�p��̃�	F�h��\���X�b(^~�"ac�c��Q�ں�M�����î�
%0X�d��Sh˳{&U<�-P��Yy�Xg���ӑT֣;Js�Qz)�"���G��r�������"�1#j��U�Vv`Q�t�݃����Q���Z3��mK��,f��.M��*^�c�_����x���wa���Z���a��gC����.r�n�Ӄ�� �1W�)E�-k�>T�N")V�?��n�/Bݨ��&'d%l+��d���$�ۨ����3	�gI5���� P���4����+�1�?t��X{�fO�໶�-i��%�F�̳_�yBOx�@zw �hg�ǆ��+1���#e�˵�l��R��FL�����oD]G̢%��`��Aͽw5bv?փ]3����FC^A��i&ϔ���'���'��[ڼT�5��l)������~��m���˜��=%L���BPןjL�S�s�h�Ypǁ��i�������eg�h�=M|����^�^K
>rd��m���2���ZW�n*�U.�@�k�@�њ�O�3��K��k��.�� �aZl}w���9O��݊N>�}\��R��2�����+NK�b_��C �D��kA�>[#���v�`ر��0�C��w��k�5�;A�h����Q��Ȼ����W�K��T��xl�Ø=2��)J�T�%�z"��1��^��5��#�a�v�)W
�Q�N��X���QN���7�	�{��
�a<^̀L�.B~���V��-yP��ZxE�L����sA������^_�C]<?�c���v��|м4k(@1�*�!���n�if���Z�`�]0�Y}��r���G�ĺ�f�"�L�<��Q�w����L9���M"�N�U9��Z�*{ǃ�a�w��2.h��تԝW�u�eܝ���芇�a�����	�X��j^"����X{_���AL�p���7��S�Vi�3Ƽ="����v� �	�KobSW�!�����+��-�`bn�u"��g/Kw������>�-HW��_lP^������Í
����/ei��Oǧ�X�O#�P\���A)�!��k:ֵ	y��DZ��~��Ҳ ���T�[�	�[��y�_u�.�@�����sHm�:�b&X�/:���U3G�����ۈM�Fm0ӟ��=@�_ն�(ų ����>&Ԉ*Q��.�/j�7y[�d,\��8�SI��)�����pv�p�\w��A��Z���@�jܔ�7z��X�ZЬ��*ǆ��N�?h��f�-?;���R�.J�N=�W�9?7�������a�e!+�1�k����C���?]ȳx�N@�.� �-c1rk+[�}�������%�=;~<����3N�V��Ӽ��G/�]�E;�X���V����5��cʇ�)n�68����������f����ipV���V�rf�\�ϭ{z�;��HU�|���M����K��m�����}��ą�Т@M�|�,0�m����W&\��ʴY��@����,k����co�i֖�2�ݣRR5}+~R���n��ag_�2�u���1Xn%2_�����y�R=X�7��\b��!�����|k�*�'�b��FLK�=WK;��9�	%�\cCm�x1�i�������ѤTz:q`�q��&'z�I;�V�ΠF�bl��Y��i�-Y�}�:�f�m�v�b�����)�2�2�)��=`�ub�M�3���w~R���Y��R�+�fV�kS�q*{�H�u�*�z2����tz�ϒ�0��̻cC�j7�K�ٳms.|'����YU[&�9�� ��մuoOJ)�炝���kR���kT|M0��(���ݩ����r;/�o�.c��e9��1,o��Ƈ���]�n�1��&��F�Z��[2(_�V-�TI�a�@&&o�����MUҋ�,d<�Q�����y	!��C�T6	ZI9����A��Ƒ��ݠA���
��.��<et����v+!�rC��[���RR�Aw>.r9M}����EBސ�,��*�����;R������/4����*��I�I�\����D��,��,~};��퉦���
!NF9bt{c�W�/n�P D\���͋7B3�M�5����ߎ!���?te/<��}y�'֗��٘�G0��j8񏨄���=�$�	�yD5Z)�x�p�=d��\J]7�q]��
�7/S]�Da:6"`�@!�I����ϫ��h���5��}� ��P[��ˁ�ٻc�kCp%B��u���36���TW��QVW�3gs�ٸ��_UNћ�T��g���]�뎕��n�xk�t��5�e��04ǭ��P��bF���HRȄ�.�n{�+U&k3Xgom�aW�l[TU�2SJ�xX$�T��f����\��n�*Y�����_JW��&�+����������w�Y��$���7U��X((�(�gK(�ϓBp�q�/�3ϟcQj���t^� �-fd�r�$���I���h�GXnҡ�M�:�Hl�q;��Ђ�|T�l�+Q�� �F�(V��lF�(�����4Nn�Ѐu���Ʉ}W��%�+s�mҙy~��$�� ��a��NE�.��H��!�T�U��~֩�!��i|�ǥ��}�Q{����Z̤Kͻg!M�����W�D.H͓����_X�~5�zy�ǀ�����b�@�>G����d�A@ߵ����"�;�H��5�����n��O|xk�%�Ĵ.�d��g�Ɩr����e@��#�/�:�j��]z2�=j��ִ�{��<�x��lؽ����$�f�s9��[Xu����I+`q&��-_�"�ʹ���V�J�����_��t��a�~*I�Ū�O��t�6BSb��@��m���I�&xB2�+h�S�w8�;@�]4K��45�G�Qv�<�=���H���>��F���p�t	��� 5�b��x�_�BL�����'�B���m���tzɨ�W'���4���
6���p_�۰r����^1��ٰ���<l�ٴ�.S�l!�'i�oq�I��;��au�+��	]%����i��<R��1\`� ��A��{W��x\1�y�F/��Z�O�Z��**L漧�&uS>��H�˵h%�����d\���H�Lf���G��#��,L3�zY,�⧽M�@��l;�Y�ޙZ����s�L��zb�4^q���Sk������m0!�b�WF9#���!;΍����_̍���@s�y�1�Y��/ꅡ�ے�i�ay.������r��s��J��08I&�) ��<�4Ky^�(�Y��:rޞ뚲�]����)�?����OJ��K��w�{aL���U�-յf��U�d�T[�Y�D!p���Q�8�8@��~edt��Cv���@��%���nX�~r3J|g�[�S��	t|��f^9��Z�8a*K�4�RO��]�����ЫlQ)D?��������,�!"Z>K)Pv;�x&̊C����r	Wp*]/�c���|zb `5�������R����Y��Uo��N,8���K';����ܮ̖m�?	9�$P���������r�7< �O��ݚ	;X���;��L�?̢P���o� CZ��\Z}�j�T���ֹ�n�3P�m�Gd���I��"Nٻ���F�NuN5:ܟ�E��q8�Y��J�#�箜�G�qRt3'��~�wI�ua�05�Q��d	�T��@��6e��"
��Z�E�!���΍{��9Yϧ���"g-UH��-KVb���n��D��?Sn���a�6k�.����{�8�#�>Y
����P9��.-c���}?����d�%+V2o'��2gτ6Z@�?��'0M�td
�00��R�K�j�sNd�9���`o��oP@u���:5�n�y-�����" ���r�,��A��"�,�G��0J�-o� *�pY��6[(��g����Y�(���~���y�kͽ{��,�����[T�3��sIy(k���Xz�v�e�y��m;o�#)|g"N8���)=V��I�Xc�!��Q�$�
o�%�	{�|��h	����T"N4��Q����ѳ�+
�b�׽��ef���p�Ue���. k�#潚����hJ%}�-g`=rE�H/�j�kT~�p�3sY��wh��7*ح�\��"2��؆$�b���C������K��"�iٽ�Sum�l?B��o�{?l�s����W(O���"���c��t.X1J$W9"�$*}���T�/��'f�::�.Y5�͡y���PDH?�ɋ�	F�E΀<y�{�\$�\��h�ȮӾÕ* ^�ݙz0�x�k6�j�9�.�*��rC�ku�j�S���u����r�����+��a���t� ��^��5٧�U��i�H x�&7�IࠤX)1��R10ߵ�����
T��Ѻ��7�l����l V-a��ՙ��F؇u_��\�_�fYt⽰��4�4�.>�
*G}c=�0r��>�5�Ɇ��6�)Y*��^�`w��±�=�N?�j�?P�NZC.+U��;�0C�;���s�.X��vv�����.�}��/p,�ް,'9��b����6��*�;^I�#��v-��x,��N��ɱ��0�ϞV�%x���WtL,]���x��E�D�Zc�N�iN© 颙�\��z'�
tA`��O�ە7 �٭P��=Mb�q���I}غ���r��V4�٨m��Ő�8~��h�pJ9�{���|�g�JvLm�[���+�:F�uk�$S�&�ewn�b:tg��U+�y�Q��)��"���z�R20q0���_1��A��3��G0�5��t���Lx��A�j6�,*⤡����$�s��Y�����%��o �KVd������<�ś�c�8{� DtX '�B�]6�h�>�As ���G�v�N��ҍ��Y";��]���3�.�:J!���}��ޱ�Ր�~����2 ��n��72�:^��uYx\$��V�ha^[#ya������Cn:�+s��-��V���o����Þ���ƍ�3
r$+���nkv��׬^ˎ?��a��l�t�#G�+E��88W�ز7O���=��C����
D�d���/�2>�z��Fg�!ƂU��Ǹ; nJ�wբ2�̴���	�BQW��Q��� =��UZ:ޛzYj���mi�Q>a*zKf�r۴�}u���GD	d�U�l��yfdg�B�>���y(2ܘ/�9
m���Bhŧ�$���U�_�]�
!JGG��E^�|������x"!�j�u�
(j��y�n�[c��r�($��ut1Qx6�ӿ$ҵ�~JQtu�q���kS��v�̀O"u���ֳ�%���e�K��i�fQO�]��� �<#��@ew�T�=8��� ��}mF��%?��0z��������;&ǋ0�y�%Խg���N1��=��Y&��5�N��n[0֥�}�h��4��&��=b!�HsE��7���-�$(�G7m���ƪh�{s�b����`(O�Y�?��>��<"����AjL����<�6.x:�ީ��	 ,�F��r�B�>S��>�^��1�$�X7�ڐ٠���y�e��S��C�of�E��bͷz��P��Ib�$��G��M�����s��#�������TQ�b.�����[���Q�%�X��H4�t��,�Ql��e}����ԾFm�ut�$�>�i�	�����7�eD�M#|`�s__�%qr,{�?	^W��̷}�vh;�j"��'���b��7�@��>�c&���/&�h�3��(L���Cd������+�Q���Ly��yN[C:�`YG�j�쮂r��s����f}�{H���g�[�p{8͏��1��K�<{�-�'W�
�c�)h�rh/��u���0�䥔�E\(�{;����c��2�����I_�ɿ��VB�Fs���%hJ���C��#��tDܛy��3�C`ar���-��"|
�/�ُލo��s)����آ/�T�,������*�u{@)�D��ƅ�w��/w�A>�-<M,�?�xӘY�@�Y�zv&�D4OW6ƴM�.v�$ ��w���g��2{F9�=^I��>�&V��S��_��.8α�K���P���aOv��"�\h�T?b�7��Ѽ�o#^|�9�&�$Jq.;�Z��{R`ѡ��K�g[�^��`?N=j���_$�Ж�.x0�7����B��z9Ӷ�lA���L��6�,���Ƶ��}��_:�}B|������e�-�\rU�\��������8~7
�;y��2�Ň�;@�j�^5��šVg�H��S��h�����{�?���m��1�I�Phe�q����V�����9fp�较���$��"�!ʀ�◘vd<Hd��TV�f��ރt�߳���DZ�˴��*E�s\G�W�W�=R�S	�d?��Z�_xS�~�I���/>����6^Z���$fL�(�>�}y/��+(z���DO��[5��S����Ng3�V����q�뚻�3�v0!���"3%���-\��&��#��7k$��b�]HJ)<3���E|�	��X�%B~�������>t!&*�5������ʨ0�ɣ>V�lv����B�Mu� �9�"N�����^����?��C\;�g�t��l�J[Z�'�����عqs����W��RD��`��qdyU�X���!	���ۿ�Ħpi༕�kH��ŀa�݀�q��ST~�6����&4��>�����V��]�<K�g<�U� oOo�b��+�>��[��/Y��궼+�M[r@�EU�.+&`ķ
B��ġr8��@"���'q��c�r�;'�k�6�;j�WW�aK���u�J)�w�^ٙ�r+���-�2>Bv��t8%L��]ֱ�#��?߂���ݱ=�Bȱ�V��9�I�.8R�.Mk( ����X�;��%���Q&'c1f�}�f�X+�5�۰6�Rxj��dS-]lڱ���	�,t�u�Ě��|��,�n�i�G����.�iS�Qt�n:}:M����x����Y���V�p���~t=�q���-�D����o�9"�IJR`b f3���`_��`E�ڿ�̦���oS ���K��5S9�a�)?�#%}�^K���]�Vˀ_+����Q	x��^�F� \b\ā�" ~����sp��mN�I�dZ���(,0r3��P=�jz�f>�з)�k��N#w���磈��7._r�՞��u�m��_*Ozs��� &�"͒W�
i*���4��89���l�Ggj�um��a��Y9
�`S���s�� �'ɊiG剭�����	G� �<�4�����6Zo��}.5�m��`�Ty�������'ܦ�||ѥ�c�W���֪lRm�/`�j�V��F�h5�B����%:���V~��8W��t��I�8��MV��jA�X:�,ͪ,����*4��*,��x3��h�*��k�K���(!�{�9�4~*`�K�a).]K~�'���	l:,mK�&Y�G�Vk����v:=�W���d��^��U���n�$��ʜ�����e%�QV� ��(2�Ǚ���c��A]�{)���q���	5�В�>V�����Q�'-���7ܱ��<]m0A�S�<�+f<k��Q��?�_��I:%Lэ9� �?����|��;�zV �3�� �(0 ���?���[`�Q�I�T|2-�o;2�W`��ǋZ��`^i�ƞ-���b�r8@�IɌ�o��r>�(mcCP}�o(p��w rڽFi��@t]�8��w9K6�_��Tƛ2��̮J
O	`<��V�w�O�e��c����B����ȋW����Z������ʰHp���tO�A=��!���i��ٔD�����8`��Z����:=~K� �	ʁ��;��d9�'o�2��Q{���Tʤ���x#3A_�Vo�1u?�tw����pnv�j-��D�j�?�%�q�E��>��E�a����]#_9������˯�DyT��������M��L�t3�4A�Rv�:��P)s7�8�-�DX��d[�򘟆tyNn���ƴ�WR`�L�9S���I%�,�&%�����K/u	ji��*]�pW��|�&�L�#yd�� q�߷^֪���>���,�F�}b�dd���(�=��ǽ{���W�)&0s�;��J����Å�`*V,Ҟ�q�1zRI/�r;���,<������Pgnf妶�$EⱠ���9~#[HF�1o2n�%���	y�D]�a�,���g2�A�f���ҏUy�KŐ���x#F8�jC�?k}D��W���gX���~�'�� �HgDf<b{�StJn��$*���
��+7�����������x����R���5�� �]����o�8�,~��5$q#�t���l��"���~~�y�=a"�[��7���x��lG�J��&���7�Ĉ�#����R∢���x�|��j�tJ�9F_��O��'����@�����}9��FLâՄ��F3��>Vզ�~.*8��K���V���t�2_���IG���n�²aQ���_v(Ry�Y^W�
/28���pY!�0��j�����(o��dHÁ"�k�'G^`n��f[˗YE@רGI$�-�0P�5̓FF_�P/
��	'��=�A�p�\��W�<g�I��S�۳��R8�hN����VA�T��k��0��h�F8���ӝ&��E���k2�H^}v��LHjW]Fۙ���2���Fu�[��� Þ^��q#�eɞr��Q�b	�~����̤2#��q1��J	�9ȗ��� &�����Y7*U.\p����t?#i0�~��!��Nz�7.�{��
��v����5l��������=u�,%�'c�����"���Z%�y��:kz;飯!��\!c�(Du��l��1�۔,YH��>�mPѫ�1:�����6Ҟ�}���a2*�U��W��x8W!�|�=��E�
S�Ը�6�4�3~�L��㼉~xS�n��b���A!�Z�/5 ���~;��i4��2�D�fS(І�O��Рm��0�����EÝ�e�e���w��VU|�	���4�S�v�i6�C�5��$k����sk����	I�G���VbK�9&������5�=�rpSb�[�d�i�\R��n���e��G=#�[�z(������n,� �����F�ޠ�%�
t�W]HC���͎�*�럔|�f��:��m<)��y���3�sB_h������ӑ���#OS��n�S�p�V�1go��L�λ��y��"�+� ���"��]��C���F}k��Yd�$T�f׺��*�^3�l����yu�:O�I3Z�5�Fm���d>��"}��W󵿽n�H�f�N����5�cK��[0l�����F|��k����h,+_;�w���\˖����N|�D'js�QPV{h�$Q�ԛ����� y�Pt�����ܱY��8���^$�e�ώ�qjOⰵm+w<,}.����.FT�{�>��?r�抠��$����z��+���ゃ���+n�
�c�t�͓�
)2��tw�Ë$ ����\��^��]�ɵ5�W�0a&k��_I�9������"�4�UTP�О����� T:IQ ���</i�~�Bd%M\��\�z�����L��5U1u���;w��QPy�����n���KH�Y�O�ۯw��d��0�~�i3�笔{$Wv+�L�Z�<�=�/�'~�i�i@�Ϊ;2m���7��u~kW,��5�"юP���j'�I;�F��b9^-�0��Viq�@�>��䟮3KP7�W�uSzWKX�Y?GW߲�&��R���h����^�%��<#z�����
�"^z�)��_��	E$����H��2��	�!����3�iQ�H�$���l���]����\��?�'" %aW��q����M���4j�!'����rIY|�s(�J��&]�|&dq��c�����LǊ�x*0�
��K.��%C)2�a3!oy����`I�h�1&���w{[�(s
�5_����K*�=$2&���_BLy����y
N+2#�ϓ���
	'Ξ��5�;���=Ȏ�3m����P�m@3�� ��=��u����e
�h�Pφȁ�A���$�)�E�X-��!a��m�/��&l���Ӟ���m���X����a��^�2{�a]�~y���:٩�8��-Eu(u�.��N��`�>�a�40���F�3��6؂%���(�u[G-s��9���CӶ��f��5��8�3\�,�H6�V��.���1��5�Xz�W���ͨ}R;�N�I���6�*g7$�����e9������q6F6V�X��s������٬���m����1*|���}D[���`:��Cֆ�X]�On��h�Z��"��N|1q6��־���-UB�� �b�PS��'�ϖ���$�dVM�(�kϢ=|j��>�v����S2G���r�h<c��v|�7,(�#ܛ���^w<o÷_Z(1l�������:�1���F|�����W�L�VlǨ��ߖH�w�S�W  �-C�[�t0j���Ka��N9d���9���1�drJ2���I�E$�<��Q���es�h,��tj�S&��|¹Wk�=#-��������������:BA�Hy�x��bj�A�(�h�����Kݠ�D�1Y��m╅|�M��k�7r�*OM6r@��ї9����`l�"{�H�^������������Vٶ� Ҟ&W�MK�t�}lTp��R�MJ���"�+�Aa�m�\�Htg@����ɏ�]�ފKr��/�v����9�#�/���.�a��O*�li{�0ϯ�+4��_B�E'�+�H�X��l8�q�l#�*VYW���j�ʒ�������é%˳�3�M��K���J䃄���2h��e���x(.[QT��T��]�F�����㸊Ǽ੺~6A�%w9h'!���w��e+�l�G����3h�H�=Gg�bƌ�ak�s4���1�`+v��`Z	u�*�����F�9�M������;��P!8��/���)������\6#�_��4�������Y]��M\+<9+(�e��}+�H/IEp�����wY���ǻ�E�5���q�U���@.��UQ]���v����J8�٩�G_w��?��'�5\|�`�9�T�� �΄�a�ЅU�7R5�N�X�k�>�Aۦ$0��h�ZÈ�P=�+:�F���'1����x���Tx;��j�Ŧ��([�5�ܿ����b��<����*7Jg���6���+��4u��[3�L+Kۓ����U����wU�X��\�8�@�	�#%�+��$��6�D_�O����X��b9�w�!�Z*c�ʡ���"����4BQ�:����/m��%���<�P*���P�]pnD_���&X%>���c�uѩ/�����A5����6�K�����g��9�n�9	��i�~J�7�L���h��l���i��;L��ᣡg��o�CT��0����&w����8ZF��K/� HH�E��������:!������C)�7�O����&����4�\�"�D.�7�����&
K��vz|�h_�<[S�p�a2X7�%=���W3�O\�Fʗ�%|��.��n�
j\�_��coVB���T��ưkԅn�W���� z�'�%�i�v��M'�g$��	{�����ڱ<-w,�y�qrj[�{
��(�Q�h�LL{�Nm�Ɯ��fAI���;��_��*�)y1$�u̪wT��&�O}G)��ꑰ�g���A��A�P�̀�GT2���f�|G�E(��ߙ�=+��������VV�ci���pE,<�> ӡ�@&D!ψ&U�g�&x[� VO_��[a4�X�6[�o�d샚��ww�6r�7������L��������Ȝ%��h��Uo ��*ks*�#��a\ټ�+J.��/�l1�S'���N�0�@�P����l��2�Ew���cya��PM�0�����g�Y�q��"�9J8�b�D9�0'G��[w`����ۏQ+�:3>)����ܣ�|���95��u��
��Ii�j9��G�("�����I��q:w���p�k<�#��	C3�����+3ν�"˰|]���6�W���~��Ke�N� ܲ<S�̒q��.����m�qX��\d.������߮�%�B=~	~xmh��3��b�)o����R�fՆ�冀����5��K�!���n�sNS��U��ܔ,��N���wI�?��Ј �I
���IU_��;2����\�<���!���$5�f�L�L�����T����j���9%�����FTT�[�B 󸼷c��[�D�.�2����I@a���J�6'��rB�?��<~f��Ο�T�� �Q���X�g�����,Ml�Q[�ߴ�/���Eɟ1{��%���hΘ\�)i!��Ene�I�q(�14]U�����µ���I+8��Z|`'$!�|�]���P���|_h���>C�Sm���nӮ|�J��q�p����
e���Řx@x<�İ3��]%~1�2�ܧ$ٮىnY1�@���ϩH"�=!�
��ὤ�d��8Т�+��6/��{Rڰ���إ�&�;�,NnEx2E��g��l�G����Ya��z�:Q#cϘ0�t��$�����y�~��v4pڿ��|(=\���Q)��9�9��H۱W���e������γ��Ȃ����j߾|x���&�l��~�y�xSGa�i��y3D�ΰg��`����4�&��9��@km\%��u-z�o�����dr�c$ލ�x�[�w��5�3���:(��� ���Aq����s1M Q�3PVc��E�o�>�,���tTcA��}6uv/���T�`�y�����EfO̺�y����u�ߦ-߭	T����m*7�9��ޟ�y-4+d��|V̦,�-X�};5�����p������fE5ǰ�SA'�?Ϸ��B�^t�X&Y��t�D
 &�pu��3>�XǕ<������_� F�Y� ْB��flC��`jRb���uQ͙G1��+�����R����r�e��J=�X��
�Ӆ���Q�N޴��R�*�@7��=Й�ϰ���9�#�x�V �S��=W��~�x`� ^�>=d=xP�$�6�38ajD���|�Wy}����W�*D��1㣚1@Ə��Qh#�� �J�%k��S������d���� �`%81�rT�_<�.V��8J]��a�k�vp{�3����RUĜKP1	:Vi[��y�ez�z��@�u�'\�Y��A���Q�,����h��6���W �}�μ;���C�� ��b`�u^��J��'��'�E���-������`��+N����{b���/"|%���:K�p�y������O�U/^0�nOy��Ѷc�N0���4x=�ꏣ��j���h.m�ŭ�EqAq�~o�y���2*^v6.�]�q���{��daIρ���	�K�_�d�0L��ǵjU�4��זz~ׂ	�.�}�:����P�K�V�-���X:��Î⷏,�	q�Q5=�q�����=���l��<zVg����/$M�\��P�vg���c���k���,@��J���a��k���F�!��8��Ih������)lmS�2I��3kR#�!:������moS�O�N�)���+��������g�p��l��Hw
)	s�A��@g�7�|�,���|�1�a`��nmncy'*����/0���m�b+E�����M�ܠ�c��g���mZS�|!MV~W�6��<y�����Y�����z;5�{�#hں|�ev��U��\iH�/.�k�c���{��hS���!�I�Z��)8a�=ܥa�#��e��.�kz��z�5rK�x�r��w�[���
#<�i�,�q��@��Z�]��C�?�(�԰��"�/��j��CG��]Fp���H�A�Mr1��J�i����_<�_�F>��|gh��dj�n��0<��}��\F��@n�����"D��Typx\"�]��AA1�Ƭ�wRΦ^�2��R�O�g8�u@7�IW��)�[�5��T%��	�(��_���B��\��o���q(��U�V�RT�e��e�G)����|��js��jZ�aGO�qr���k�D��$R�i8�ub�W~W� ���=�,*l@.�-|��Y�Ӈ�e���EQpK�l J� ��Q@�m\`�y�h���v�5�%R>�`k��2������ú0�s4̍�2'��Z:��hz�a�۩��4���J+�(޶�.�uzꡂF��tN>�D�"P�_ݎ�P�����,ѥ/��윕��~�$�eُ���q�58��Fkp&D�=n�Je!�&�7gMe�� �s��} a��W�Fc��8���e�wm���#UU�I�+Nz,�9�����C�$� �h9�ӕEw��GNIF!"�_�af��}�M�EH�:j`b{�����:�A�|�\�P+��]q0_���V�ikZ�氙ϓ֡J`�+�C�Ȭ�����8�5w�!�$!�5�$�08��)"�1����8��lq�T�h�ާ���	LF)oO�;���l������W+�(#�̢�t$_�
>����	�th3AU�j�2�c8%be	�� ��Iz)+G��Z*���O����gq4�{�>D���d�fZ}�?x��Y0k~h%��x��}?�/(��ҁ%�Y��η�ܜ7���n1�HB�̑��T*�l޽L�����U�ի�Ѵ��ʆ�L�Ff�����K[t��(�'��]��da2�o����R"=�O�Ke����x�,��$<h�6�v�W "��@���D~�ԃHw���5Iu�$!e#���@�o5~����e��׆���ǩ*�~�1:�W���.��̓�n�:[���ӨsHxQB�<�mѕ�&�E|hl��GoK�G¢CTkN���?�1����d%~Py�Jҥ���Wc��;��>"��p�r��̈́*�^�j�j��X�o�j�:�~�t3ފ|��O�T��{��}�w�5v��U3ET!x,ёߗ��u���޴"�<�jxh�����š��,�1���j�ji�Y��	`;�!Q���y��*į�ѿ3���xt Ċ~Z�ud��me)�)�}0,	3�NT#��ܼr���ؾ_'�:��D���qt�62r�|�%YԀW�r+� �2IH�'��C[�B+?�v�[�������Q��`�x�hGf*���玠Q2T)����s�����@��K�td</ߖ{��mN��Beb[eW��]���|�ȟ%7$d�½Q����P�*�Ty�����)ߛL��s�ц��@Sa�ْ[���~J�a��1J�m�}<�/i7�KZ��C[����C�19�ЫjJe��{��g`_X������c-�~�l�;fg#,&�|���ǌq�����'#	dm@��4��댌Q���ʖ��@01<0��,� ��25�v=g��������u��&���t�����M�z8~���w0,�i7��]���z����9��hg�m[�*�+��bZ�����S7��G�s(%YL$�acG=�2����I�K�����U��ct��� �wd��J֛aOx�=�FN�ք�<~V�PK�#�Ib����Ν>�q4�Xm���yV~FU��޷�&���hTf��ѷ�xo7�?�D]X3�D"61|%W|��V���O�:��h��`��DJ���-�E;!?��*3�8�ꁦ�������΂fL��9mf�2� �U��t�#@?�'����x)Ū�*�"]�9Pǹ�� ���m:N� �OOfq�ͳ5Nܼ�0�8�R�MF�o�M|x������ �o��	k�$��_����Z��MY6!c��g)�+-�{�[`�0�E���g4�>w%�RA� %�9�����U`g��!RV��G�=2�������L�*ړ�*�z�Z�rR�GȜY��x	_���Ӱ�0�8Y���f�5b�5y��=����ۺ�2[�������Y����8$��Xt���3Mꉹ_g��wuv ��V�^��I�f�I�tdB��Q ��uZw�����c%��4NR��4�iq5d��pඋ��?3Qu����Y��'��)<�K���9�d�$���-1lt�1��u�,�
���;������-RC�0�OSt�Kux��(1�^�2(]��3ɴ���_>��"ì��UpA�vʞVJ*٧�QC�5����	G��ן�f�W;T�l�0�I�<��=��X!�בD���9I:?A� �۟�eN*nqg���2�A@Y���� h�\�#A�.�j�K�#��GL��"&'��"�-ؽ���Wf� �F�2ԩ�Y����"����)�O#.*8�>�˾��)I�����\��i�3�o��8�R|��IY	Ϳ��^\�#	����D���ɐ�-�]��H~�%�n�7�����V�"5�Ϝ�IN�ݞ�u�(�u.�4v"��@��+p�[ C�ٍ�����M	�� �) �����7�X\,�k8I3U�B�'l8�y�W�@8����ڑ�~�Q������J�҄NB5�d�F�v��7?���(�`��8�5/Z���٭O�A���S@�DVyu��C��,���d�)EZ�;ŀ�� N�u��x-�l^�6^��p�q��H�Y�D>�t��<,g�;�kM�K�X�@W��^̂��4"Ft��!�O��t�G�&�cRA�>�V��:�)���KB\�5,+�^��\�@����r��/�1��U��5����(R�J���*����5��N�4�&x_S컂UUq��  ",�q�{��)�~׬��]�泮K�	��Ks�Yͺ�C#�6�Nְc�"�x�^�V�@f#��fU�)��0;mZ[ZL ��Xt~;{DmP�Z����м�� p��&Eh e!�I ��
.B�V�1/���8r}tw�MpHn��νt�0��j$hݑ�-Gz���5�t��&Vq��p���y�iM���MCM#��"=b��0��x���S�*��:�8}�>q�D�6T\)w)~����3��h�`���Ƞ��wM=����Cg=TƳ����uDWa?j��R����i��к��.de�z��[VmQ�J�R���
u���2���8X~G��*�y��2z�V'q?\���[K)���b<gJ�5Y
z��.�3	EcE�*�jLw;w�
�,�ym9�R�]�H7����!����"B_u�D�>=��w��Юo�Pg�GY�������də�Z��o�&���c��Dtd�d�8�f��fsBB|�@���d��ʈEO��{:|HL>��h�6W��w���bÎ>��~yh/�b��W�B�&@\t�Ief�NI�pz?�9�5.��R+Xd�
����b���Ω$rR�!�"��\e6� ��w|����������Ȝ^ܮc�q%ڝ�?)��Xi��X`�XŇ:m����;����`�FX�ѰM.��G�7PE^A����H�׃A���5)�Ǻ��t����C�v���nE)Vr
*� E�J����N"�{��>+ј�J�[G�2��_AH���Qk�Ϋ3YXLק���d̕ṁk�іБ�]��/������i��GA9UD��p8��d�Cr�&���$���ȿ���2!��s�ܾ� �1s���r�ID���T!�EW���+�Ѳ�5��@ȶ+~P�n����r5)WV����-״Esd$�A�f���ȵ�R50���4�܆-�L���d�.��G�ѱ�J� o�o�,YB�d<z��3��B��k�{g���1Ƹ Ǵ��"���p� ӗ(�	!R�Q߱���_�8)ҒƐ��.A��F��M�������<h��F:�e������!��VHMW);�=�f����-��$#���:	�m�����L��},K���|�4�wY5�"Rx+Ŏƈl1�H�j_���N�Y�V{M����ulZQ���j��NP�th�/i\4�̜��r��3�� �&�C�� ��b���iӥn̽<�(r�6�mO9�F �/]*u��h��=^2���iT���M���v0���~���:��VI�eT�
���G���tXj�T�,�*�xO���PE"��ή��~�f����M�,u�jX��I��C��H��y,���7�9p���r]�������t���;��>�(�y;�8T��2��4��pg��B��%�c5�c��@И'�׻(��,'�+�b|j��@lr�%�/���fjŞ��,�<�U�qT��9�hIRx먦~po���>GrZ���Z��� K��[�vJ�U|�}H�^���r�i;�?��6,�ʟ�|���l:G�W�G[%�y!�Jw]8�e��ݒ�d&����^�	�����ZFhR��/2N0�5i���}��l�U]��C���X͓z�`��$��ط�����Z�n9-E�z�����f�{�g������Ja��(g��B���ShO&�Ee��q�覞ֻfxج<e��ꢘU�>�0N��d.���{N��1T|�����=Y|R� Xi5e�1<�H�^�x��ѕ��y��\��ߟ�x)�-�Q%obO�x�ZL�'��-D��2res��>Pi��v��E���:-,�@����5D!��"oF��W���˷Z�Z�p`�b=N�����sT���K�r5i/���-�'Ɵ�!�\�)Ԇ���>�8���5o�,"0�b������M�G��_1o�䳲�����&�TƎ�n%'w�g�g���j��.��~�ޅM���Rr�u�U�t�Q7j�R_���՗���� Փ8�c�?K-l��ͤ'O�pQ��:�zW럅�oj��;�=�K�[��7�S<����Xi�BC�G� 2��].�)6D�T�}�ªI(Xkm\2Wu�Ǭ4���၇�y���1[<{B2���y&���i�&�f�Y�#�Ɗ�;h�@7�&b�2��P?�hOj�1����@�p�������>���fV_�?�(ZL��)�����b�5T{0O��;V���If�I篽>W�2f>u wţ>��H��G{=]�uBZ�L�|P" ���-�}��u2� �w�/g�DN�m���y��]ڊI�-K_�,t�S�E�����Cg̹?ݫ�·�*�^ܗ�?0*��)Xl�q�T<�qy ���ye͖��y�6�R:TnC�^�:������gS�b���I�%#�Z1c �2�3������ ����q7'M�2���=�ث~�XQe�|��]�K!����&�R�����O���T�CI���sYo��2�b�$�}X�'��%ȩ孉s�����HgA�7_1{Lӊ���I��ST,nB��sT��(+�Y>~���� Gn���<�/X-{�!�V^Њ!��,��k����+z�_����af�J����~'���*��=��E�����X� "�J#G��gn��C ͊F�����ޏk�S�����S��R��:^���d��HaT�������W�mh��[/&^��dwꇟh6[�^��$�r�Pe1p�!2XP�J(��q��I��U�q�,�Ƈq�_Qx�4�$Cف�s4ٸ-m� Dc<�@�6h���n��,���:%����r��o��XVؾF��9Jv?��kS����rë�� ��~��[�SfrPb��eͰ<�nv���I�A}T�jO�?���w�p��
^HE->JGRF�&��$�5�|�^���vʡ�WL���~��<t\��x�T'6{t�����n�(&�+6�L}=C��U�ih$PG�#,@�t3TׅS&�7�U$I@[�%N���= D)A+�X�kW:r��P>��^��ޟ/����c�8Z}
K8�G�����>��#;Ph5s�{�h)4���i�n����QY��8P6*���S���R�#�8-tU�G��f�U�����(��V�膼���O��6������'s06�c]F0�coe�Y��q�Y����ME���u���T�;��_��|�4a�aZ�On�o� �.1��t��8��)V�P�f9v�b���E�iٕi�Ox�m8�a7�X�.@���%�A���_FE�
?8�=��-�W���n�bC*��<bTI�=�h�Tɥ��/��-��f����b�m�9�-������Qۣ�.ӱ�N����Tl���F𧲘~�堾�3(p#'n�it9QZek� �]�;�q��݆��:��a��U�hq��QS�7����<)�7�'�x
\5����s��/=���%�R��U`�/e4��,Gv�,�?E\�lY?������da�C��|����� ��T��=s�1X�Qv68��X:�w~?�V٣�d� �n�S�?&+�v-���;�F�C�r:ؾ�2(:��Y����{�ϩų�p�@&*MR��x�F�ˀuڇx�:�*�*ր,�>?/��ߠ��: ڟ���e��hfm?m�qc. �BG`F3^
"u}:	u��ED���O��i��qt~M $�0�Gnk�8��
�@䬻�i{��]u^��
جP�J���l����K%�iVWσ�Ά���S�J�����k��$���%��h�&2LI�!����p%������[�L�r�X.@^����d��@k
^�h>A� ������)+�P{���t����Z��[��+6����ɻc>ٻ ,!^x~�1����[�����4i����.-���d�g8
~=����x��1�������61��	�~k*�2O/�d�b�)�s�.:���x�%�'��c=c ޠz{��[�rb�Uq����Ƽ����~�q���+`ǻg"�>�������U�Ŷ�ϳ�cfFjf�DN�:�N�@2�{��|��;t�/h-DA�:����圽��+Nc<�v]����d�����5F�m�O��5s�)/�&~zfuw��6<*='�����ŷ��=U����������"3�f������6�HBpk�;�3�|�r@Wb��f�.�K�N��-I�����aoİ$��+�2�����#�D�^<k<���yE�Jh�FXe�����C����r��Żq�kzWI 4�Y'���������)�Q�2�B��2��툞VH��ݏ�cVF𯁳���
�F�;~�7�W�ٺ�F��@o�k�g����OF����e�m�O��D˔��i34�Cr�z>*�E�|���~൫�9�I��Ey�eN�h�E��lizW%�x?�brT�!�k�a'�N��'���-�ɰ	�����")H`�BaiK3���(��O"�j0�t�܌|r�U>�B�NM�T���D3ſ�r�����K,R�r�� ��$��"�jq%<)��Ll�9cdB��P��	y;[��j����͟�lF2�j��i
��.��&��]�m$՜lDkձ$���2�d��j�o�砵��a�a_V�Uj!'FS���ZP̯0eQ���)TE��k�|���򗚪�`�K�O�RK���@G�;h��'�J��]�O�JI�sݞ�L��]�P�T9��lf(���=�������e�D�Q�M�s+��Ew��:��@��ZPM�O������F�\jz�B�֊�+f��K��<K4���X�4� �y�
�'�@�p����Gm�Y�}�U>V��0�0MJl-/%��i�z�mce�@�˷#m ��%SHLi�I%�d��81�	1��̲� d��nXC,��F1ڟ�Α�X"s�h�w�S����p���kO�`h3lǦ v$[Ԅ�!�J�e��!��S����2����5�]P:�3h��	f�G��&-��W��>��(ֿ헩8	���J�x،�8��t��:�E.A��}�=��1����L�U��Ν$�����I�eXݨCc��1*+�(S��.Z�b8j���ӥ����}��X�@?+ki��Q�MBBd���w7 �V�J�6$���lg����%��_&�x��O_(����@��`��-b�GV-���J�3Ⴏ(��B:޾Nrہ2R��C�V=�$�\����YC�pE���;��h���a��V�w�^���VM��D�(V3r?�t�C���\���jf���� 冑�+]��h��f�$bᴎ��~R��>���>fv6��Q�|�.&?Q������w7*�^)�i���FތBx>�z��|!9�O
f�Ɔ��$􃠕($y����b%�{U���f���|�s�/������wT�Sį�i�ZX�r������b�J���)h���;�c!u��j�=^Óσ&y�e�PY�'�i�!FM���8!�[Q8�!4?!:�\*ཀྵQ��I�}�C0�oJ˞v�(<�z�-\�)��+��u<��8�ZzJ��Э��G��(zW��,˒�I�ƴ�8��z�q���Ih~����E��Fnm�����⨎�l�F����`��K�5ϪP؟;�6o�5k�ʛC�%�DP�vY�S�x��g�WXw��ܞ>�!�%���ͷ�
U@7N�?"i��C;S�:��ݧM�K,k��<#�S���j��G�۸X�Pĕ fl:��^�]�qȨ��j���E�Nz�T-���^`�E:�p�,�6lK~7�7�0��a'K��<���z���n�+�G1�t��p�	yʁ�����!;��D�����׷��Rg�V�����J�9��F7����q�=��v�l#_���e�O�� s�5��K��KE�b�����y���9�Io��y���=Yl׮I�6��(���z=��$I-�
���W������(��ο�ZE[�,�ċ]�K�TS� 씡�S���Z���P~��EƲ�gtԝ�&�[��'�u��[<������ػΝ����W��/'��V�+�'��Κ���C=y��"&!���yv�z�g9)�aYN6T(l��}wd?�o�5#)_1���q+��6@A0�����'�d��MlN���l���jYT�\�;����"S�'�W� �������9��J�:ɓ_n]�ދ�������@Ӥ�ڽ��>^Nœ�V�5��]�DN�)e�o����.���-_^��@�h)\:\��9k�W����ecr�/010�jr���1��*G�]����p�l�#��)
������$0�n��K�4�ta�{�k?bQ�N��|e��S��cޏ��]J9�Jo�U��R���5̱���p��6�ܓ�ͤ8�L�bR5v���1�&:�v�r���첝�r� �&t������*;t^�y"�o���&��J�
��5^4���1S����b�<,l��Y�l�1�R�%<�c�`�V*�F�g�t[T���\�b�}�>���Xv���
S$�`��V��?�q���uc�G(W������7E���v�[)����|�qI9����Uy��v?2Ȳh2�r���Yg3�/ۺ�E�NM�Bs�-o�)V�k�Yւ���^q��ғ�/�֟���7���:���?��#:
�Pc>�����K�����\�4��O�zoo���J�W�4ѩ�x�����fw/���	���9c0'h�Hxl�A���Ut�Zi�2������4g���fi����z8X��p�Fd�������
���0���iكb�Jћ�cO��B�iJ9 ����FpJ��;Խc�(Ьد�NE��Ԋ

6�vY���x�\��.��0���.1#W":��+\2~��t9�Xh@,�X뒨q��
P$�)����w�N�������͟�ꌯl�7�#��5��U�����.��dc���oEȎ�P@�4�6�U����l�C�E�+���%�g'�%�E=�{�n��*ơ���B�����b�����8�Wx���;)' Ko��A���v�p��5��0|	�D;�i���41�	J�d�hd@R���=��L�Ֆ��
�����5B�u��*���-�kC�c|����<���<p�/�:�v��:���Yy����v.��-�hs4���O�#�iv�\�XSR;�yJI��(��y呙ã�1 d��b����vɌ��EN�.=���v�u°�g��X�<��~�b��<�U�Oailx0�d��݇�t�Z�Դ�|��;�U!�'�Ú��j;���/���Jf�ɾ���L '3�V�"��q�B+�nlI����=�P�`V����b\�[����9v���ɼ��k�`��3po������Q�@ �;a���a���y����+�\��<t�wĲ���6h�E�Y����G��{S �n$�	�C����Џ��(>���d��6����*-z����j�����,f�����K-[g���bvh�0�YJNU�O-�d��t��S�R�������G��,5`È�S��k�6x���.�9�%���`��i�
���0��%��ʸ��/G��!�C�°߉8�}Gp�O}0"<���� �ղ��D�� ��r���60.=�L�T?OM���|��@�=ty=�È��s��s��*D�L`M�}�"�q�;q�d
��tB�y���u�-㻨m�j���3,}�4PoXζ[���8�������\��0W�Z4_��4ͥ1�)���G�GS��>�I��L���)���r�k��Z��\��K�aў7成�`ʶ�;<�|Խ�J���D,�Q��yJ�!�-"�(���ͩ��=��v���c�_"�R��5� ��uv�H�8�c�#��7k֘;�\l�vx����9�S!��)�i���7�L���󍁘�5�ĻN�����y�,�����A�����)@��B��$?�Z��E{��$���&�/)�������N�F�W���ō^��96X�?-���l�;��YY�GK����E�R^R�W��.�!r�p1���R���R�����%��(���g�݉�?�n|4���4N�Js���h�Hsc�lo�k�,�}
i��^=D]��9O 4Z��]�����S�Jb���D�^��S��2�V�/Q����ҾG��#Q��7��Κ��1�7>���Jb-��,n�>8e(�y�]��=�z��i!�`����kl�i��.N6�^����84��\�d.�s��ڗho"���C6(�j�� 5�p�b��Uq�VA��O����r�r+/�E�����QV�M�a�[g9�7	��_�^���g�����R�L��J�
��U�R�K1��1x��)�R���R��<-�k%�b~��j�X�>�aQ�5�;Mcm!y��G �+��Jw�F�+�������am|ta�s�q�h�љ�c����(�K�{��1���9�)�Am��r��/6�-���C���փ(�5����Z�N*7���q�F��H�j�<��0��a0��65��G��_Q�ǟ�w�&߯!�
��7�����wa���"�����vt�Mc��-���2i盂Y�b7XZ^!��x�M�EI�|� Yr��L*?*��c
[6NÃܼL�j�%�U���Ѱ�
ݝn�[E?��B �E������>�����ю�b}0��͗o�udZ�?x�c�dc������~^+tBgM
�S�$�IF�*_Mq;/!g"mr�����xZ�L�&R.��|p����ayK���9wl��V��������\�>p<ޠ�6����<ą�G��%�C�k��S�E�<R�h))"AJ��C,�eL��7������p�)\�g�t�gW�Ĥ�Pe�,��t�"r��#_Y��t.rʂ����ٮ�����C�P�JwwMjqk ��p�[|v��m�I�<-_�-6aA[+4]�Q��k��1��uH��)V��u %�k^P0gV��F�Ƒ;9SqS����&��?K�����f�ԱU��`�|��W��i�;^���y�&��ډq?���KL��F<ǈ}���}��Gȋ�1��*X��&ƹ4K�q��Z�ь%�'R��Y�YAh�>�5eG��V�-�aS{��j��u���5��)�D��pz��lw)�V�#,�������k�Kp���%�~T��J�UT8a�E&<�ײ��O�	��+�/?<~�am(o.8���	E�)�|]�^!E�4U7�N��TSk��_� ט-)01�\o�Z�R=�
�y"�ڑjI�8�m��aq��kvT=5=1�4��ú���WHY�B�3�� 3c�J{%VE�_�*{��C�y�a堄���7�����+�������qd6<<�2�W�[ke���R��uJ�G���m���'���ň�w�v�k���c�1�؍�����N筕FO�7Y����Y����7�=rm"�i���'����7b�)
���|������<���{>Y;�F��Q4r�2Q^�nQ:�t��J����xV���1��_�[�U�9+t��7՜�q#���E ���ӫ��@�^��Y_34��P�v���Mv���j���W#��G�4��k�u��*��Rs/TU$�ѩQW�)��W�I�z��^Xޓ��eew�Np�=^Z�s8��&�PƖ?�[@*�r�!��/u��rtR�8u�T�L9Ȭp.���.��1o������u�=�_.g&��J�ᜫbQ�<L�P3��?-��V.��3yj��;�_�6�Yk��¬����^ (Pq఻��^�� u��Sy��<X^@!WU=�3�hߙQ�D�n�˃��Ob���uΨF���?l63B��Q5� �YB����9+����l�@CC)zP�)���6��9AlZ�]_sh�J0��sg"�%[�v@!��,�k�Ll�EQ��D�f^��_t�?!>�4��3�=����2�	wd�o��l�5�t�7��Ej�tb6��5ږ�wU�0%�#Z�
��Fo�#�I�����[O�<�g�z/BH#_�e�Mj��e�i��V�X��O�u�a{���?�E�w�!�܄aͯk�f��=5��t�O,�'L��9B�c|�),E|�D��mf��aR���E��5$X
�BC������K���W�����8g):����-�����7��L:������a���]��v���k$b�N��L+�LB��70k4�O�Ԅx���:��A}uc3˵��5:b��t�l�� ��l���0GK9��������T^xO֮��8����O��E�q��v�`m�O68��ɴR��ɐ��Z�Y��Z�@��ejIyr�vt���n�,b7k:܃�7V2��\�r��;B~��N�3�2*��R�.�%��IG�J�`Z����[n�;墩�G����nch'֊-��j�N�u�7x�%Vk�������L���B�~�(z��P��2D�r�k�^� �U��Wa��4�% .WzI��.�<�x[��.*��ઊpG�� ���U��	��"�3q+"aX���g=#��?����~��<g}bV��fp���~Cz�=����Xn|:<f�eFe��K愚����m��Z� ���Kɏ�?&"��E�!��0zz���-c,꬘!iI��H��fX�Ra*!���"��|��N����٫H�ׂ.���b��ò���T������m�.��M���h
�~���~�v�h�0
�@و T��k$��B���f�B�v���G��1|��g������x��EpPɗ� ��VK��A�p+��\;�Z��"�\�O�*��嫴d��#�<<
t%S�B���&l��ѭ�̻��$J��+���dy�W^����O���1�%^2L ZMdb_��Lnͺ5�+���_h圇���8Ww�[|�C�E,z�P�(w��b�,	��M�M1�Z����˯��+u��*�)[Җ��>��3�I�c�T1e��H�#�����` �
�x�m���pB�n����r�BW��P[�����. �`ԭ�U��گ����5X�d�XQ(<;*A�������iQ\�xo�<R@3���&Y��+2p����ۊ�|�"�l-�g��r[��a���@~���p#\nP������;X�:��(��+�ʓ��:��8F@��P��T
	�-��yŏv��������Rv�u)���}h��ދ��m.
��i�3��&�C��'�|�
�2cH&�Y�r���
���E7
.js��"tw�gO�n�:��z�ѓ�:kuj�+Yb�3��Y]�}�b)0��~�piLx|Lp4�O��&pvk�2�$��)�d|�L�[��^�-H���c"����o����`�hC�ٴ���aK�Gfex�/,B�AO��udQso%�2��uo�u6�N��ō�o��Zs�C��`ڣoJ��op^y�s錀����d�y���\��p9謹 ��]�+��7:#���ȅ�Z ۞2v�B|ox�' 49�
�3&�QOx�?����""���Ć� ~��)�<�Ӣ��ӌ4��e@44 8#�.�a3R%�b� ��a�� �?� �h�L� ��
�-��[~�_��a���B��߈��/��L�y,��K��.���6��Hd��P��r�NK��h?��;֊�h�F��U�T�uJ�-�9ץ �N%��$��t7"f?� }�b��k��AZ�Uy�����ݽ�+�ٟ�lS�'��â���<fb�Q�K��}j2'��r\��ʆ�ŷ^��1������=V#\].,���Sk{뾛|v��9#W�I���iK_{,��m9.)�I��4*mw�U}��o� ���am��A{��2O���6��A��_b�[a��x�`�>0���|XAr/Fw
K
����ϸ��@qgU�]z�#8�o���&,%�ֲ6����g�dׄ|R6��H ��36&�i�E�͕ׯ�u#G��������2�(�A����Ggjk%�G.��{���j�i�����7�h�=�P��?�����P�Wb�XͲ}� ?ޗ�T���}���/��Q�����_�y���i����~�� �l"�-�퇇��z�y:Y�k���� ���M7����'���ӡ�TmP��b9���u�)6��a���1�B�j�M2�J�&VVNyg�(�g�'�!E�&5�����D�^nӉl$Jp�/f�����ݧ��-�NT��PF�"��[�L1K��0m\��O(�'�6e�f
�tE;5 ˖�X�pZ��G/��vMpp�ʭ2�Aq����Ű����n��Q܆&]���>*��;�l\nǜVo���Z�߼{������{�%��`��<��uɞ����E�8s&Q�"�����K]?�4!�Ub�B�R��j: ��@R��;AE~=O����q�j�G{F �jW����9�v1�X�z��6~Z���L�8��^k|�`��B�l�
�e�4}˓0�~�E�p���l��Er9�x)��t���!�����F�a!�7q$�' �^Q&����m5��4��nc8�����5+�V뇐R׭y�o�~ߓ~?��P�����>�T �����!أ��(H{wܠ�J횶�: ��Wz�R!��03�!�f���g�EQ��&k�.y�Ƃ� ~�����_j�~�E�Ьέ��]�z4υ��=�\���`Q��"_������ǦH�2ɆA�N�����	|�M�^������I�$�υ�[����-	�M��+�3��F��ݹip�Vhc=�-�!�� M����:3�R+џ	i�0��Ƭ��E0p��ڭ�j�l��+B������١�M�1��Ak="�\tHb��5��J��y���M0��1���Xqإnz=�w+�B�A5ۃ�s�h�����=�ަ�<�9�6gM'{���}�Ǥ7hĜ~�i*���	l4�EU|GC��9���2�9�KAd�^�����cϽ��SUFmZ	xnw�\��,UUE�!��M3G�%l�_��C��M��vj�뎰������(�M���>2��H���5@aZ�Ixs���?z[<�P7A�(�tC�z��br�;� ��H0y	q ��^~܇�Q�c�Ah�FL�Z=��yr۩.�7��ڰH�0:z�=���^O�zK;l A�v��8>������{�����g F@�mϰ���2�r���A�'��5��AGd�@�%`:�d8?��|궦� x2Ìo)�:�h_f���o�Z(�ߓ��gq�ɓG�Z��+@$�p$䦊�&��i�Ac���b5)�缅��{o�"W��p��G�l���G���Na��w�����s(U�[���)�lȝ1�Ϩ]��/�`�\T
T��`̻/}�&x~J_1?}�8oy�mis;�Ky�l�4�J��4�O,a�T��p��jop�6Q��v_Cv��$?�l;���k��z���ܩ��fBq�U{��X׆��Ŷ�Afh+��)#�-�3�K�7���	�~a~�{�����>��T�)�yGQcb纹4�/:u*<��8ݠ�M���_�(:u��|��$ø*�;s������fK�pK��Kl����;���ωG��7أp�=�Qv>�7�^s~� �|��"����@YBEվ(h�ꪽNInsʻ�TU��'m�%N)}߀G�PG�@��d-A�0y?��/��M������pzzf����2k��j7(f�:�h����������Ö�n�J7*[+�h9��Ӡaɏ�
�ɺ��%�����墟��S�� �_��#�M�3��x��+)������L���o��i��'yT�{��&+�{Μ�����t�ς{b�_�5!`��T�:V�@L|E_h����"m
L�)�\�X���
�׼�$��D"����a��yu误k58y��ɷ0��$r�S]�٩�J�1EUY��{�I�gg����]>����z���[�;F��9�(%������и��8΃�����W�d����H����W�1C-@��6��n�/
cU��4cȅ�L/e�D����T��-�63��	жE�V��X`g�r9KJlq��@d�����گ~_��F���MZW5K��.y��9���^]�NE� I�;M����h���W&A�C� ���:�V̺	ZT&�Ʃ��2TM���To?�O��0��Ҫ����q��8��S�'�嫇�_@�Dylȩ�P�E�]��6t\�F7�B������x�"��8lN�����<2���.'H�ng�#��D�F��Ks�]u.{�|
&��n��H(W��6J��;�E\�Qj�Ŏ"���s1(���� ����VnK��U#9/�Ǭ2���˴�G��և�\-�"�x8e�c#���r	*�F�=�CMG�n���У	���-�k��q͘!�[wZl���X 8��W'E�w�8n�������A�'a�"����NB��16#����U܂�۪��H�
��]|(�TH^�KL�"X���	�`��uǧ����<�>�ns_E��[�&�^.��:25U��.�5��Oґ��m�Հ!�I�(
��#(O�6m����DD�7~hADx�iX%X5еham��ذ�ң����yX�\{Ȟ���U�*�3��bWmg]�r��OKzĒ��|o���N����X?#g�nC�t�z��� ���h�۲R���qu����k��Vh�> �����9�L}�n_�t͹� fCXO���́�N�I5pƻ�^�z�W�D��͟��� j�mU2�<0���YRy�.ܑ���^��8S�)�=e0��/(Jw���?dއa�Xp��BB�L���<�O"�ۚSHO ��.����ќE![��n��-�]K��f���~@���x�1]6���=+<�>^������U9d	q}����C��z�z�%�C�.��f��A��K�E��S�{���l���~9I��T�n�3�ޕSY�D�����)I*^\(E�C[,��Np`��G�߁2�}$\���H��o_��ˌ$�H��v\����� }u�
3?gU��Bj������.L|G�����@S�mdǃ��ؕ����젎��Z��>v�P�8�w��\�䂋Ľpj+,��p���EQ0f�|�8�R�L���}�@���a�"���}(挀Q�������$��p0L��͑la;물�N=�o�5��"��"'d]�Vx���k7¬ �?#�$]��)K��R��PMڈ�|EV���+�84XŪ�b��p���3��MJ�I�b��-��,=a���lF�Sם�,'���[�U/1{�J����:���4U�Е+:�g�����矃���,f=��O�e.���.��Y�3ca_ŭQ3D��4d�g����յ�$���C�n�	Id���t���h���~O���6K�#�(V��D����@D�ۋ�%�΅ю�A�<k�g���G��f���r'-����.�+�!=�p)=)�>��g�� n�/�Q��|��w��b�U"���B�2݈�����,�ΎQ-�K	��z�cWl�����}�믐��8��zY�{X������N���߬W���%��(4AS~�:~�E����v>������I�:AI�j� �2���V8Â��n�˝���A��Kb�"C+���Q(��l�� ��o�?����fО��%�����\��k�I��� ��Kّ0���*���Ţ���~R��c�\���kcv~{�6��Jn�fV[�R��N���5V|(�P���N�"^"�&�ɱ�a}ٰ�����d� ��90z09��m�`w|�{_2Gu�#����P7�˛����Z'�=j#G��;+|"�Y5���� �O�?�����.�\]���Y2�ڃ�䂣m�1�?J_����n��OP7�1�w�z�EEM�۰e��5���{�[�_%w�U����E]6�&��g���|�NU�!|�J�����Q��k~�T���8�M���hJ�B�'����Ҭ���-����%J�ewB(ca�PZ���=��z���.����{ńLF6���D�'���2�1KӾ5	b�6�eBKx�!"`UO7)?)?���Iz� �ԉ$�>���
G�2�[T��x*Q�pު`M���o'-���[���8w��£���|�����^c0��(t���M�x�3v�b�8ĭ
E�(s�����1֟U0#j�'"CH���w78�
h��(���rU%Ƭ�k��n0�����g��0o<�'���1zy��^ٍ�:����,	��n�%��D-��e[�)��eQGp��;(�z$|>�,y��	c%��>u�}��waO�D��	_�_�޿E/A����̬��R��"4r�s��O�G��R�1V�J%��r�3Xv5頑;츬��l�"��E�2g�����Dd�0S���7��rc^�\Ȫ��n|}W��}
��a��Q��SeT&d#��W�	u�m���8�:�>7�B)^���/$�g����X��wdK**���M����v�i���r�[�h��} F������
G ڨ]eb!�$�����'�\��16a��]C��5.)-�B��E"�$sZ�'����[bt>��=�5~�'��l6*d��% ��A-�mٿ~�dN/��:���v	�b��ch����.�i�^o:{�bpw��0���j��Y&�Ӗ,���:�ag7'pO*:tΫ	��MY�ݔ����1
6� ��t0�3i�1���˒i�<]{�,]�[������@"J%:��SY�Y�ɟm�_ ��MG.������rLUIO�}@5��û<�;�:����7'	Z�#5��4'�r����\�Q� �!b`����j�&t���%aj�J�r;�c�Rc�Z���1��^�t�/V���;��+���#���W����.�QF["F��]��G�^���h��_>�;���T�Icd�������#@�\%�%��)�!p�o�c�
�j�ba�d�����N�7��K�v�w-w�=�
�Z��z�mp@�G��$I�.�YPy�6y��u�5_�|�����)��4)�
�j}ɣG0�^�kXA�\�	>�����&ʌeh��
����}�o��ܐ�SR޹�zS�H_$!�?�r�qۯ�YGc�X��sV=������ݧ��:�Y�æm�(Eqd}+C���4�MD��FGn��i�fFZ���⧣����N@�O����0L� ���k��o�$7�޺�$�ը��l"��F�6��k�z5���]�u�a蠟��{�)3�;��Y�9b:�Gsb�#�>}J���W6] ZA���uձ�P�lAQO? �k�͜�e?p�3��rh��ɯ�V�
���\34r@%������<�xN��18c@��[��[�M Q�|��z��iֺ���[�2���FkU����əT}{�������XP��l���2�s�q��`Ԟ�~��Lo�>/��?H��N� `0GQ�n�g/�C�Q�#y���z�h͠lE�i������1��j�\9S&D�Nb�[�只��lQ�\A����g?î�)x��=B��y�;!Ņ�#i<L��T�Q���iZ�N�2��e]�m3~��Ok�����k��1�h�.S^�H��L�h��5_x�|���0��G�b:�0�N���|p��
�H�h�t�/��إ�j5�W�)4�!9�n5즢N�W���<�]=�����.=�kK}Zؼvn6n�씎B#֞~s3�j��N\���}��#1�#�VCL�il~S��+"��И�J�z)�Ze .�i�Ia��+|)�0C��*�d���ݒ��q]����2vV�_��RvP���A�厽.����������U�#Hs1��D ��
�ofX���@6�!͜>RI���msj�������=��|�<���P7�Go�*g��i���X,E�K:��z��m�ƅ�Ԡ�׍�(2�����"Q�������zΓ�в;ϙ�C��x(�r�;�N�Dk�!�ȶ��<�>:�F{.Cy����yǕA�۞+s=֖����.v�~vI�ƥ�,�C�(� �}�`/��KC��A	��'��9�m��M���Eɒ(~����<����w�v�7��PޙC��)���7U�9ρ9 ���쀑.	u���� ߒ_�n-�BI5l�t%�e���y�9~�(*���4
�1J�3��T�`?�q�@���rqm}�� Ԛ�46�������>�9"߫�y!�yy�u7v�ѐ����a�?�ן����/ȕ��1#D�Q(���Ƅ�U��hͣ���|2�6I�މ	+���a����|������O��Wf��D�^��P�W&����n8%��>'~�1��>�wnD��_�_Y�(r��<DXZ�d�}����z��(�H�D|����������;�PlR�F�0Asj�) ������DX�����b�_F�m!yg�������������KP�[��fy�9AR�G�)��R�փ�%oG2�J@�� �.(�Ƴצ[ypI��j�x�DG�av��t�.�"�f�A7�kj �y�W�������	r����4�gl�l[p�Y��td���)jg�8N����Ҝ�D��vn����V��/�ϥl��^{�>�\��?��ur���,[�٩@��M^��fw�J�k�@ŗb��*�DAe��1�lv�|�&�T�� �/$�MN�H��+�G���3$T'��ɋM�{���M.ױ��%6E��~> �J��\rb^ϫ�4F���>X��?b�Z-8�&���]Yy���y��X��U��
�3����g�P��nCDp�J������Y	�M�;~"|����Vk�z�������0]d?��w�0hlk�^���[�6>�Y4D3�)��ԥ��Z=QOM�~�QPTN�
1�,��G)b�y����� 8�`\]̄���	�#�?W�o"%|�2��/��5�P�������y����گD�g>�zq0sH�0�������9�/ל˚�M̊�'�i�4�z���b�y+rO[�s&�{�w�&�=ܘ�*m�Oڴv��3�a����ۮ����=n�2��ﱎP���W�TG_������T�k�x�XC��@����'"jbu�R=���L��~�^hKU'���BI{R��'�W����m��w���tG媐�U����+���c]��1S���t��-�\��V6B��d��LS�v�s�N���*��:��$S5�c�.���D��O� ���E���%���⎣�x%؊�xl��L�G2�63Jh4sj��{���G�k}�'!�� ��:��pMb�A�9{|�֏�K�]Ѫ����Mg��b�~���6��g�B%~��E��j�m��g��#�Y���بF֓��X8�S�3�l�.���w_�/Y�%��3�v� t*�v>%����H�E�^�34���P�ʨ�X��&�Y��I�����v��Ӥp�f��V@�p��Ji��N@�j����c�;�1��a:�	�G[�c�d�5b�ι���SE�YgxQ��2���dC���]Wu�?$�| a����쐧�G�{����f>3;��~1�[�yMN�V)m��$(cyw_?:DU/��%���^���]7X"�%��Di�w�|Ǥ�]�/u�ƈ�bd���� y��
F�xU�4#�Q���rU�� )l����S�ˮ�<o�� �Xأ�DZ*Ď��=��Gi�t(5:t)\i1����mݱ(������Z�;��SK�oN0��7>1_U�]��,����ʺߚ�
��nѨuۆ|���C�հ0�К�,d�����x�<���z�l7m*d�˿�\��F*��>�Ak���wI�[l�Ƥնl��[у�?���:��U_�L�׬�f�W̏r�Z�$S���<�q�&�r�y���;��E����JtI0��#�x����X&�����m[W&��`��"��0}�.��4��qp���g�#bG'��b,�o�e���Gɪ�rH_��("���^+�a�� '_Y��D]�֚�����������S��Ië��zk:���S�'�����%)X�(��M�ī[?uQQM*�<����u2�_#�d~յ�݈���\�A����IWUQw�ۯ��|��~�he��Q��H�έ������Q[����0LF���/r�Sj����6S�\?Q	��)=-Lܿ
��A�J!��w�T�z�l��S����y��=�U̸�֨�8'���Cb5O�7O��'�5Gs���|�[���i�7��� ҭ�V�/w����t��VS�-pg�
���4H`�rs�{a���'j�=H{^!�z��c"Ok~��c��Jm��iMAK���8��~�(�SBnu{W��	ܣ���A��1R�ź���yQ�y^��k-o|����Yt��7Y��iU�k����@O��kҠ��ZP}m�~����?p�B65�y���#P0,�R�=��W0��D�X:��H�`G�/q_ՉUٍ���Ɨ̀]T�>�s�)���A~lJJ+���B��tV��D^�D�,�d�%�K+g��m�bػ(���A�5�>,��MP�&|����V�V���Uj˼},Ц�0j�>�8=ᝤj�I���̝,7��#�� ?h� �Fk��������~݆ǽ7��K�ğ�d�؊1���,��ɉ)�gĄV�i��KMq��7(���jrIP��%�$�k��W�ȥL�B��ۇ��2MVN�q�+^�!iҳ�[���y��nT�"�&@�K}����j׽��F�/\�%�c���s��|����i����ź>����f�-�6\����(oK�hƐ�P�>�W5�q�r,�D%<��7�����4)��^��҂��,G�D��j�0�ׂ�`68�gds�x4t��;n�@o'�e*QN5���{U���b �q6�5y�i���-}���e���D��]~-K.�SY
�D�i]��N9#�����=�P�@��ˆ2?Y	��)�uhB���5�>h����x�qd�k��{���?�rr�}�L�ll�u|�2Z�0�爃�<�4���ĶN<�}��D���e�RK��A5#̆�"��Z��nt����z�vɴ=7�HÏ���=31�A9ܰ��|���5P,���`	x����$)��=)ab�llb�PL�ant�k��6I>���2�O}�6�xn�:6Jt
�d���[ާ8���u(]*h��舽ͳ�|Sl�/�T�V�k=-\?FJ����Ƨ�9G�pO��:go��FظY���f�i	9/o��ݷ�
�}ݛ�{\�P��7���^��A4t#�����=�ZT�B-�������<�9�t��&�i���s}��w�ź�Ia�q��7���H�{�����:����^'���ㅪ�M�Bi�ZwD�yf�E�!}�p�
4�Gc7���|v벖��c4{�myzN�v)��X3\�[��/��=�,�b���G����e�ظ������q����M+ζնFW�Q��"�'��A��{&�<t��5t�����d��Rb��p;����8�ܞg�ʺ�L�]9JegL�e;N�N����7�����S�Ѭ���n}��>SO�am���8�����r�ʏ�ZcV9��!	�ȓ��Bi5β���c3欢=�Y�Q5J1��c��EW]���{�q\['���_����X�]HG���-Z�6�X� d��j�Z�HI:��I}m�uH��ڲJ�=����{�b�}���Pn~���I�j����
�,�MZi��>��������2s�u�ͮaj�=����u�'mƨ�z���z�^��B� �����O hcK	
A��lMP�A�Gp��پ>b�Qca
�gH�o���(����:�Aw��\ڠ������|��0HD�'�B(��)�i	��Ț~*��U��u��5|�-���K���RC=��u4H��r]M@���hc��S37�?W>F.k�,�k�,��`�n~Cq���[�.�HT"�=�����_�+�Ӧ��ãB1E�dl��f�x����K�����mw���,~��KE��
4���EQ�s��]΄O�� 9��?n��9���Q��Ʈ5~��F�_K��E2@�$��e�X��q�,������:`��=�&5`����l ���ƶ<�u�#q�w�^17c~�QTG;>Ez� �Y�K�����h_����N�W^�p�MAW;�c�X2�2�iH���KO:���{�n��$��iM����t޴,Ox���߾�[@6Ш-�{�a�6)�-��q��z��p�3=���õa��+?���Y����u�`GY7=��P)xW�9T	�C�i�v0�0��Xlӽ��f����s-/\ˁ�c�-ɱ����&��6wըR��'�*�{���6r�q�@?���:O �M��-6�H����a�Z��ք����̥�������������b\��3`�m���q�u�v��^�LZf�'��k`�,$&ˇ�~D�����(Lk�� H�Ǧ���Va��3;�N�*Wn��ixf�1��
�<����x:�O0�k0������j�5�\����o����k.ܛGF�9�~��W{V$D�F��õ�gK&��/����ܣ�qf@��-��V�>��iG�i�l��Z��ヮsw���b!��y'J�:,��O���"��t?3�VGk�+J��M�*�3V�sɜ(
�d�`���Z3��}Y���R1sbx��Ͷ�,T�誯k�2�ŅzѮ�w/��4}�}�ڇbDWr�����.F}�G�1g.Jf������y��Bޅ;sC�;�z��v?�!��p�� ����6`ep�D�JW�R`��m���b����2�&��I~r�MxОx�������s�P��;o=j�������ݳLUe{��g1�ş_����,�}�^ͦj����h>'���C�~z׳��hg�1��6��P>*�}��CP��uI�;�s�ݙ�ǿ���c���e��ʊF��Hcx��l�&����m��SJ ���;1#f����w'�vKtF/,S�jq�:b�s����G��té�i�����8�Ӹ(M}�u�ߖ��LҤ�Ы�SF&*�!^@��U�ԝ�
�m��_L�'r���Y����%��r"Y�b�Z ��Қ���L/�1i<��Ո �[�p�I�v	�
�FW�����u�O�,J����B+)�<��ӎ(F�J����m�d�������U���2+��>���[���T� %���I[�o�&�Z��P���v�A�	+���QL�~��R)S�q���{A@�c@N��ǋ�k�%Z�q2%%m	o8��}Xo?n
��\�ܱ@$T]��x >tq`a19Ku��j9�-9pkg$H���pΜs%d"~�;J����D`ׂ�[���j�Р&��|��.0Îy�j��SəX��0��=5�ş��?;��dI{];�W�au]m�dhn��g��KFX�x�<����~�C��z����5����R�Ö��"FO��'��%������'4<��S ���|���>��?PL�ȃ��BO�㱁�M>p"0�ϓ�p�NW���WL�'� ܚ��܂�P�	n�㙝���;U�ȝY���$����g����M����wO�9K1;c��v�6���=�}V0X$�5��Q�A�nсG)Ŏ	������=��p=q���a���%�v^��6��K����yӢ����@q�_/�go�\���0ѹ�T{2��m��}n ��W��i�XG7�z��P�>�È��;!���v]�ERR|M.Z�ed��>��A�E%\4�Jԝ\�t+��RA�	�:]n>69]48��2�J�ĭy�^]��\ϑUW�ʎT����y$�6&�f��j��sW6�[V��!5�<LD?��ܒ�{���_jcw��eߚ��g8��l�9��1A@(6�m	�`Nw��Ο��nN3wF1o�I�>}S��DK��X�s�g���h2�j^M<�K�V�MLc��������W�bVV��9U���]2����g���>{(����?���_� �z�
:��u���Pm|}�9�F���@k0��u���@���qT� �c�	���Έ~I�bN��t��ق"1�� ��@X��>o�>Q�~ؓ�mfq�?�\u����ql���Fx*�E4$Jg���Χ�y�;�@�k�n=ϻ^Թ+���[�7T�y�H�i�3��A���������~n���ӗ{�(q��E� ��)�(6�B��e_2X	�*�(?eb��p���L	W��@��Yl+�	�RlU����a��0!�`-�ŭ��
r�K�r��{�Ш2��Z�Yh�x��M�����s����������Q��=���e�dH���~zeM�����B5�3����\�+*��b�������'������:ؼ�\��W��C#�.O��QŜ+I�"؝�W�(�� �A�y<�.��b����p���څ�La��O�����&$<�M�"�ESa)�� ��][�S>�>e:�����TA�3a�����H)����X���C>�H��v����s-r��+I�Ѻi��B�7U�}y�U�iXZ#� �gM�w0����ix�b9��2ҝ�E��'I�Ĥb��m���4�;����h����*p�����s���P�H���0����t��Kk��m�O���v���SzU�R�z�MN�H1���A���E��3�'���˯|�*����5�Of\�[I�\3�?x<�wT�`��<IwP�U�o��BG^���?DX��9')���x�x��������z�g����<�c-��e�HF�+�!��r�����!������a8\K��u���w��#L�9�Q1r71xx漵��2�(��l#�9����PƉnذ�_$��9f���i$W�.��. ����J����vX���#ə�J]�����K��7[.Ez��V��F���3������>�� 0���5a��j�»nf� |O�&��?0�X������1wQWXNB�`@�{5��\n.Y��ශ����ٹh������c�G!��ӝ�+���{����r?TET0�1�a��O���n�q๡�N������G����T�N�(;�F�	[p�H�a��޸n�eE�ah_���N�`�Ul��V l�_���㚵������Q�V���4$Q�NpD��o�W-�k�p�C�~�@*����4�?I���=�.��Su!v�W�� �@6�$�����u`����DoUM�p�e	�����-)��i��6t��q�����ˠ�i:��_}ksSvV�6	ܰ�e��t����a*�����hV>�U�{� X�-�IT�� i�3�(�Z˚�6C�U� s���'%�+-'&�=�q
��d�7DZ���p��zG�h�+"wLN�n���"T�M�]M���6
t��З �����n���P6�J�7��I��Tp�>���nl0��߯l ��
"q�P����K�p�4Z���_K=�p�<�G5���)T���R���=�r���+�2?�(�(���o�	xm R<�� ZҬ�'��wI����0U��\�)�T{0z��7��o������8%��T}��~:���f"ޙN�YG7A�v<��N�Rcv�����uOE�{t���R�>E��su�|35,I�[
��.��иҡq�S��5;(�d�"�C��j<�7V�V�:��hli7	Ōv5
��=V	B��J���]����E���)P���Z2Z�����3�xc9��C��670ie�q3.-RH�h����lƼ�uB���@j�������M�B��yv�ʴ�čL��}6���W�a�
]�D��EN�R���|�ܡ�N"����ǿ �6g��{��-Fg�uB��OHU̲2��R@߅2���׽���=6��g�f���&��R�"(rAh�@��"�*�s�}YQ�֡�����S�Twh��u�H�0-z�� J`X�L��}D��ym��5S�����tr�bj(:��c�"��M� ��i�;�6/�u~�|~���D7Na�2%���� �[KS�.��.���՞^�NY|��B�����_9m2�1X,�}��Y���1㘐�`g���wi�=�BNj���i��KLф��;B�@�q��_��~՝\n�\Y�y��6�NI>��+T��;�{×<�{vX�C�Z=��e�n�Q�݄_Լ��[vi5�in6���օ�0����#�'۪2&=�%�l�A�O�����uH_m1�e���b'�JJ�[�P��Qs���l5�(&� b��H����c~"=U2#{qӻ\���ܷ^�F<�OK�+'��7���3�}��p{���<n�o9�?���mdݝ�c��Wd��UTRM02����5��B�~����V9)CK  � ����� ~��seǻ��-�%�>����4�a��ti�eg��6�����N ��G��Rfc}���ݱ��Ju�ﶜ��*1Ź)z�z�����J����Mo}5�=�H�ȥ���Y�JȜ�D�r'�C9"���i�"Ծ]���G��>ew�.˙�M���W� ̘< Wm����Ob�!N�͇Q�i#+�Oy�ǐ���d;�-�2bܝjh�|Wƪ�L�'A�C}�%QI�ԅs�RA�@��_�����{���ǒ�g-EE��1sڋ@a������^04�y;˜�}�!>�����~�Q3$$L`�H`��xׄϛ��c��i�c�; g��[�-�غ�J�ӢK� ��R���>�)�_�VD�\/i\'�&�2mz�r�=4�:k�&7����Ue���!�_9Bc���m w��V���?f� c��H��*VE����6\�k;�lP`L�t�M}s�Vß����
HP�c�����۾s���w�,���,��I�8���-�}+�ăX�L7�Y�������QS͜}fu�\��G�6"��
z�e�d)g�C�B6j3C���%=]�XILA_�� �Q�?��+Z�W��fa����u�=�#[�I�e���)��{�@���N�#� ۞�|�&6/Z
�����ե3Λ
�6Қ���0)���	��"(��� �ar<V�E �/+8k����/��MT�(�$0�C�^�nīK�4�go>F$�\�O��&����r�!,�^��h�kP�nUa�w9a�Ë���Z�#�P8ǭ�����3���p�o�&��R���i���a��J 
�I˟5��rRu<tg��k��<��\F�E[2:#�/�~��nΨ/��zk�{���5�"�Ѿf?Lwic�����������cJ���B��B�
��=�0����¥����o����#�Ȃ00k=I�	������r�z*�[އ×������+eܨ���ӷ;6�2���/T:�����Ř��������i]0�屳\ǳ�F��G��#��E�U���Tq=V�war�bJb�.��u��[=3�*^�)&R�e8�e���y=�Πm��/|��{�@j�蕈�5��r�����tҊr��'��c�Q�
"�����a}���a[U���� +�]�O>�A�\ñ���͗	�B�-�V^//��\���D@"�Vt'��lُ ��ZLs�3�OP������|sAe���f-%o��D��Q���$�h��' ���_
��H��,	��(c�bw=�)��S턢?����q����!�(�&(�}�����n�T�[3=Y}U,�4�\ڝ_yRqP����Y����� �M��Bd��C)*zu�M���
\�_u��UpMZ��a�-I*��pv��4Uz������'8�6��Ɛ���n��=����a�� է�s)
���⟡\�9�GL7���QM"L`�_݁+���0��? d�ì����Fzh19􂕂0:!�6�y$�F�^Sz��#U/�ϠC�kǹg�B��x�;/�~�V�A��_*4\2� �`��0��Eۚm(lQ�O�#�7*�{��E�(����	��Ϡh�*�)c$#�� ��-��<KW�ĬeMvld�񤕦�+)���U�j���ɴB��~��S�p���L��ӯQ=�,�v�p�FUI2&��c��?��J{�\��}/�>����N�{���,#W;�[��Esf�j�?+�#�W�v��A-+k,��2Z�����u�<(-a\U�#�߾~�@��%C�/������Xx�.[S���E�m	�OH�k��dm����o�wk`ぉB.i���O�.�Q�k�5�.X�GÂ˙6�2����Qe�t�����D���9�k��E�$LyuX7�����. T����E�O�r�)! �`Ȟ���u��C����`���}Ƽ�U6�������@��~�/�l�d�	1J)Ur��!�!��ىr*q��k��]Fc1UґO�=յ��\��4�������<q�f��PJ����,Q����o�Tm��D�G��Z�Lٕ��{��`�li�œx��m3��I�!A$JP8��\�f=%�A�w���5��cQ7m�fOb��bᓟv�f
���,|����ơq�}��jb�(�]��~'O)�ݡA������\���1}W0�o��\���uu��6���l]��ޒ	�UŚۊ�V7n:2���db�
p2��:g��6��y�(&�)W���^���2�d��Md�����Q��6ҏYE^Fu#r���j�+�!F�}Q�D0�K��<!�v�\�O��xV�&S�v�/qc�mT��Y�B��W�2 �gI��re#]�-�|���z&�&��ݫf"����ځ�1@��8�e�M+��Z�I�u��0���r47|ƪ~~���a��n�&���
`��'-����Č2�2�9`�]2&Ϧ ��7l�		A'#��<��Tr�	���h�"\�"�weLm6+P�	�~�Wo��l�V��8)V��6?m>"O�#��ga���"�y*z`M]%_>s�h���f�պ��A�*��;�L �w����,ć����>�L��յʆ��)B���߱���M�ѷ>
?���?\r�+:�.:{a��7ڳwP�M"$e��*�X��`I�M�>Tb�N�Fۅ���Pq� �ph�q� ���S��O�1_�����W�o	U���`U�o�Tp�,�F��3Q�i���z٦��"d��:���t��":Cy�v�%O���݌�Z�nC�&Х �6�k�5B4Wn�ۗ��`���8���A:W�y�!g!� �=m,�@�E����"���W�N�Bg,^�	
E�]��I���G
"kPO�q�|]fz��;	��A��^��ω���aI,�D���C=�����gMZ���O Υ�	�49�f���%+��K�rm鹏)0��?XAj�Z���k_ 0����5��D�ˇ]�q#��������>,�gRs�*U�y���:���|L�}���^v0��;aWI@D,�ۣN-o(��]"�0s�Y5���g��hN��ٙ&R^L��a����w��c>2:6�#�,@�a�R����[���:t|z�9�k#k�@��3yd�BIe��{yW������}pU��]�$�� 4*Ʌᦖ%	œ+c� !Ԉwa*�$[�u�J��2j�H���ߵcL���b�/�����a���S�Z(������ڙ�\H�G�牲D�`��-�d:���ߚ��%GN�D�����$��Zl����#Ƙ�h��ƽ�|���B�Rl�H�$�S*�[a��FP�I[P��ႊH�q2R�B���ٯ���C.�Sm-�-���҅�_L
?�e�żV·OW�&7`���`��h�jjLg3�s��Үt(��@�#�'�w�� ��~�������0Y�K`_)�иV렫0z��'�@�Q{顠�`&+�@��ׇ�/�%�Eݮ�5Cɔ]��v�1��>�	˻�n�?mH5��
����1-���^:��|R]D�64~1�q~<e��l���E�P�<]�O��_
���VY3+|I���#��h��[��NC3��m���V�B|��e�+����i 	�#8��'^���n���L���ǜX� ��ղ�I4K��Z�_m�����{A-�6>�������T$��as{3Qf(mcZ0���GR�=C��7�M7\6؆Dd:M�A�4�Y��N9�F��tt(� ��_�=ek:�.�A^��WhU�z�"�n�s���p�L�ܖqSCG�7����H�e��բ��D�z$�(ډ&C��P3ޱ�Lݺ�[֨��à�7-�.P�EZ��6�>�P�	,��*�$>)HD�o��d��k��5�n �w�U~0ـ���l��g�T �tvm��<�6���c
 �%�"P�C��k����������nD���%j̉{��	[��P� ����5�_п�u�a��%��g��lB� 1'���'��ּ�]rI��G�
l�0��ᗫ�� `�K�<G.��4��������'�>j�o�G��l���%Rg�� L����sY����W{��\�n$7iM̧�̭�
��6��t�����=���u�l�Thb��L^<��(䢶�҂�ϫ�tN�������?�3*����~��N:4x�N95�r�4|}�X�'�x*R�����'y��æh6��i����=]so��� _`�ߓ���k]����Н4]��6RW0�����=n�]M(5�.��H?"o�@���������>��b++��[��mn����*'��p�� Ea�_��"�Iê�y�]�Ҝ���Y���<��M4��o�L��c���_�,�ߊ5= ��-���3�0,�<��ۀ�p<<�7u,R�žI5��N��k���GIT
/������7�(�T�%qS��j6/&#���V�x��=�u-yi�t�|��� �{͚vg�Q�=�D7�9&�+����o�y#. �>�c�|lΊb)�J즙 
�<���3iv�vգN��$q4�jlލ�=ԁt3ם/n�a��_>O2���8���%!q�.�t/E�ZƉ�#���#ӳ�,��	������eH��I*���l'S���#���Q�Z��is�{f|RE�-Y�Es�_IQR��]Dh?��_�i.����'���I��x��{I8Z-�,����?��P� ����%&,�_)�6�k<�P49@�xѺH
 e�DǍU!�a4��o�o��^��<S&��f��h�k�Զ�������6,��ofp��m�-�Y���<8F�$ֈGt�8&�{s��AV�犸3���򳌱�)Sm�^�$�i���r�G�wQ�>&���f,`�����g~lS%����;���XB��3
8����R|��O�}؆S��s�lV�.�֏)ɬ�N�����J�B���a�j�30$���O;��ՑP�R�����ׁ�xw`$) ֗��o�u��֩N��*9�0L�h�ҷxM24�s�$��l�M5,���u"u���Ϛ�����\�gΣݸ ɟtpI�jH�>j�o����`@���GI ^he���9s�@7٠�-.�b[A��1�]$�`�@D2��{�p<��)�H�G��4e+����,4 &[���|?_1kڲ��f��Y$e����X����d��
4���r�`�c07L�m��ͩ"#w��r�1n����E��&��RU�;���v}�}����}JRu|H���-2�kYf����s��.�(~E������>�� �b��@v�
V0�с)��p10��ZE���rb���q'M����� �A)~�zIq�I��LռƸ��c'�~�zBFE�e�q�Z��͛��ԇ�z�����FF��d�n�P^	Ű�=�=C�	��(�r�=�^-G�b_*��
Zy��J<j3²Q�ͪ0��v	m-����%�>�}�z�� *�Q��V��h����Ó�����p'��|�L��Jv��,k�	F�70�R��T��
v�
3���7;�ى:G��k�9k=����զ#*EW�6�w��e5�U�A�Մa�ke� ʑARsEs�r@�lX�WhY%����#�ʏF�A��Eg��Dj:��7~��Sw�`��&>w$=������y6�0�#�GF�}Q�9R�6��V⪇B���MؿJ���tB�|Ig��V}3�bv1Z�]>�&�0d͆��o�0���F�}��K@CKT��S96���ס��R�)IGe������\�!˭�5�a��������"�,n��3ĵ%4!���ve�d(�N������l>����#�`2�RK���#K��5&rn,q���Ec���5�����(ƶ�_��pt7�G����hc�ۘ���M?��vC!!A �=���u@�y��VA�wCB�e�R��p�4x,8��'AS\;ϫ��.o�[���b�mE����{�WUNq/�e5��L��5�Ǧk�9����7T��R�I�'��+���U��/R�&D�f�4��v��HD︔`+�s�_
F�b�yX�=	�p�L��G�Wlh��g��w�j��80B�f(���u��z ^��.��7��������2�4k@|1�G�~�ޣ�~�$.h�ZD�2�`'����wtj?xa�q��ܑԞ$�A�B�������eF<̴Z�b�iHĻ���,��6g��<�4Z�>}�z!�=�ur�e��>��{٦� �� �YL]wʠW�0p�N]P�6���J�6v�a�"�y4)i��{�b�M�!mB�X-��5�:�Â3��7ʅ�B����[g(�����R�d�{��B���!�m JT' 
����
�:�����I��a��#���Ã�쎰�0�������S�,�c��>�J�]��	���ҙU?��m��!��vvgm
�R��c��l��c�3-��*~+�_� Bc�c"C�K"�7��#�(&���`��j{�T�fP,��p"3�~���X5ml� �h]�wRr#
�K%��$����Z���˃�8U`�AY`��*!8_B����H-���53#�T�� �[�(�A(h|&%`��*�C���ɹl�H(�8��&��g�'���Q@��Ǡ9��R��}���Q�ts�V`�ƛ��^
�> ����J�qz�f2V+Ҝ���;�aca����ߜE� Ƞ���/��������"
��a���jo#�O_9t�T�Q{�.G۠�V$�=|oB��eVE�ҧ�Dzb>�J_�{�Fz��
���?��pe~;�M0�C�P����Y�.v�Ӽ!EU��H| ��2	hT��n�D0���H���J���� ��a��[�����%�L� ���fo�@�.J�H��+������!E46��-���oʫ���s����=�~H��n�s3�]N�tOO���az��}��S~W�c!L(�Dtp��ȭW<���-v?L6	���7ACQ׺6��(;T�k$�j�ek3��,�x�	�Z���N^��9����Xڧ���i�g��#�^�qr4m�7:#��^�68�����>5�]C�����4(8�[��x97�&pxB�8o�]4�;|P4��+������*��,�?&�z��B�R���zG�9t߸�H��F�J6j���=3܍7B���1qt���)�Q2�i	nN?�$
��������OO��̞�%�bE:��}�v�]m�b��1�,Q��9�r�. �Y�z� �/������s�3��l�Wa�bA�m��y���&����Y�ࠧ</9�;i��Pb�0-�̎�"�M]a�?2f��SA�J�;�Q ��_������HS_�ݳqVe@ϯ����V[#�����\�����Po��2;�*'��422%��F]�GU/��W�*k�M^
�a��8�򙊧S}uW���*��ibZ5��O߿?ˉdY�(��������7��<	B&{)�F��{�	�en��?�����BMQ�	T��%t�Z��ʙ�����I<ﹺ����c�&R8�<rP�f��մ�ƭ���˂����ԃe0���+������Ŏc4眖'�Ms�f�����E&��u|f��2�������� ���vی�7�L �BK<7ؖ��K�&2*�b]�f��4�u��N�5����&rM,�?���:��
�Ɖ�ywh� Dr�i�ky���8t)g�
�Q�>*��n�(��6����&��d�6���Q�iЏ���p�ij"�b��$��(�X�KL;R@���CC;j쌻��q�QPs~��$����;b���z�\Y�ۀ��(Jd�s�+���W*�2�v�"�g��ڇp�m�����	�4�!������MLiD���1������Ŏ�"`zj͎�q���.h��!���&��!��J;�X? t�����N��]W`+��U�V,��z�,|��3ΝEnqú%_1L|fd-H^HC�]D6�4)Т�fP�z=�SX���� y˯Dn|�S�w����b�����![�������(�*���ã<&K�Q��{;����D�u�����"H�[���>䨿�IF�/Ho�wQ�O������2�DWq�����i�B�Ӫ����.��lŸ��[5Ks��Q@*���h���dߪ���,�����o�ـ�tJ}&����+RrG�U�#񒬧��zo��Ҷ�Ԅ�,��^P�վ�ܱw4`'�-/������D�	�$�����sʀ�&oW��n�n�E�p���`U�1��"�U�sI��6�A��|�z�c`&����aJR��v]b4�ua+2�of�F�G���m[e��tr��(�̸(���+��N��z��*#�i*hӭ��3Z�;Y�&�K
4�2i�b�5l%���<^�����;������]\����t2���H^�p&X$�ԈO�a�.'��Μq�k?;�(�^{Z�����aɑ��V� ���v��&u#P<��I�*����?��O�0¾�)��F�a]c�^�v	�g��_ަG[�L�x�AF�����Uߏ/2�� �%h�(�7���ŁW��
`ۂ~������v�g�,�J�l���jJ�F��6�b
�"��jԽk���g��`zY�/V�f������dY�U9��������i��4d@�k#~�S�A�z6n�ږf�W���M����˗����^����=HŜF��l��g�&U%ﳠ�]��	�SMw.���Ni�S���cB!�lnoM�y,P�9�̵8������B,[%w���|բ�+�I(�,nf�v���MoR��<�K��M9Ğ:�8/a*��M�)&��u�����P�ȳ:Eq��J�������g��L�/g9���%<�W�ɾ����1�*���Mx��H��yWIu�-˜��ĉ��$��N@����J���C�1R�/_�MS�zrX�\A?^J��r�j��]��s�\�cI���4���G�M��-R���x�W�2�����<�U����/*�|=O<���G�A�?��kخT��o*cM�ׇ��{�^�,}�Pe�9�z���/�_o���| x��2u��!cw�H�q�<�'Sn����BB����Y�V\!�{׃N�,�C85��@����rJo�6'����
g�C�l�f3<&8N�淖[��Izl�֏���O��}����Ե%����6�0���Y_Y��r�O�Kf�8PT���?�V��ʔ�{�J�^��jwj�$6M�O10���T��`�Ԍ���6�{�IHְj�-jR�_��	)g�qK�\���� �ޟ��~����y ���LU��֒Cg�?y�W�4�5AIT�����F�x��S��!k�;�'�B�T�~�:J�����ć��,�R�S�����yH������i�T)������"Rdίi����T�3�|���ߕ1c���К���@���KX�^%�}P��Ypn�K�TzU�|H��b�z8J�m����WճֆT��HN���@�oآ7
2u��N[��y�tCBR��4h4K�v��3E R��m�  ��1B�VGv@�C�z}Q��e�������Cs,��c�A�;m�0����L��(��o�v�~[=�NF�Dj�O����|e���
T�������e�����C�gn�m
E�s��#3�T}�;xe (��m^Q��<��E[�l/4*�:����w��{_?
Y�Ri���A���Oͪe�����M`�Y��\�b�>AR3�v�v� L�'�_[;�Fe�\�6����3���g��p�a�7�+�,��|�Ϛ
�r�[̓կ����Y�"8�lÏb�j��0RRaS���R�C�v6�%�$⷏Tb������LTx}�>r�@�UH�.�b.M�f��£�Lá�
��
�Md[b5��ndD?*�~#a��H�O�y^2u�P�Ȼ����Jė��$�˓�QD���繡BU�O�R�� �N!�&���'_�1RU�񻇞���i�5�ٔ?!�+�wg-o�+��E�+f���!�<�T�_uO��܋[;7�4@cH֖za.���#�ب��U�h��e�=�N�3��x���Ҵ8p��q�K��[���+�V�u�IyO�%~�Bݶ���=7�6�ܾWM�.����H��ӆ�J~o��4���G��e����e䵋�J �Vrĩ@��!+�>��B�iw��8�k�R��@���)�m%��"�-0�Y+���"�eL�"N���L���-�x���a�r�ǅ�D��5p�M�R`!o�4%P�T�Vݷ3�_@/�E,p�CC1��1��}�뚀Bٿ�T�;��P#��69c<�����E�l�����o��	ˠHm�↘��4��3if@b��v	�aϲ�!�����E�.�l�慃wW�ǉr��\��W����w�4�\P���i��.��y\�'���^ԯ{��`u2�t���Ӿƿ�����,���)W�0Ԣf�Q�<t�r�������|����k�N*���V*��K�<�[�еX����gdx	UD��]W{��J���.�P
|(���k�h��56Dh��`�vS.�z_�T/���c#ڃ���BmKK�aZ�e���	�a����E�t/Òn����
T�����(�y}��I��盳gΗi�[��tĕb�i����A[��;`��s�i�yt���Qݢv ��;J���O� !�]Z�I���<�j�ø��.E+3q�/�bVv@����9H#@[;u[ܽ��s�8�GV�W&S/��5��NY#�.��<4�5���ĝ�I���@5�D� �^���Qo��$"V�´�3N8�	�0�ye/�D����$ b�Ѥ�V>r(��m���SLQ�\�H�s�GN����#.�"̥Lg��Cη4(6�F�Rt3/zS��Sޅ�1kC2��p��}�7��#�8UY���z�l��A�����Px�6��8�@d�������B�^�X�NpИl�Wݭ��}�Uc?�'�Un�4/'���I��˿�,k?k�9nG��-n/�,{E������W�qg˗<u:n�W�|��u,�o
���|�W��V"�u)��������	��]O�����k��K	4���^m�'KP�R��L+�24{���c�q�C�ې~�_7K��V&� �����K�G�⹺���[Y��D`(D��_��{vz��!'8e[����������9CB@��� ��!���Y���&��V���O�x�F��*����hzs�[K?�����_�.���t�sA��������O3�}E;��PU7z�06�_xJ7��n��R�m���OF`@��<��@��x��PfFWo��B+���A阽d3w��悟�ƒ��t�7��F�)�+a�!�X��`�T��Ǻ�aݶ"G'�ⵖ~�wl�XtȲ�o�P�v�ɼ ��B`�
����La֨�V���K��@���X.�ȉ�g�"�˄�WTο�d �9C@\��n�~�Q���9D=F�q�	��x.�-:g���ARG�G�s��na��~ֆ�E�V2�����w��&qY�����W�.�k4('�FîX�V=��c�Xe�"#���.pZ��$�~���,E��F�����G���7�y�r�~�Ac�� �-�9�"�)%�,?0�ZR�'J�ԁh%�C��[�Vd�����-�=�X`�X���i=�����kP��]=\\��V�n�@�Lssm�4�/��յ��ä��
���(��W��c��_�oSC���@��kª$;:��	�����#��;}@�Hѥ_Eؿ .�?�b�m2���O~Tq�Y*tZ[�1R��"�Mv��a;�T����p9����� ���u0�c5�@��i���f +{�]���Rf��b�a��%m��y���:�s*�KUG]su�tGm�-���W����5`��r<J�0��S�%&�`��.qp���7���Q��Z7�js���kAQ�xBE���)�Ǵ������D��T�L���:�qs��e=�YO�������<(Q/d쒅�d�B����lm���C��L,no�������S\?	�L������+?�a���)�r�j$�I�O�P�I!%�vJ����d���;�e�H`�U��4~�G���0K���J�:N%�M�zq�y
���7�~��OoEc�%Q��@�$�u��!B:���V1Ίl�R�OgH7-Q_��1a� ����X�y��L��^!�,������؊��
t�[|�&��W�U0i��g&B��x&PzƆ�,.|���2Fg�Ǣa�c��6/-� e�Gޫ�l�Co�7D<$���J��9�]k�$���y�F($)�?��)6rU��#��d���K+��.�R���6���I��YMzN��{�e�Da�H�{ȕ��
g��Po��dpO2==u2��3>㳭�l8Eθw�������K�V�����gx��V����!���o��
��Hz��q�瀮� ����ʋ-�ic��G~����i#�1ք��;)w�bU�'�؇�lv�����j���lS!�}@��%9����4M$Jt1 ��Ա�(�{?�}����X^��yd3��Z��0ԑ$S�.!�����''<;�R���}~�!.�sƷ���\����4w�7G��,b*��0fǁ��$�}�;�B��A�?zj�5Ƈ��p�&1O��05b�W�R����{b�"�˦���)S��TF(}u�7B¨#(�e%�����T��Y)1OP��i�?��W4���Vy]�v/b�FPv���_��,g+uT����B7p^6��,�܅��0d%���!1J�є7�J�ɹ�Uj^�^�ۣ�]�A�=��%�n�-��^i����j��X<�4ǲ��*���Pv�&�.?v	Z'�"�V�����e�i&�#�R����I���
hB��ڼ�������6�*�/�������j���t�,Ph�7���B�����@nW_�����x�Ȉ9�-���m,>eh%X�
"�F�/��p�4#��WN+_�.g�̓��"V��Yl34��"Y�?(B�i�e}�W�߸��4��9Gɱ~��D������'�Z*N�VM��#��7�*���s:��DJrĺ�	�[��{����̲��ߐ�����(�k^=�����P-��0U�l��9�O �_s&�Z�a����t�� ����\�BL�,F@ ��Cź虝�*1��*�t��Y0���pլ1�<�ݎZ�uYIc��R>�-���<aC����:�։^@�Cy��S%\r���n�ڒ�N�uT�gQ�7��"�"TT��	t��PL��2V�Z��.�ܖ���,��µ�\�\,5B1W����5H��A)Q��������m��Ր���BC}�%��L���Mc�L�6�^LD�5�z��a��B�"�k�1���)�wt�jQ=�ˍ������j���5C�/���_&2�ӭ��>�H,y3�����'o��6��3VЋ/�Wg�{�(j���_�|l�NRr�[K��e��2����P/�Z
f���P�E^�fu��1��=��`���ޥ������T��Zt7�V�t�
*����!+Dg �\PfE\���tVV�e�����@B�@=!�o�WH�G|�����XJ��"��($0���ڎ���妽�J=�P@t=WM@���Y���ŤR�}�[W}bA��2�`����_�����q��G"��1AjDW�JR2y����ZB>�6W�Z���굚��u����V��u�%(<�aR�[�VY��|#	�M�ur��������n߁g�	��^����o̒9��R՘�M5�Tz��v���k���U��Ւ�7�-��c�D	S����*�Ƅ�&����k�����c_�f7k��g�v��1 �z&Uv?�rԴ��2 ��KeO�sq�ө�<�Ə�,��{�2{W���f���&�u�.�z�R��[j�
�0�E~��� � m�y<`�Z��W�S�����gE�ģ����g�K�����xF	���
(5Q�d��5=�tGA��#/)���qԚ�U�]�-9�,){f��F뇵�H����<��n���ɺ����U�ϛ؝.\Z���Gt�gǣ�O-�����:���c����[댝w�;!Ѫ��Ǚ���/49��������}�`��!w��\
|~�g=Œ���B���K�8�����u����	���$�k���Ƙ���5� �e�5b��W����4���Gy�C������ML �<�?��vw����Y��� ェ<��������!�5�ڂ�M�F��05�]ϝƨ6�TO���ϐ�a<Ӛ��@�v������
F�p� �E���=v���C�$(Ĥ	�J������R�� �F��o�������D�|dG"��a����iH^=i�51���q�ۓV�ͨ�8c~Pi>	邍�k��yW�ns��?lޫh�y�L��^�Kf��k��qk����:-�0b{���k�N�ʒ
��f�e���>ĞOa�yxbo��q����^�"p�٣	8�KVo|��M�����<(�$ƴ����\�����4`q��oj|��cc �ѸQ%��9��X�ٕ񈍗}� ���o]��(f�f��ws�:.����BE��s�(�=K�iX��X���R'�-��eq��؜<_�nQ1;�����Q��N_���0��_�dg;"�P�&��z�V��dS�1!G�e�Ѱp/�×�s��xo=.�CD$���Iv�M�n����T�qg���6/	>�fGx�RI+/I�(R+�{M(��{6��]�jNq��g Y�b�����6�O��	#��T�w2r֕=F?Ab�ű�MA^kM 7Z�^�`���!�%��"�����.��Ŋ}�6���.	��&��	8�S��x<�_l�Q���bU0���.6> ]܀�l+Ϸ�Zy6[U�Q<�"�e�����1Sj���_~���`��{��D,�
�t��<`�5���\b:����v5	��:�dn�7E�7��,�Υl����Y�6��/-�9�Jz�4�#r����p�NT0jUE0�,�sV�G��*
bnBGU'��9e��JL�<���������R������F�K�W��K3�YW�t��x��P%�C������-��3�؊���1�	����/����������o�'{��U��<�U��Us,�I]Wi�=��O���`&�ȫ�����am��f�)Z���U_�c8�t�Za���S��t�%�0 ���`䙥j��}G���P!&�����Bt`����{~'�\�š|�����CD>�B��P�|s$�-E�=��w�:����X�ɜ|h�Cٯ�S�\=�c&�R���zO`�'N<č����s��q1����B��C�T�!�yñj=֨��V�B1]X�fc����,mT�l����R�� �2Z�7��'엂!�$.�Mr�z�5"`$/m�˼�˘���*���Ң�� ;Y��wN�f��9m�7������\4jd�i N5�酠&f�Y��k?����,���z�`������FY@��F�<,�	�T�����@���-+��g���_ع�%���$l:�
c	k���g��E(�:���;9&��c1�e
:Z�,�׻�YȞ�*�-����̋��k�T�ҥuf�&~v޺�X&	ܨDW���^)p������s�h�#��(���Ʒt�ի�K��v�b�Z<pĽ07�Ej&u�ĕ���<�,Wj/�ŗ-:N��{����F�8 �S8y��֠n�!�ZSw�v���%���gX� �� �-׹�Mt?�*�[��
~�B����/����`�3O�xŰew��3F'���\��\5����!o�L4��ϰ�ڱ����aB':�����������F��E�0Y[a��~��:�J���J�����j�/�.�{K�Ϋn�wG��hӾMTK�
����YւZO�z�g�V=���p�s-w�0�xA�]~��-#ٰ���̠�җ�!J����2V[��ͧ�P	S9B/#�,�!9���v��[>` Y6U�g��?`kv|b\�N�����eQ ��0�)� U�m�b���L��5�:��Uv�*d��5Q��"��pG\q�a#�go�~�Ym�<6��#R���������zz#���}s$ݫ)��@YŎ�1����b.%Y�:�x����fFo'w/Q�]�v	�/�d���1ݝv4�h���|�� �� ���-�>����������G����Vc����
;ѧ!����p�?4ٍ�Xб�E0��z%uO_ǁ��x�զX TI��v���#}�Y�/�X1qΩ�F���㶼`��($C�'p�̱� wׂ���dUZD��I�k�.4=e�݀m遾�ރ1���X৛�ħvn� }E���1y�604sr6�g�OeG�;:wIR����[zԃmE��·�����o�Ȁ�o��,��P�6��,�:��<�.��V���c�=��I�R���h�DIɤ`��z��ef�?��KZ㫉�� ��3�k�?��aQ܏ި�;y+K�e:?Bv9��ϋ ��v�R8�ʇ]"{\0��}wNuۣ��1�8�)т�Z���!t"�S�#�r�m���|e��d#^򭌺�|�і#G&#����.���b��9:�i�-��ͼV�NV�\D�R@O�7�������k>W�ҡ�L��;VC��Wۜ��`��2����u�/��IF�ycgO0҈��K�ӅOL��-�L�E�N0 �Ubݘ�1��i���#]�/,�V+�	SԘn�br�W��Qw ���N;�@B�
���[���?���������#���[���O	�_�taX�b1�_��&�,�s�ot�I�R>:��O����=�I؛'w!`��:
__ۼ�e�^��	�1�q4�B��-`�����!����Ua'=HW�	��Mk�B?�m��N��߾u��(:���h~Y�#�9�Y IU���+�:�b�9���ި��ǲ�]��9��k-<�噤�K9�zrB']e!b����i�t�L�=��VH��0�-����V��^JUgY�Vg�����:�t-�*��\���Zh�rN�:7�Ђ�1�im�L�Y_g;�����;{�q�׈��qJ���UQюOKc[@��;ף[��m_s�}B��{���(8�/,T�1,(Wt� �{�:fp�<;�Đ3��((�iJ�)�C����t���,��
�*�J��K-�=���������4�h�G�1���YC͏�2i��"�X���?h�f����{��Y�*9�=����P���@i��D�ĩ��D�z�x�9�V6 ��6&��#��i��]����{����a��LMB�`X�?YC���q��!*�#t�� ԋI&⳯8��yq����nM6�`6����