��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jåا{�\�u�?߷�dn@6�zf��r������;�������Ϥs�����юN��S����xZ)z���T��[�o��-:;4�
@��eP���5Kf0�Eo��1Xn�l�@��ȼp[�lG�E�+|Vz��\��/�0�	���)Y��
(,_��2�e��r3I��慐��$sn�s�S�i���M�3 ��Tx�lQ �j~�1�%�A�5�1iGE�&3�~�ȬZx���{�˚�S�%��Fk�9��p��S���.�N��X�򡁊xn�m����VI�A�������?uRR匚�.�*t;
��=��b��d!i�w�&�}j(y�MOZ�dS_����E���22U܍H�R�^y���% P9�F
����0�����R��{X{E�+�CE�&h'��:{H�(�&��)���]v�d%�� 7��W��˥�����wRBM���k߯�g�T:U{hΤ_B�EO֑��Rs�R��2����t�G���ӻ��F�)ː��(I�ݞ�)�OE�&�\�'�&h��ӎ1��If��\&��Vo��H(�o^�&o<!��I��Mz�qz�N�e�r�Ek~�+
فaAf��硡��2u��C6��?fQ�HuCB%����ҧ��$�|ֿ��ʹ�Y<�`x�E�,����̺�پ5�V�Ł=����`^ �I<���JvK.^�D��57΄�`��h���9.3�黤غ��i�$�R�-��b�%yp�R��mY�jX�/�'OR�V��`�G&>�L��8���/�'>?c5s��(��ɖC����J��tn�������D�$j�	�s�9���e�Lyo�ƿ琝��1O?�n�?�#s�H:a.�Ue�}8��z%��Kzf����3���aDh�1n��!l�D�t%�zM�t����Y�1\#m���wAK�`Mjg8��@.s��L�7"Æ0X�����`pL��I/�=C��b�T@�&���ە��U\k��7���P��K�ԯ�e���=P����G��x�%hB>���|~���<F9���5��.�=�+	��]�|t�z	3^��p����<u��%8����s��~�޿İ�pO��(he�5�z�mC�u>�Kw&aXN�/T"�m��DV�����Ҏ�I�m|�|^x��3�ɵ�r�-Y0Xߓ�qxo!AX���V�t٬���S�0�4`Mơ��]R��\n� �P6M� �)���G'?�'"Eeg� 6I�����G�)�fT���)�ַ�jE^����R�kqX��O0��#�7΍���Nݝ����l~���wJ�Մ_ثÜ�	@� )�Sg�/�b���̉]l��b�_�ǽCثO�	8��S�o�_���j�9���s���oIޙ3PW�I4�E>��<�:� ?�gm����Q�|��%A}�Λ������k)�J����2a�:��6x��� Wm����sQ	јz�6�w
�;�#,�Q�a_�L�vsJB�������ڌI&�Ǩ�Bq�6��Ngl��|���WWVT�*
F���A�� ��9F�	�Q�u�E���W��^b��:oӠ�[m��x� �D3q<��
!Z.���� ��,�`��e��I��;�$��)�^���g��m�|T�g�����Ψ�0�ŔT��Ց!F:Y������可O�!0�D��Fz��S�ׂA�m�G�#������:�oc�NuS����>����|3����T�R����]Mդ�Ws�4r`m�_�苊�$��|&��n]�|��&�?���I������g�v���注�V` ��U_���(VN��� ���R���\X/�m3�����}r��
Őg4�nE�b��n]�<�jK��A��=S5Cױ�}����돌x�]{�Ƿl�)����F09&����Ҩ�=�o8W��sT���7�@�ni1���;M���� ��U�P;�kp��fT��, ��c���� ��m��|�A�s��t��ȫ.�-�_��.Z���9U�]d�CH_��y���$��������������)�s��`B�eTt�0���<��v���O/mw��j���-8���j-��dj�o:�ν: �,�ѿ�;D�st90� %��{c��i�ԉLت�����{;��xo���"���ˡj�aj߼��s���S5�j�[�m���O����X�ʶ�9ZPx�z�)P���G��Cc���S%�oM�O̸�ꙛ��X'�{&���{�s��'���Li���N<9; B�	�_TI"�~K�Ԋ�$�� �n�N��u�#zT�Ha�J�(F��h�2`�C�w]><�����#�U_!���]�|7��RS9�P��ܯ� �Au���|�,��l�]��U��׉\i�9dG� ���
�j��������B�(�Ne�A�<&�J��0��2���V��"���i�I_����G���"��m�w5^P�:� tCfEM;#���e����u�b$�L4�����,����݉�" ��^�[=�i���겈a�zl�'�"�>,6�fR��/M+I��G�&��R��D�*�$_*��_݅�^bS�m�z��B�1+��-���p��\�OT��g�,C--�Ǆ��L�ҚƶcO���6L�h<����g	�3�L)�����Ԁ�'k�M&fa���gj'D{eFT7]��7{��׌�2�L����>�\��xћl8թ�l=Z;ݤ�a�8����:��%i_��'�5�Q!���J&8O�Ϛ���V9`螼D�-{2��yqE-]z?u�Y�L��HR���H�4wX?��S���R<U������� o�`T�P"^JGS�>��?����ݙa.���|�*�W����U�ѼeǬ0������i���K��_j	6XU:������0��v�$��/Ѳ[)X��������c��0hV��o���c�#;��Rf �T���"���(�zH�	��p�kH���c<�~��[KR
=��蒻��v�u��:��[d�#)�OQM�޵������E��c�]��E #e�	�r��`��fFO��l��K�@���3�p+�D��A���w��I�+�p�A/@�n�``����u��<*�����g�j�'�<X���.��]�o�MU��|~��Zh�_�n$r�}�+`H���}&� τ;:j�:D�[�f�:�߀1<4��$�j��9W���Z2��?��"%W��<�=/��aQ�P���s��}~-�/RtF�%GA��(�� ,�	��T�c�(�_T��%��~T6cn�:�bn�.r^J��������Ģ�z��Fq�<}s��Fx
a��N�?�E���S5X�Wk��r3.��f���帯�,��y�W��v�a�Qq��7I� b�A������J|Q5�=���Kj솮J����x��8`I�i�c���_	�!CJI�#A�Z T��Y0ݒ�����G"	�*vSt�|��`�r�����f$��r��\&9X>V���{�E�"-�O)9	��b��};_"wb�p��mp$��z����7�
�-�nI��ss8�mZ�(7�&��^4��-�sM@�g����զF�=�mdj�Fġq"؍8oX��=��Wt�hb%P��__N��B�Y^a������g�!a:�5%&��C�s��i_K����g	�^4�Z��*-���u(�<
�F�n�Y�SA��BX�4ɴZ�O<0��-���4����f�ذ���y7�w�0�\�����=W�O�*OU�j���T#�F�Au�?�n/������0s�<������O,����߳1үq�xGY�b�6�$oĞ�}��,�RƋ��E$@���A���]9Fޗ�@{.��;{gh�hz�A� vBڋ���� 7�����P���Y��%�׺���}�����|��M�+7��[��7��G������	��������a�8V�Ť*
>�2[`���-0Ue�9���E,�v9Ov���~��ι¿T�2a:Ʌ�a �-xA�LN�A1�� ]'�*�|=�3��^���fz*ms�.w�q�?	�KE�k�%���#sV}F\G�\����_����X��vKu�,xG�͛�f��ô�A�+ ������8�I-����J�9π���j��f �>��y\�HXJ.c"�L���t�J��*q�J[I��6yw�(4RQZeg��N�B�T��-�D_����泟o�/8:�"~�,x������F���iwZ��鄌��;�>ŰQU���T��Z�r_,t�憞��z��:Y�V�)��v�dnqc�P��O�Gg��:5z�Q$�#�u�~-�I�H#N�؍sk�H����)���D��[��H�����@�[�y����'6{�O/���pFQm��Y%���#x�G��~���}}��B�d����'�CSk�,��>&J�Q/:��M���|�a��z�yM�=TA��9����r	@g���Պfr}�SY�ڬ��t��H[�ܜ2�\��G���2���V]=��[��y�"�]�\���{��;փl�;sA�����#&�U7��v�J�M��d9�d���ߏ��JL���b0�п5U��	���9j� 6~�-��PIg�|�ݵ���d��`P�O�ǽ!�Y �=����A�*�MdD����z����R�,�V��uNA��aZL�g�Do,$��~NS2�<KIYgM�X4pϚ�gA�ϋb�V�uŐ_c2�)���P�N,�~���i����w�� i��~%�2��B��^2+�ˍ@�:�eq��qy7B&9Б�gNc��&������Õe����'�Sl���ܒ5K������e+v�C���t�B0�u3�b<�q����i$����z�*YP�0�0��9�ג���31n�vF\
#���1-FO���갖5$��XF��N8�8�v>�F�<�`�V��K���olE"1&���sP�ʹd>�!l��ٻ\R��t�:3���=�cѐ���Ձ�Iϩ[%��ڢ@���N�4�o�O`�W�{�C�Yd0�׽URC�rsY��u|�9�`�{Ƹw&}� ��Jc)6(B
�w�v�`[�/����s��+��2��b�-�-�
�N�=�e��7��s�z�ۦu$�?^��-1h]Y������+���v�����_�­����ϕ�\�nKY�SI��#�P;��jivN*t� ���-�N�bx�q�f�XM{���O��׬�}X�g�MW�H]��H��7��'<V9����J��c�T|JyM����zW��Rl���	�yd�±��ƺyTB����:O��1�6!����g<2l +�ntN^t�[3@E:��ַE ��5є���v�Hre����,4��x_�E}�v�ۦ��+sz�
��Ɉc�h�z����+"��=�$ϭ����N`�zˤj��0�����D��C|��V`��w��1�����P�ȜA�V�W��V��χ�N4�����*�h�N ��~U�~>�A��VG�#�0f�0v�|�kF���E��P�Xֆ���rs�_�"]lY�ab̃wN$�ٽ�o>�3dk~y��lJ퇆���m� ��`���*�-�[k��L�_.���p����vM�3d^��G,�\�������r��<��H�h���c�]��P�����N0i��7 ����u�}�7��5�?�<q�:���$����a#Q2W����b���.��(���x��jd�#�),��o߬@���]ۗ��m�1�p�w��XءðYG�~Xb~i4��|��\��FnС@q@�[!�_��?�:�b�-Tͳ���t�;�2��_|4.w?�%�����@�� �=�?P�h6�6���x�>Dcp�s��T�[!s)��g���f�4�J�n���(���Q7�����Ee�[-��K�Ɛ����+����{�5ٗ�4v�զ��S�1X��͌�6sR�LB)���y��˜��?�WY��Q����*��2�h�ѝ����"H�ֱ���}`TQ���K�P+�6�;�0WAc<|I��`,Y�����C�C�3�~u���if�B�f�m�k"ҋrd|���\�4f�&�gU4�����H���ؠ� �k,��:to�m�F�'
[�+���D,���,�R��$�I-�7Y���*��*�A���<x�L�j�T��b�ˇV'wF�F|ԁNq��\�M��Dlt_�m�R9�c�Dd�`mc}�	�V����S�"�H��1݂�Nhwgy��҉�;d�`�U35��E�t W�͈��Ϥ�('����s,u�/j��C�=J���
U����^�{���E�vr�_��������Ӿ|6����M��{�V+6�8DƲ��j����o_����>�3p��Fj��*�,F�Y�'wŦ�u�5�e�կ 0
�/|Dpi����)	��(�� �����ȬF~Z�.4>�ڪ?��UK_�ίxش5w!�YӃ(t�~��j�z�m���+�1.����f�9��������4���7�.�EH���cA��u��$R���Zߝ+/��o̯/Ck"hOeorJ�&&���َ��)lY����`�bn���R�.d����䲞=���^0���7�L�ʋf�)"l��#C�%߁�:��'S��)oU���L@�b*��&kp����8�㨄8����h{�s���ɺ��HďK�h�سN��_��J;p�z>�>�mv�N�x}%�C����?e�� ��w��dĸ:��2�и�B�����̡��/LD)R@;|5꙾cT�K�W\��2���Uw*MM��y[W�+�}6�"� >��7Y6�6��{%%�L�d<��`ʒ����[&�F���@1`jL�I�?�NvKK���/)��ger��&��M�������bb�)�^39�e�g�!�ՌD�{,vv�q@�BaL�iB9����M�r٣���?|)�]�E3%�3,��]�8=��]��_	����u��At}
W�5k9��h4�S�˲q��m�s��"#6'%^����:�Y]����u@%�H��'~T���|��l9�4�|�	�����2����?�y����V�TpUdt��4���B��<3�p� �)��Zi^|�~q�&D V�ɝ��a�/C���v�8ɣJ�%��7gb65�b�(�1g��`Y^a���9�!2p4�AJ��+��=���t������q`���}������bed�h�n7�oFrJ����/����l^�����XMG!t�6���Tg�������.5!@'����E�b�'J:��t�F��2�럒bX���֨qT��2�SՊ�o��0;�����b�!�p���g� һ�����A�`(�g@V��u[V��<���aJ1�
�o�h�ٴ�?u�ll�e�ͼ�;�S��SMR'>z\u���C��h��1�n{�ޥe k=�CmV]�?�kmP%)I����ʎ`��jpi�y�2T���>WSC(^�f�П�VA����ӃgauJ�l��#�v����%A\�9L �������h���X���h�;��/P�<��"K�6v%Dm��DVاi�<T�V��JQ\{��:��l>�xC�>l���^r���>���M�(�*ea�Q�?ku!����->�ȫ�@�Tl����?�Ɔ23�PP.^��E[����]h9~�p#�F�yg=!��kĉ���42�Yˢ^���*��S�,&��@`[z '8���+�dLQ|�����ܳ� ��A�Dg�]��2����m��_"SM"��@��5X���n��!w��C[N�� �U�W� d�T�Q�n������jp	���j�Q�ls�O>��ڍ��rnM��eQ��ջ��`��Õ݋<�z�����4q�wM�����9��ОkН2���Ʈ`w[�PO��a�Pw�Nf3�
���ߡ)�l)�m�C7��$��o��`%yP�f�}ml���>��Qك�Ƀ�8���$d�yom��.u�H #�M�?]c�&�[>���hO�J�֛��>q>�{E�K��Ј��uӁm��;^�+a�`J���z�!����R���͠�� ��c��٧����"�:�*FB�\����b�^�up��s����uB.�]4c�!�*���`�t3�r}1����Y.�ݽR�۩'�)�);�R1�(�]{����E�:ؘ�ʊ%��;�R�h��}�o�I����n	�vv~O�p�VȌ�ҢACc�q���.�n߀����JV`z��F�ƍvt��59�<
-^}���ST$s6ۤ�u:�k�p��矠H���ً&s�	�4�{Gb����6������g�I2������'��-���XO�~��~[K�c��u7�߽�����K�
��=��Ȃ�&9�G�z-�W#Hh�upX����sR�J�E$`���I��Mv�A�h�����7'�:4��Xa�]�̤���Q3<�&r�6�9�j�(�]�_�xneUc������)�p��mڒi`�z�<3�`k�Q˝����C?�����E4��#���^��T�
���o�"�<�K=��]x��#����[A(O*h�����P�-W�v�����┱SHV��_�u*�4�	�Wc���df���l7mT��_�+����n5��V2�����ߗ�"^�!�wM��\�H曷mr~���/b*;��]��[gU6����'B<�2R�9��ap=N��T�X�
�ŭ����F�j�5f҄ZE��~��fp%0?D����@x.X�&��|&yT�U�F��S����C�r�����Y�f'+��sp�X!X��s�퐽#��u�m���kQ<;&1�-L��c6�w���2���+CqǨB[�|E)8[U��o�����rG�>b�����`���n���Z4]f=�]8�4D�K�y�7��k	���Qn���N��g���1���u\n����;<>�Y{^�l�r�f� 9V;I�*}���ʩYD����w/��g���2wC��4\�r���~X�OU�u�6����_�Yp�_�A��{^��/s�i;ӛ�M~�E�Τ����_��Q_��êU�Ү��������`��?�2��A�����ˎi���V��3�w+u4�����	UeܹZ5�n�͈���4 �Lߥ�QK�7�k���}D�+����(���W��M��A�0�F��M�!<A.��7I/L|��3�0��!Z>�I��g��+��xn�a��ʝ�����0)u���V�g?�4��MoK�%$O�띙&�J"Y�:�������mg]#3_J8��د�6q��LH�\���t�M1ϻ|�$�'�8�������E<0��.`j�T���~�O����5)[��.��F�K�e2Bm ׍o�$6sҝ|2z/E���� ��ƚ��<6�p�C+@���fA%�#���S 
}�5��G�"M]��L/��`pz�\2��hK�v�*�zǓǝn3fCb�����`N���ZmI~��]�k�e~��w��_u�r�~T�-i�2ײ�֟��cu3�-@�[-�8K�Z���T��1�|:�5 �.0�w�Y�=]y�M6�^�!W��r{�!�T�x��)?�,��0�q"ޢ����y,m>w�g"�n5ߢ�o�: fH�6
,�
��ݓ�=u3�Fc��;B�aɯ���H�fw��G�昋�%k�N|~[#�a�S�L�%�yl�
�AcgT6ۖ���{��!f�~R{�1j_�r��U�F���-��ra��Ob���~nE�\���߲��3���a�r �wu�8�U<?���U�}��U��$>$�ȸ��ѥ��1���njW
K,EF�R��~��$�w!�gn���>�}���~���]K4^0xfn︊�ƅ;b�i�I�^��%2�� ����xZ*]e`I�#8.?�����EΞN����U��.�ܭעs�3���9e���׽��a��^|���ZbG⠂_��$!��~����Y�|�u���e`-�2����W�P!���Ϗ`�}���Z��_�t=5x
���ղ.��,��O�i�ݾm��,�V/*'V� ���>l�[X�|�$�e)��P��_������솻Y�� /?ɻԎ��Yu���	���v~�T���48��v�*�������@��<6>A��nW��=,p��SM$��{͔����JW��c���2�,�7r��Ta����_b���X9��6Uhe�o�P�=V��x|��0��a�(�),n8�p��=�B0l($6�O�j5� ��n9.r���,T-wj=�Ex���z�̖,K�1w�����Da���j0��Ğ����	H6�a��@�j�ڥC�Gf�~�X�����85�q��U&�l�k��T' ea6��)\N���HN���j�T�гi'����=�R��OoK���9RA�̓��������e�X�������@�6�oK�6	 l5MD����C�}�vJ��]j4G���T���/�CGI���.B������O�	�����辟�/ �r�N&��~�;�W�t���}�z�*��>'UW+�g,��X|����2� �Jt)4Ԥ7��A�lKó�n�7	��X�%��!?g�!$\Г�٥YI�}�G��+7�$ϧB��DVXjB��aMJ��!�T�����)CIFy�z]m�GO�&��K����DC�i��`D��q��O���F %_t�������i�V'�{��wJ�'VP� �g8\��y~-n�o���PMV��wJ���{&����p�:�W�2��pϑ���g׬PW�f�ڋ-G�~T�]l�D����d�V���ZY�g`?��2���\�V�ڊ�7��L<�	!3F� �����46�����%ջU�8,K��8џS��o�~m8��⿩��U&���:�3˒��23$~O�4k�c����]��Mkف�Sa���-�1����uRǾh�8�|{L4�y�J��hA[���(�)T��cv'�����~�Gm(�|���+X�jgL���%(: �
��yyC`��/�QCxdCAD����J��-RIs����X^���ҝ)�Y��1�Dd�M���̝�?�!