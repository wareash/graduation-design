��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|��V�^�Z�4�n�	ޖK�|���DZߋ_f���*�H�d�s�^g�!&��u�$�T��+6���B���gRȵ��̂ͬ�՗�u�z��ZT�s>r�g�P^�VBo�\�z�����j@�MQP��2�Do�����.�✸����r
��F�O�a���`��oQJ%�����<vg$~L'v`��:	{ٗ��T̛�Qh���?yw�����`���A�����@֍ƴ��������/�lT��E�Ot����m�]�?~�+=��'�G%��'�+�S�	����q�yT*��
� �=�,:���4] �`|v�ѼЮ�S津N`��k���k .��T齥3)փ�3�����2�D������3S�y�㫉�w׎���O!�K(��"m����9�L�eͱ�g�zQr|;*�{��鿡�`��yL�3�ÞW`�
�]LJ*OGv�z�Sa���L�	k�G=H�ן�&��.�*O@�k9��I����4�b������(äȥ�4��{N��|,Qf��4�4��gI<=��V�HO����__��#mhL�I��9��`?7<'��&8j��x���C��S�!YWqg�VZw�Z�a���6�ܢ�����+c��ei�(徭1yQ"+�[���Þ�s�,+�
��:R�áX?aNy�N��Z���;ɗ�#���.���;����n�v&	��?�c�Ř"|�Ki��(S`�=��F#�q\��,�h:_������T�!%��u��l�"�9��Gb+b�Fm ^��`e�6��KPK�����8*�Q�}�Z[ek���aEB��"$+)�g������ ɍ����K�UŊ,l���Zy����HQI0ar�ǀ5��&�ԧ��I<ʔ���d��ˀ�� {nv�L珖���J9�1º
�KAΨ|��M����*��%i�+YZ�f8�[�5��1ٞ��JL�� {ti��rhF�o/��)�<��`nd{�+��/z
L�-�
?��lu�N�!u���ԫ���F+�n�Wg`���� X�7�IN&-Ǳ���xw����QLXx��gS�S�m�1?&uC����?�K���z���+���!]��C,�#�����p�[~k��D5�a����X���HRfE��=|�_���C����&D>�dL����w����T_g�0l�0� YxTUM?�A3�%��n�4<̛̐��R.]�!�Q`=Ut����)G�������H ���h�<n�D;��R�Z�g�d_�$�-�)�<#GI:���LDT�*cR�ò��Xn�b�(Zc_��/
�PBN��uщ��m���A�a��=������SC��0*�{��=3��������b7[�p�Pϰ:+-�/5M�D�,"��N����Cx}�yB�����)��;�xM���^�bE]�7���p0���Rlh_g�T-)]Hĸ��K�։(\���^��v����AC9��e$4�'�u���ES���d;�/?��� m�{՘�ف q�M�֕�������!�ȃf<��C]Ƈ&A���鿛G�4b�he|9N����\�qK��O���^FH^�p��q ^��@0m<�@�[�][�?uc��V�� ����j}���\���y�)�ez
�ܜWTD���ί����^��$+�D�0�v|3��2!j9z�<��o�`���dT���v�|�P��]����w8h�iT�P��ۻcs�G�WV��HH�4���]e޵;�٨�x��v�<�"y��xz,8�~�`�,�� ��܏ �*���%�';��cur#�ֹ�4�_wɖ�(��	����y�n�ױ�����*`8����&)��K�5���O9���]��jTeZt]/_��T�~�w��3O��(�`g����&��}?��n�zY��ԛ���<��7ioZ�+҄��g�_R4�9�w��Hŀ��v��w�ȃPҒ������fq�!�c**@	�H�C 67�cl9�v-Ζ�s�ߝL��Ϋ��El�o�&���*�C9�ˑ6۶7&�m�Ԥ6����mƊ��;0��8Yu��?�وh���f�Ӹ�?&|VU�KI���"�v5��ũ��/n{O�uXl\+D�;3n;�7C��Ϙ�����γ�@]��n�	�a�,,���7����w� ��G��Zߦ�)��v���<ʒ����;�I�rpF�w�P�@�����HbLìXƨ�h�yFx4�a�U��=W_�L��8a�}���c{r!S���DAS�n�N��Ѥ���$���[�ȓ���l���dy�J.�_����AA�-����w���'AԞJ5"jo�;n�7B�1�#f���I��{J�}�~��h�����$�Yd�1��;�4��z����9q[�����{c���|�%�����:NF��r��q���(�X�\��klz<nt�����1>.��aL��x��h�Y6�/�U���=�vk�9���i�x;��E;��K%.��a�d=ms@w2zI	�7� A�!��M�b��tH S�q�:�[��j�j�� k�]�1�	�wF��s(����懗	�^����Qs����;.vZ�	o���r;!yN��;�3��]U.�+	�u{���˩Y���5�w \�:�NI$\����:hW�S����t��W�%\(5�k+�q����$�f��=����a�퇎�\���V�S9�<�I!fhk�qn��!5�YƎ�2����uԘ�B{:��yp�¿�td�<�V����ӽ�ެ�r,p9u�T����!6\�I�~���G�6��=��n�#��$�7f:3�^�i�����@��������ء���}�^Hp��S�?Mp�*�Z��q;Ǒ7�3�£�T>y���(�E%:��5�ԖKtd���.�|��������������^s����О��@��+}��{�<�ɍ,h�qx���~G������+f�e6�8�d�񜡍��0���H��"��\D���s��3�����n+Stw����tQ���Fos-o��-՗��c�.�}48.�y��X�֬30�TB��N�#�BX+�?���HH���'��&v��E@T߆��1X
�$Bu[1�)�C��d�x��˱�Ũ�0���n~��|�:#g��|�ONn�K[_�o���f)���<�G�Y^^�6�u�-3�V�w)rא����,�}����/�}�
-�r)�9�!��j�V-g�X�I3��]��Z�N��c&���C*MK����|+gy�~��"ۄ�f�T�fa�9:a��?���X!���A�w�C���U�����k��ܗ�(�+K�B���+"�4��e�J|�7�j$uJi��+�>8�U�� ���.,e�*r7�ǜt��L��\�Q��O����r��D*��$L)�^0`�\w}�:q%�>�N����r����p�i�|�����:�Ut4C����T�9H�bU�m�)u����*Z��@�y���@����}��f�ta��=�:�oM|�O�].5n�w��?
W�x������.�cM	���S�s�8�{���N5��%��m�?e����rj�����R6��4��gP��v���n�K�:̊d�M.����#�RiS٦��fO�jY<\v�J�󧋙s�S�L$䙼#+�dCL�T��ǆ�ؒWC~^�\�Y�!�����N�!6��Wa�N��ݭ;|���`J�E]�N���u��
�µuX��;Y� Y�z����o�绿FQPO����}i���M%13;�5���`J�y��'ѧ s��w�P�x�Մl�W�j_���p�?*�ŗ ]K��ֆ�m-ŐDPu9��������&#MT�
,0-��^{�̗�(�y;��,?�����6�
ћ�'��3S=�R�g�Ab�iDNU}��Ö��
��4���d0ﬓ���b�����Q{[G�k�G�8��;!ҁ�n�� ����̓�ј*�� �cV'����Yޱn]�iK��~�4,77��>4��醭��=4s��`:%�J]mę�����*���B⃯��c�Һ?y������{��Lp�L�-_[eU�����`#���ԫr�ӭ8��eM=��O���qt|��T��ˈ6�Z*T7B^����IaC��М��,|M��m(��sg���S���R��kq^2��w�%,�4^Z ��gK�{���Հ�
k�Y0�K��
W��~�l�$��z>Q�@���L-J����K�(y>�Ԉ�V����� }�=V�Z���\2�UI���(\�i���2�*b8���=�
�֟�K�~��5��RY"����VMދ�
�M�J(^���U~�"��|�21�n���Ԫ���:�P�O�p�� �����`˾���uLC�y�X���%�5B��^5�-T*��)X��$�b� �i����W��E�O�I%�a��GL��̲�X�?&���(_���ߓts�̬'Q�=�o�nƖ�� �6Y���$!{�k���SIjV�'�[?+�;�)�U<�f@�ܘ������<�V�i�@a5�>�!�����/��(jMyI���j	�p�V1��9P֝	s�0�8c�r �G��K�䡹m���*�r�LX���%(�v[���2���G���J��F�i��"& ����k��-�wϏ��t���1]����Z�e��+D;R���]w
y�&��P�?�:��2�����b���!9_�)��\9q�w�tTX{Q����y��*����6�&���p�4��YB�����6�O}�G���ųhM$�Gr�'��&&�~�PzBrhV'����X�� ��L������H�fo״�Ȧ��Sjɤ�U����F9����A���Rn�L`�p�A�����'�5'H��$`�ݾP�vY��ߥ��g�Ϥ���x�ߦ�*�"��?OsVzL�Nc����<h�B���x�B�AZ���f?�3�'q0RMc��� �,�)�9�p���Y҆�
`z�������j�^ჶ֤�c���_`w���F�`
~��K�[�὆#k���v¸j8gb4��n�+�8���h||q;����2�lD��d�|�3tB���b�MCl%m<$���wŅ�J�B��:�6��h���ݳ�bE�
V�r-�`°��w⥼���Ի1ʍ{E/S(��bGc�?_���2�a޴��S����q)h���"���֎m�a�)��QB��a-�����n=��|�Z���b:�I�@�N���}>�x�8
��y�ZK�7�?�"X�N�A)l建�)��:�D±�z�����J`Ԁ�U`�K�ȳb�L�ck?��#򠋋Vh�?�f�W�E���zH)���5L��e��F"z�F�-F���"�#����O�kRܾ���=�	�@I��`��O�a��i=�`a�^�� ���>6��N���71������o�Q�Cc��H���[�v�/�!8J9�HY��ǵ,�KR��6���b��g8o��>U`mM�v �Jou���^�h�C���Vmm�+��̯&r9��c��B����5�S皦J�X���l�~�+�	��aQX2�,U��훾��U��v`2c"����f0bA�B�l��O�
�N�p�+%M�md^�������@�lG�ί������+q���'�e/H;g���H�Ou���^��g��s�K���yk5#�uB��/x-��A Ҫ�:x�DJ[J55Kc ����č&"L�B�Z���1�&��>(%���;�?��,p�\�g�oRpxl��9����7�}0�_#
����/J$�el�<H�w	�Y�)�����O��S��}�}i�D��]u�j���Pz)8\o�������*@RH0�p���2�����fqt�?�D�����;�+��V��H�������b��_�=m<��-��+��N��X9�sMnVK�4�ָ�"����B���
�����1��<A�4�@H\c�����ÅZ��c)��ej.ʓ4���w�"gJb������pvN,v�e)����d��&���#�|z�BY������;뀮��1��梧B���p�tI/$m7T�e��E���(�}�sJt^n��v}'4�,+:�_Qо���cz��s���sQ�}]O(����k��ڈ�n.հ��K� ����1b܈p��E�=�|�jE�x����gӯ��	�l*f�>��9�ʍH�:Vd�钬�n�1nßGiӵ):��H�NN5e��_��F�A�G��=Xƨ���0؜�%���|�n�����%��	J��u��I9����t� ����!�w���fr���&z�t��wR��i����^&&#�z���f�J�rA�����`w��g#!P�Cc�*��蟡�Q�t��@۸��l%�㻩�Z�#�QB���}j��߉��nVV�22|6�`t=�����t\�W��v�R��8�W�Z��GO�Z.ɪ�}��*�D7E@��=���>El��8��T�"M��-�+�x����)~W���P�A��-�_!�!,5��m�(��;:����I�l0���l�p�o�U�|4c�o� a�b�S���,�r��\j&���͕�t��hY؂��aLR�¥w����e���Xcw(:�i{̮fn����20�����:Y���[����^��k�.h΀̻r��A��ߍ��jN�]�⤇��ƎV���Y�Wv���Rr*t������`^ք��a@˷�/<q����#c��	<ހW�%�-9jZצ�QC<���t��9%��lGQ�f��q�F[i���m��@�3�g���՟�s��s�cnde�Ÿ��r&��ʤ-R�\lB�&Ϛ�x �Hz2F�#a�<Eg����n�|k�K�����`��H�h`�����7I�*��R8��SO78K��0�W��?c��I:G����*�-��`gq�n���࢓H��Nݍ�wkZ*z^��#�&f͛��*������K���q�6�)�S�:X�r�GAi^d8ǩI��w'1�y�ֽ�"�*G���i�����#EM�&�^5����0�$!6�q�ް��a��L��֞���t�]�]r m#��Pl��Z�q�V��q(JU�<�
����Q俙�=ٰ�H�x^g���-���X?V�h*�I�-�r��Ǟ?޶2w\X`iCT�Q�*^P�(�P�T~R�N�:������#]~e�85MŚhGJ����C>�w��P�����+)w�2�p�����7w�zK�R~�XMr�#����4GsqAk�10��mJ��G1���z(��J�KrWo�����+ u#�@��r�P�S�_�X�r%P	�5�9��h�:���	5$��Pr2~o�������O��)n� ʡ����3@�mn���e*pYXJ�1���ETW�Ewߎ��E���A$]��,3G@�q?�`7qGJ"�Qs�OΛ��hGL��A��Ӓ9Q��u�� �x	��g����Æ᪹���r���W)���Y��� FAg��Ôə?�V�:f"���y�xZ��ْ�P���1��bI�`�e9;�?\��ʈ�U=��Wz���=�A�{k���娹�vqӥ9sސ��po�
�j�^�U;��[�wJ��W��˫�1�
?pD�L�e?`!