��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jåا{�\�u�?߷�dn@6�zf��r������;��1��BIz�ĵ��P�W;��Q��7�sY�$W<���{���յ'�õ�R�#+�&TA��Hu�ʒ^5&(cm�غ�\�7�����b�.�u�:m�+���A�b�RXooҙ�<�0��3��?��3�Ao*~�ib����ǧ�48*:�0Z >/��y\���?����wZ�(^���Hq#��t
��|S� 1C��:��<2�$����V��&�qZ#��C;U�!��v-J7UiD�DW[n�a�� M�I�_�dJ�����GW}�i��Ӡ1w�L�F4���@0A]�7�35@�"�K��)Rb�m�U{���b��uY␿�PF/�F������8�y�nR�^�¶���G����Q`rT`�"&/������F��։8��C4ʡ��}i�g(\��j&��w�b����JE�}�H�R�(戮G��� >�`��V#yc��L�}}�/t�%���� �c�f��?�x�A'~�i� ��
��֛���Dp㮝�������M8}���V(~"L��8�W�R�$�Zwv+�����B!�ӻt�g�>�X'�rvI�sqX�&1o]�zKa�O�T�EܸndHh�,UpՓΦ���8x�8��T%U���SA���5�Al�fd�����A+)+����s��q���z�O�p�&#﷮]F趫�5��9����1ϱH2@=�Fp $�������,�[�dǚ��5�����$N}�����7�A_b�'��6�QD0P-�`nä4a��o��pp&_g���d��{��<�f� _�1������V18�}F�oj 5/�*ֆ�wL��f
�������P?2���x���gw3�,���ҿN�ה���*�P����,�Lא49���C�;��NZ�!�&��p$��wG���Zlڙ�efQ�>+���Us����MI\u���U2"��Qۆ\n+�+���2�簘Vކ=5���'��:"{D��e��iՇ�}¨��	��ԝ���d}Ԧ��@�&y���CT�.��۞t@��=�(�;�������<�t�U�ME/�%��Ω��ϰ1+�ϻa7��ѶUC�YJ6I4l�8&�;�g�t������L}���Ң(�l��N���X�I��_@�22-����W@-n����9��/-Y �b?׵���77�R�F1��<�[�b���߼��aE��I�F��������W�S���Ƞ�����S�\��9"K��ۜX��~�}g��[�X�4C�'Q(2�yr��~01`��ύ3!SCG�#H]l$���E���X)x���?ŵI{"�"0XUw���Y��Ŝ����ؼ/�紒�
�����kw�d�Q�$��3z�q%R}"]�Ǘ!q:ԝJ�)@HD"������@2���a�X���s����6��n6���mc�kê0w+��j~����x����aV�:/ �$�b8�.j������I���K,�L���j�ih������ɟM}^r' �����NH�T,)��eɌ��s��c�l��d�ng�IP7F��#�-U���O��K
)���W����̜�S����F�N�E�j�����Hd ��f�R�esu33v��o~�4�m�l��*~��	�v�E��T�_o(�9hV�%N'��>"0�w���X�� ܘ�®6��?Ǐy�l)����9����a��������C�o.�Ȁ�2ؗN��?�ֆsu.@�~l����i��aTh_&�@�r�@;�GܬM�;�m#c�A�EFf�2A���O�5��,��'�������^��S@�U�z�� :a������<f�6n�0LKߣ7��s������*a��-��(��3j�a��{�6j�l����Z�L߀R�C]���V�P+�S}[ꉤ�\�ο5�n��wdl��S�߯OO�����e|(�Wb^O��B?��:!<����c�
�Z ��H+�i�PW@�������@	�i�3�O�F��
�Y�U���򨬇��%����#^�Zd��	J����h�-���s�a�Xf��s���ޮ�΅�Z8���6k7���"l�pP�Ճ�"�Y;��њ����xs�!n 4��� }�9  n��.���ڍ��o�O_�wQ����7������?����e*��m�����^J��%���[����WKj; �`��� �=�_��a���.dڧ ��b�޶�YaD��6 �?�J�4H��,� [k�D���+��8�usn;�C����7Q�iCqk�IT�ח��<^�֭�������4)��]�t�Y&��a�my���
6�:ɝ��f�F�;��HD����E��1T*�^Aj����׹0F��|�~BG���Q�DH��a��IfTI�6��Z��f+s�ֹ��F��O?ѣ�����Ȗ^
!dK�FgBW1U^�6��?�g��1?r��B������QZ����<��y\);�������U�DG@O����=�Ip���������=���x0��|��<���ũ4#o�^B��C���J�(�U�3r��Q_����u����O�ڛ��h�W��u>�R�x3Z�G�U�D�0Z�T*��?���	���h�B�%�ʭM+\2ZFV�r"�Z+�jDN�T��!�]�� �%-�8���G1wHѴ����肴AW��Dd\h\�|Ϝ^O�+&�ǈv"ܲ揢B0o�m���;<�.(�F�x��44-X��25/g 7:�2nS����zc	�T,��d�%v#�����E��-Y��4� ���N�a��AVgMK�E���ٰ�=>���7SbC���ʵ�
	�5;I����+WCH��0�S�F��8�]���
>���
�x�l�!�q������+8I5$���k�t&k?��k1f�Åy�g����
�$��Z��f�d�J��Z�I��	�޴W2E��Ҿ�����|�*�Ȉ|k�T �\39��s�*���ˠfN�4w}}�M�J�����h5�P��F�D����q��f��9E�L���p"}4����ϞzJ6��=�vKM���M�n�C+f���ބ���vb�A�p����3�ڼS��rw>�no=πs��R�jpm#^����q���z�|�|�̓%��F�m�*�ϡ�MMF�.$ܮ ��j$�7��j]�O0(� ���O�(�'�9�U��۞���.(��(�J��u]r�)�Rn��;�������9�G��v��*{Ҿ����z1��Z�-np�P�;[T�2��q��T����7�u���/�]���5�ZtPd���B>۠?��Bg�=�L۵7���i0�iY�VĠB����5y2���ʶ �~pA��^+9y޸�6�jK:��qlX�!�"ۮ"Ŗ��'���+� �zPb�i9ޕb�Hab�9A�^��X�x{�=��ھП%&���D����?�5�6�C5�yځ;��?�7�M�*)s��K���&F58l��~�w�o�̢>�7p�lL-�;�(%���p�����
<�^�����!
�X����[�4g�1"�����f����s ��2Y�r}�� �R��R�
����	ѓ2�0�ݰE�?����@G�<���a�'	�J�������3t�ȼ� sI�]�6;"��+Z�t��г8?���6F �;��x��rX��?�L$��YBP�ޘ�]k�ꏵ�#�Q����x4�>���mI���
�j�eq��������=��Y��y�w,9�P��ͥ&/�; ��f�o罱��%����!,.'��>��I�>xy	�/���ι���B_��F�#�D41�u�{'K*�,�D��<��;�zFJCb����0=1�)��#F�7��
WD����eo=�E¥�񥴴�E}KBN�<ކ��up\s�����Q��B�Dӆ�ls8fւEZ���������pZ����ٲ��^��D�hW37HY����Y����m؜����>���gi\Ҡ�����1�����U�ےTR�Vž���hD�8��EE�R�P^lt��*�4�*��h9�������+��/ �R�}޻�����|����ew4�v� ���}���P��}Yթ�v���U��/#)	�F�(�/Ր�b�1�ˎ�wj�N���WC�ۘ�צ��ſ+b~���`��imm?>�22����a�	�s8�����V��hl��ݥ�F9�Qϗ*���lEBTw�4u��_�|�c0�ƺ�!�4Vj\��i�·�_�9񻇇�4�f�K��^���3>����Z��]��1V�*Mv�|UHRO�`f�+\x�~�<c��M,���O�ڰ��$�UP|�Y� ����AS��T+V�tM��t�b�Kž}�i)<u�#�����GG�h{���d����E��� p��J�{+$�3�D�EU�� �l��=x�e8qyVK�-���S�;	57���L�ay�jg8�ߦ�7T8d����!�Ol*�!�.�UOM$Zn~�/��: {Ɍ�	��z���Tk� ��xg~a6��R�3[�®���$��Q����h�ZZyֺ��-�_n�1+���F�;=������Q�N��5K⻆��:c����;�\:,|hbfx�y���f�/�ͬ�g�������%0��߼��B��
�H�����D
]#�t�<[,^trylҠw#��Í)'{Ț��"��W8Qֽ����'aWU��L'`p��#?	=Oo[C\qN�Y~MmE�Wt�"�^#�[�D�
������X�C��O)V+O���}Т?QKϙ��ʋt�l���=���.�D��b�ʌhO�]@�� �TXc
�	�p�t/�XL��Lv.�ď�H^��aQ�I2�"qAŕx�H�{�Ժ|�4�n�����"i?��}q�n���)W�Ξ[=�rU�^�.PM֘ၧ���'�a{�
�5�$���@[�2���Z�O�b�X,,�,� �!�#ei1kAgg�®]M�XN'�o����^��W Df�����f�aSb���l��P^��P���&��wcE���脙f"8A�ع[�&�KZP220��s�-��?��A���I�+��|!Rs������C�m�=c̹�d�F� 2F����*��,��~�;mԡ?S������
i�L��kk��_p�u��G��xǐ<���R8Ĝ�����;4� ��ص��/Q_ꔒ��� 'P ��V{�@sW����*�ȡ�qa��<פ�k��ﺫm��]�ddV�6�c����O2b��ԓ��a�z�Q		�
���7�����*@�j��,���R�ޔF�S7�*���,���Jj��F?ZT��8��}w9|/�I�HO�Q��r�s��u:�i@��h�	>VbwG��\�m/��M\B�uEO\�����z%1�uc�]��v��شy����뒳;�4Z_[;�/���m'���@�(Ha�v"<P���@ ��=�^}#l�aMx�	�� �B�i���^�Da�DOK��X���eVI����%�Zր�d
��N��'1Y���ܹϝU�����1�!��%|����b�m�[jAu=�
pA�vr�.$�R��Wu�V|�!�@���s�?	c�L.��`AS��{�l�KM��}�3��I�u�n͐�4�'Ѱ5�G&�d����LK�A��^������$�R�j��[b��h7� ������k{e��D�0@U��y��'�Na���$ϱD�G�E����L��V���m+�ÂV	,KI������@mo~d�t���������.��ALI�.'
��5������Kˋ`�,Ǎ���#�%����>��#}b�|�2,|5��,e�1�&)���N�9��LO_W��8�2����>��T�BF�Ni�~����0���`�G	����Aܙ<�g���YGX������?���}�KV'���@��+>��U�ɽ 5��E����(�48h��s�����xs��,8}A�t�gz�[�^1H��P��+��:�]jK���mv��p8���
��!_Æ`
߳�7C6�e ���^V�����ΧC�n��
?�58?�K����*�r.u�@b�>���G6V�X���%�j�Zu�Pt��D���_z(�_Iy�\�����S�Χ�q;C@�X��y9Af���^mŧ&8]���SM�G��5y��w}q��f��2�!�[��3�%j��*,��)�[�q��_�'S3�Ɏ+n�d�r���e����w�V҄�#� ɕ��?����U��[X��6�.#vV�e�V���=F<�P�!n�f�� ���R�H�{��7ү|&��}����[�=���B�$����j��xCx���%�ņ�f+ٕy� xL��NճJ��J��_,GJ�np,�|�2(����jmޓ��H#��^s�x�#���.��k>,Ҵ챷%q6���\,x2wԟI^<�7dՑ.�?�P�8>�D���`מ�P�:��k<��3�9�97p��HzCe��C��?�A����Uéq�IB�Q䠻mj�U����{�@���<�̑�Y �l_�#[ϲo�ZXe��C���X���}�#�*l�$�4���Z\�tcr���0�TCm9B0���Vr<��D��C=��7L���$�!�rw��֔�r��Y��S��"�۞sy���	5nTީD��7��m�\�n�I}��W�,M�	�/���aH�g@[�F��?	i��Y&�ŬA{��Η3%]��
c�l����֝�z|��ʎm��*��� |�=ۛ��Ea��]����글�+�Xu�y��d���3b}�ŬQA��^�$�=�2��BJn����a��/�
�J5ۼ]��Ib�U#�I���-G��N�Ѹ������!�6�o!i�DWZ�8O���u����&�$�V�LƸ�;�&OH���J����N����Oa$��,�b�>�8\���=9��V�q}�+��cB#�j�����/iО��f��m�@���pkp�f��Ƿ�h7e7��z����ѩg)�y����'Q, �+u�po#��l��w� �R�Y�`�d�=��s�߇�r��1C��l�e|K��Z��_C��SzU ��������&����`�N��bm�]���z�~�� C�K`� �r_)�%"��lq1c]�Lx�D���d���Ĩ`����G����3@�2nZ�����~=�$փ�P��yK ��UV�@/gaT�1�`޼R�O�oa�G��#I����z���H$5�D�>���R�a|��������_"d*�����YW��+R�Pz&�������^nh�㫪�gp�8��G��]ﻕ\��bzpC0�e�9=�9=�٤-D�G7�4��×췴�3�Ky>�D��wۆd�ʶ\��~Sq`������N˗4���if$G�F��n	�#)�)�U���]o
��H��|g�ʽ.q�)��X`�f��\^��~0��m�i�֙*r *��� ��h$��y��q;��IV�@�Q暔S�������!sgY��g(��w 2L��
r���E Rܷpy"�˰�"R ��6�z��������DqH햎Nrt?����5rG7������ ִi�
4�'/W�J<�^�,�El��ε|��%��Y�oߋq9���㟞6Z$�9���1����:�=�T-�^�Qk�MU����7���VAX�t��y�~l�i�����u3\	�'F& n�gP�^~�m[L�x赫B� �v�Z��y�&�w�K�����f$���_� !5",��L�Bu��}�H�PP���}�R�W�zI�:�R�H�#�%�e-Q;(��)|�CY�&� n�~��)#ȭ��;LC��w�zm�ω5J�-X��,����t�������� ]�굽ԇ��z���q?^LG$����E�:�6Pf��HbB��uRb����j��62�+*PH�U�� u*0��\FVJѶ'E��N�Vd ̃Cl�f���8�Z���~����T1����-�}/��([�iw?6�Z���u�}��t� +��z8��1�	d6�U��+DjX'���!�6F!�L3��(�_���Ό[9wk�{�x�K�!|�IU�RlF<LD��b�5@�^�I�2���m[�� �ҺĊ�T�'�h�7�B$��w�H�c�A_��u�!�� У&I�X���a����ݹ��`WQʒ�m��u���4s�zr��b�6㠵R�$��QX��9%�ʑ�x"�TN�r��	��xc�
Iu1h�/�q�ex	�<$�	�����Wm���vs��<^��L`���RrhK)���ƥ:�n��+k�Lրc}��nD�[�����0i��:`d��:��jFL!��b�@rs��$��Ī�~�?j/G��f4�@�0VJ�����
�}�Ka��-4��m5vw+r��rc������eb^o��9��CJ;`К,�4UH��!�Y#��\J]�srB�u�U:�0i''`�?��G=х�kH��[�`,C��n/M��&��
���Ej��gGA�kľ'�⨗��U�P� pB7|	�V�"lR���ҁ�sat�DUI��]aA ���,������az��䩵��Ķ��w^gZ=vX�R�+Ӓ����0s?ګ�煮ʀ�@<�bjY����_9Ѱ�йD���y�ʻEk"��H��7�L/#e�2�O'z�q�E�>s�a�:����+؛��!�0��H,��',ѯQo+DN���M�D���p��e7�c��-)Ƅ��Y�Uz��|����l��=M;�������@�|}@���}��v^M_�Q3�e���#F��C/܎A�p�sg,�J���5$����c�o�E�'��~�m�s��6*�<�zK�*!z@��^�j�χ r�l��p��69�N�6�)����8*�̽o7L��aa�aV�s�AZ�7�H{K���;�]nUA�B�2r&�~b`4����	6�ٜ|�Kd���,�0;�2����!
[��&��������L���X��H8S���z{,���28 �������o/���d	��	�C�M]�pF��ݞ?�_0~�Y�������C}���}�.n�	㐬�Xx��Đ�M��7Q���&��K���c���uӷmVb@E��W�QM6�FF���̓@�㎂����$3.C_��,+O/���&(�b�������_}O1�Nźx��K١}�Cy�Up�l���+,S��i��~�G$鸅�%��&\ȶ�n�u_gc+y�����L*-�� �6��SS�+��2R�x�C�vM��`m�[H��Ucu�Ԥ)�p���V؆#��2T5�QoA5Z;=��/�J�nU�_OA����Qf�-��������/X����ʛbk�`��T����pL$.��Y��v07�g����*��%4�J��0U�G�K��s��<u��W���5�f�:r} ����rڌ� ~�ĦĨ٠|P���洺0��Q�����v7wSM:��]E|X��oi�&���L�<4Z�;��q4�K��:�4K�|"��kv �ƽ����� ��!2�@64��Z4�|�BO�V5��h�m`��+����	�w�D��zm. R_s̕��n	�����B�z$�f^i��K^�pT�6!�zϰ�,���e&-���D4b��6�"@m|�h�7�� ]�����2
r#�J�=��7[u�P�~��aY��6�i6dm�<����9ߊ�۟;��_�oΠug�*�GOK���"�o���4� V���ݞ���AMᝣz�� kȃ�Y@H�O9&���]!f��M���A�&n�r ����xh��*i@���p��2�j�xU�ī��5Apx�h�T�L�F,P�ޟ��,�O��݌��oWDnE�e�b�G/L�����$j{x�_(H�y�j<F�8G�����Ol�ÝKM��{�[e�������0�'�X]9�.
H�-I�7�ڠ�^v��VI]}u�/�F3�"E�(�&��n�ʗ�V����ŴpYdEP��޼:�?�-,�4��H�q{r��6�(���Q�	�]\���������W�i�����rDwd��qWʐu��H�rd'��?'YhR+h�i���x����5*c�|X��Y��a4�3�H�TV�|�fD��F�/��s�y�T�6Щa5��^