��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e����d���f{��@����S��>���4{��ת�AO�Q{����YS􇡽5�����n��U�lc8����NP�/07}�\JY�Pg�s̡��sD��`�M�ͬ'�!U��[��ώâ�$�ƒu���8�c���/^3�2�����^b�p�9u>�*���\i�F��F'��x��3e��0���_�eI�Ĕ��Jla4,r)Q.�F�[�ά㔫��,��/!8҉��="%|���sk�h���� _r�u�&<�O=��_��R˞U�N*sx��b��6������4�XA��9������|�m(���Ջ��wl��gG(T���GQ�'�1��|��kM-&e3V���ԫ�����S]��k!� Gq�D�Z���o���j��=m�-A"p���!��}]py|���l����%��DV���5��r�NP�����cM��x?<-{��ȗvμB+����wW���j1��
��{q����d��5���[�.*.0ɤ�(����)�/(�K�m���EI��`�Y�l�r='����d+N�T�ļr�Y�#t���@����)F9��4"��8C.o�>ݦ	���^c+ij��%�i��_���%dȇ����9�y�"��%9pO�\+t�i���_���5Z"F��[f��Z"�&d �6`R��h#>��M!
s�	�`�M�M�PX��t�	�x�?W���qF�g
a^aP�JX�)� ᚴ��]�}&�X���
�����2��G���|��Y@<�g�����f����.���y��
d�W��~\l��ʹ�nDL���2�t[�H�.��Y
�o��9TJL���fń��ዌ�(�LQ�p�����ko]b�� �"á�/ܾ&���U*[���������8*>'�[�R����� �NtJ"�\�lT�.Eٲ�y��F�|d�ﵓVЫK%�$vu<y�s��M���)�`�Z-9��V��D%b�o��6AT�&���g*P�7�����FVK:_�[
�6�%����
�=���ډ~/.1�ɧ�1��6������������X'ŲT�HN��e��C�⃜_,(��Ң�\��x.Oe�ZM�ҞYxC�5d��� �!ɉP�|�Ȓ<X�b�����2(6�A,�$�
*��{�̲e�q$����>���z1��0R��p�����i<5F<*�*;x���(U��H,�|D)�>o��5�r#������ju0P��F�g@��.��ן�x��'N�O@ 4j�������Ɗi�.q@޵�	�,y���ߋ2V�I��C�JӖ�OF��+���8�G�U��4�s�������Ah��8,�z��v��F�Ӭ�6��Rmv��D����h���1��m�PΆxnb65_ SF<��d�ܗ���pțM�Y�	֪�ZJ�n�F��M9O��.���H��$B�[r��TRD�]�ޕz 8��Q*=�VS�a�F���	�x�R������m|���k�$of�L��1_%9��/��T藭۸}�����N[&�x�^�<�&SS���/��Ur��ΐ.T
�p��U`B7�F����*��fb�ؚ�f�Ǆ�<_�����!w��=���XD럴N�#g�����Ї�O��Q�_��$�Lo,�u �st��i%k���;�69�o�nF��@���ة!>����K@@v�f�mC2�-�ޮT��µ҅��n]�5=�e񁞝Eyy�%Z4��iu�߹�Vy��瘸���]J����j3��K�M���bLk��WJܖ8�˜�n����Q���a���v��nyy���hߩ/8�r�{E�	I������f�'\7c��`�~���q�g���2c�N��%Y�:G�-M���v	(�l᪳1�4����l�Vd&cB��\S�����t�_Z��ܯ��)l��6�#-S�x�)�&�I����P��0�r�W�3��&#� y������sa>����)��|�N�?pz>�&@l,�.
3y �C��"��4C�w�,.�Tr$^.��M��v����S( ��C��fL^>�i�q�M;�o\L.��!�����WO~�p�F��+!,N��[���
Q��R2j�Q,M�(!�8�h1�7ÿ�^,�Ӏ@�=\(�S�㭛��JzA�U��EJ�HI��Dg�'O�e������	2?����#��*�ἀ�LB�m�]�`r��%|�4߷�R&�q�;)Sn�F�8L#�Փy�_C-Z����^�
����}�H���./�*
����sU4�X�[|m@�3v3�9Zq"}_�m��'.�|>h��IL�75�+[<�yJ?q����_τ�( �kp����%�U�����7b�hL�[Ie�@�G⨂Զӷ�Ch9z b�s�lP�dN^ ��q21�y�vc2��@L::G�Km��#}.<z��Fa"LGS�À#�5uz����h�g��mE�yH��k9�7�h��%����;wMob	�ڵ+7�ؑ5��ꏄ�
�+���@���l�"��7}�2��JJ�f�%K�x!19�w�횦FD7O���q��&tMm��4@��K~
qE�Ҏ����s�7��e��
�;�K��#w� 9�e���:��Cw�(I�_�啣sM���lbB��ˌZ'A利�g�%{���O���q� <��� A���u�p�Qq��|Y�z���d��Ã9�����5gPZ����j4k�v��dKR��16��U�"v�u�$���k�Gz���5<R�M����x'N��]��z�ա�*��BE�22.Ȧ��!���������ߢ�ɰ�T�$w�F����E(��v1̒'Q�`�R�P��~ZœR�ܭ��|j��˱����t�x\�����N/���x���m!��I�W4IR����/3�Rs��0�]�FA��|I����<���ՂE?+|z�nm�e��&�;���ӂ�vZ>��я��*�2�\Ֆ�%�F�}*�!?��R��mƃ�H>zq!��`�*�4r���7��ؘ�Ww<]�*���利�z����91���^���Q8t�}Q�|LU^���W4�8-��,���T��6�>Rz� ��<̎[.ZT���t�2�r�����[J�V,P*^S�"�콲\���#�Dw܅kq����9}�Q����(�8�!]=�П��� 9�q:�Nh)�ٻ����3�w ���)�v
Hc��찶��Y#
��՝�VD���o	Zzq�S�|�S?�u*WV���3����jA� C6� ���gIA�WM��I�S�
t�m�D��A��
~B�>�C��t�#���*��)��zy�g��Gڥ�0,��Zg�;/o�џiK�*�4���T�欠����\3U�r�;w٧&L����`�]a:oB<��Am���KW�T��w���N�1�<��Z�Jq����p�)�����\�>ۋz�|�}j������D.�q�F�}CQ�T�����;��p�!G��d���ߟ(�hk[*�W�f�}Yk`�.���0V�|N��W:q��z�x��k��R��e?��Md�)�+��K;��F[Wj���s1��f��CZ�?�Fݭ�Ǟ�i�G;��5�.�SI�@QF���H�\G�|�7aDs+Po�r#î��C5�rL.�T�b��3sDK2���o �q�� ���^x�$�P¢��V��Ir�K��ύ��F\V��H�k�g���\��z�%�Zf|GbQ0���`�<�OGy�݄�r3�پ'S�G8�6E�$�����L��ӤI����(�t��OH���i��qb�#.{'��q��{<�]t�v�(� ��X	3�%t�L�~(4��}y����~����'���\�yL7od,���/�F�y�^���*�}��-s����������A��9?�5Y'���k��}�d�0�d��g@�����5/3�WB�>w ���Z���_O��Kn�`X��a����kuCiE��;Nӵ2�=�2�%x�r�;k���>r5��g'�WO"��S$��9�<!E H\F|?{�o%o*׷��ڞ���9��q�~*�;/�0�c4�4	.+r4�ق��&]>��	�����N땽����$1\g��D�?���rG���Wʥ{�{�B6ɶ@v!Ȁ@Cg��ė�S������/���9n�v��i���d�Z��<���RC �@i��#U�u˹��}�
�̎�F��Bx�Z7�ňOx\ۚ ��hA�����<�Aa&�2GJuc���D�'~V�Ɏ�ف�v����J1e��*ib���u2�40x�����^�*�ײ�������<�7?�O��`�?�KWI�V���bUU�[�d�-�� K?�"c���������l�{:���~*!Vގ�;���GMt����&�� Fx*nNW���Gè3=[I�Z;�x��$�3�cG�o�Sc��w[���)}2��-i$��ss5!Z�G����o�'�7��ڠ5�yxK/Q���Y�^��y�a�hhia#T	�\�.�Ώd�M'�pD�JHo�����8�a	���݊����q�[����m�F߅`��P�t��JY=��EG�>������/�3�����YME9���H��Ϧ�.;�ڤ���� �,zܒz�<�E��IU+�]�^�"Q=#u��Wc�鵸j��>M����`.Tw#�vڄi�x$2�L���E>q;�r�u��G�NF��z��'���VE��*Q��%Fyx�Q;z�V&�w�%s��4��ܰ������������:N�o��������I%�&�� N
D�-x��U��;��� ��h'$+�V��e�(3 cw�3f��ټr3��ʢ/�{{Ĺ1E��|t���笗�Z'#��b_��G��s��4<�ud��{{���m���V}#~|�"u�����1��t����>^�c �"���[.olK���1��<� ;�h�g2�����6��E��4��ƗUzE� ����B���9���Z���ڡU��X�:��O�Yk�㌶���4�'�碔gr'0G��L����hc�o�k[n�Y@M�}��;��@��v�?@�8��d�w��I�WZh�C�MF0�73r�K�6톇��}�<�v-��,Ż�A��)��D��9\'�X̣�Y��#/�	�}�BNM�.�����\y j����G�\���i�w��cN���^8�Z���Ab'�ɠQС'�:�?�ê��[�F�:�5]�}��g?%͖��Md��A��H�U��A�+���;×�]�6CS~�>�B�Xn�㛡��*� ���,\����"�)y�,�Y�Α���Σ��of�N�R�=��y��H���Q��v����|���
�d�9p���	��X^���VR�T��!�;���*A�R�
�m�a����4Ů�]A$ַF��2s��C��G���Y%O��� �b�Ĭ��b�\�?n�J8��˶��(0"1��C9f�h��v)`���ֻ>�c�y��E]��+;YlY�P�3����o/OvE�s�c��u.�y�<�i��(h�E�7�恕��^}z�����M�0�I�p�b梙y��"���oMa�K0�I'��;�l��4���g,@DN�$��?�\K�˦1�e��Ksvpz!i�A��Լ����.y�Yp:�Go��8n�,$;��֞�dL4���/� ��I~N�)zM�J�#8Ĺ���s����|��@��W�CvL��R.��'�Ko��	wW�e�:�$��2PO/��a%�`�Y[.V�5\e��ҽ�Yk�y �D%�X@�k��1��=����z�M?��0�������0�;
+X�{a������d�N��7�Q����џԱA.*U#�[''�k�o�6W�b���*�{��\����2`�,���4҂L��k��p.0�A�UJ�Q�@�K�k�V� ���n�	�qr�e-�좱������mqP���$�Vx��mٳ�n���WB��Ɋ̸TT[n�c|pA:!1��:���Ys�	;/�v(
Y��+f�2#���yМ����|N�;8���iY�=�H�$�非��!Kۡ��[Q���DK���N�4p	�R�^xB�h|�Q�v�k��V��ۉEK1�y=\^��5�UQ� M|���ěS��kͧm����OO�u̗�`���[0�9�Ԉ���	-HyS��.!˒fY��� �3���������`Z�dh ?�+g.���L��5����+�(ɓ���fl������OWАCFp��D�,�w$���mVJ	a���Թ���K�����N\����CÙ`�#��6~�	��Dj�[���-7�tܑ�#�礸��O�P��c@p�+=�{:�y�!Ԩ�IW�DJr�cD�G����,y �M�pd@��>2<n�|
�� kN�$ʼ��v�Dc����1V�g1'�@I �8�_��&���ˠM�8~������e�<&q'1�E�����`3���3�$A��0k�F��ere\
��a��=�WP�B��M A��_M_���#�2!o�9�՜V+.#]Iyu��[z�$8��<e7��P�D��c�˿�[���Y�=����2�?�ZOsO2@o����-�^g@Q�M�X�Ǖ�9ힹ�~�0L���A��[v�|�4c���*qhTEr�BN�w?�%��&9��J���)�4H�8�ѱ��j��L1�*�6���s�[��]��V'��	|Y���O��LZ�=�KEL����:s(��^�`��f��6jW�؂�C!�L��q�|���'Gk��R�����?(���s��SƂt��a�G���@��	Iۇ:=l�?��.$��_� CK�>���6m�~ֽs��&�J�z��ޫ���-1����mІ�D���t����w�,/���T�ۿk�f��m��*�#L>o�����Uo��Vm뛕�,Io2m���ѽ���'(�@�\�-� !�KG�Z�6��!�/+����9n����A���_ |4�{F��n���"�m,������C�l` ���

�0��'��T9V�Ds?pNC���/�G�j&����6��<�L:]L�)��F�����T�i����1��4
{}Ὢ �@���^��`=��mp�A�'�G��%�D�b��wa��P�졌�f��C{��Q��H~@'}���W���h��4L�k��N���J��a����������)'�������}>�L	���shV�8��T'�u����ȯ��~������X�K�<b��U�����-���S�m��i���G��h�9�෾a�h�
���K��`�1NOfC�*pbɌ�f���m�`��c��T`؃���_W{T������E�;v�,Y��| �x��`R&x:�B9+���U��Z���a�+����n�:�ǩ3_Z�
rv����M}��z�L��ն���;�:�c�C��� ���8�2��/���-܌�!�U�H�߭?�]�п	�B��l�������bg��`�o��2�;eP�/�����I���J�c�kV�W)t�2S:���}�]��K��ҿ���Y^���S�-Pq���,���Z�s"̫"���S�p�)pȍ�D˴��Q.&��#�4+_�U�6!Bc��i���G��_��;R0[��M̲�v�hZ%����U�G��/2&�NF�Y�cP�D2����2L�����}�������Fqtm��Jb㟭�&��W�U����<�,��{o%OmP\ߋ$�����:�ZQ�U#�[��*@�ٕ��@��u\RI~CF/t���Gs�/����xŭ͎�4~����U��Յ�L/ZL+���E�;pEn�?9+������ЁKŰ�JUu��Kz�*�Hk)
��Gm���R���ok����ϐ�e<���<��e�U��Bdt���"$��>^+O��)�ƈ<,!��o�9� `�W}�G
��{< s-ܝ���ln�
�����f��sQ��M�J?�}7���i�lZ�S�-@���ػ2ɩ7/ Y�=��n����@Mg��Yw����
�5%�l���#��9�3%�mu[2�)���W�uxzk�~m+��).�3�ԸF��Cx�E:d�P�1c���#�$Y�%�.s/��NG�����8���P���ă���ڗ�5+D�T��p\���_t�.3mث�\�K�)���e�d2������I:Г
^(6�K�+�+>^�M�e%Hu�+�7R�t�tu+��3oL����)��`G�>����2t}��[w���+ڴ���H.}H٣if�~���ѳoDC\��-s���3}4���	�m��V�0�e�t�x+w�g?T���g!�Կ;�5� �eT���B�	"�v�V7����s��"��t<Ra ��l�Ɯ��c��	�f"g�R+Y���
�9���I��$^s#����Z��N5��_qeX<�1J*���D^��;Te�GGE�܊;���4`[M{j�"=K|<YK@���V�-��-Λ!�%Cע�������+&�e�R���	���`��7�E)E;�������۟�a��6^����o��.�V���¥88d�@a�ǖ����?�I�?Ji�v���j��H��-�O�,��#v
�㲓�z��v�Vu@fz�"]A>���
]����i�]�]>��t[17��떈��:w�{&���2I:�2IWF7l�q�4ܲ�`b��Z�<��0���!�Rf���R������f� ��.���x�8�-I�=�=�X֖ƾUͬ�Us,8|C�H4Z2��8�ҙ=.^p'�Ƣ�*���]�zб_���Χ���g�xTf���Q�+u�J�u�ݛK���ǷAy�)U2�}A�ݥ`�+��D����K +ax%V0.�c�VW	7��2�0h�^�����F[�tO�t�Azdq�"�>#�MV��t�N9�E��9���)�?����0�@0P��ī��G�L�;H!�(Ρ3�3��U�<w:����/�����&�Λ���wt�S�XaQZ� Zh]��^u��Cb@R��.E^�+�beI�]gOv~8��%����Et��i��&�*d�BdH�Oҧ�?�~T=�}[��=�;��/M�B�H�� �U��ߝ�V� ����H���)�������Os�f';��ˮ%Ó��w����[7�t��h���z&�ċp�z��o*���.�.�D�.�]+2R����M�)(��c�4���q��FQ[����*�;�!x���^�$�Ԁ�]�K��=�u�ƹ�$�~�L�����:AT=!�E��/����T��P���e�օ3)Ә��e�����;�8�6f�ԩs�R��}��� �W�(�1�;�Cj���uYgc���Y���m8j�`Y��c�_�Ь
�[����ޅ0��:�s
Jѯ�Y�x�%R~d��x�m�|��������0w4r���s�q��̡6tFC��l�X��<��vR�x�_�A���+L������@d�;�P���'��A�:$H�H2�i�\�� �q'o8��?^#��0G����Z�<���hh$�ȴ7�Ohq�6G�t��~^�֙�ǃo`�

g����;E3W�>�}1�{�^Fgs)���1(��G���6�:��_���T{���W�
u6,�9غ�����G�'o}�$x���f�P�b���D��Z�iR}�ş=�]�D�͵����c�8៧H�����
�ߛ�q�E�9�=��a<��l�I�X�H����|5�h�x]7)����	g�y-w�@1�-
0V���җ�Ĉ��-���F�58��[M�2���*ēT
�3 �*������~i�V}"�d�3���1a{ڭl���^1&H�.�{�K�@,'���Eత���V<�+����vM�u���V'|���/���2 ��GZwsI0�ñ����,��(��I��5����4[���we�a	yw��=i���4S����[�3���}�z~�]](��{����ZUB6}6Ģ���Lc�?�l��P�:��.�`@�9���a�O ��ΊB���Y��W��6�WI˔V%ʡ[u�&5�AR������|IǨ��./ ��KZD����"PS�̈́�|<H��j��2����ߤ�ߐ;U�i����v'���ߤ���J�F�NC����ckh^��6"����:}����T���n!�n���[ٯ��rw��b]�N�����4m O�NE?�7ղ�0��"5(	�*te����iR���ł��sb���?�1�B�ޫ��L� �;En�0�t��8�Y�d0�:9P�F,��#g��߿����6��
ѩ�CČ�uU��<=N.OC����!��_�b�uQ�&��o;�����������D��L	��zA`�|O'�F�j�tWs�����)+�������x�bs���[�9LFjn,�!&e������.W��)u��x����=���(�]e@�C��u�v���u?�V:C����Ss|3�nv��[�$h.�SRbu��kߜ��܎[��T=����G�XS;gD(΅F�E���<������)�Үs|	J�0_�����U�?������F�ٻo��=?8���E���B��Qs���x���a3�hRu}��<;���+�[wM����q>��v*����ܾ1BU�|��d�p!و�m,����-z�j.C,�* &@��ÏA�nn<��r���z�k2�a��A���y,�E�%A��	'j�W������C/;�GW�������G��׆E6��d_��gp:�X� �a�N6<�'�oL�J�:i�Xi�d�z�[�(z�@.� qY�׳2�^+ʖ�q��2n|�?`���1�%<H�F?	�<�2:���6�B�	���=^d`�?[��.5g#��~궚�v��17��O!�];�e��-�6(��b	d���t�s��49�Zћ�W2������s.m��3O�F@?�)�FY<�-�!c�\�J��{�zP���mѺ#	_ؓ�WV�����t��j��	ޞb����`�\_Ǩh�`�(�bfG�]�cgY��U�#���^֋�k������pT��W�;�a��Z���k �f�l���Ѳ�bc� ��(�Y'���_?�=�0Cy�ʏ>�ѕ��}���b��-zYD!��&T_Я���+EO}1x����d�,�j���0�����o��N�>p�4�a�6�=Yۆ�ax�9P7��;;��#.GR�R���+�"��t@kQ��dgv�Ri���ҽd9�'�i4G7U�Q:�V�8������?������{X���\1&j��M��|/���*~�,s:=ApA!l,͓��`����@�N�Ţ8��$[m��_�xZْ8�<���>�#��*��
�7/RD��:�"�	p�j��ye��&)h��a3nez@�^��z~�����9��?ɫ�m�v۝̲GU�4?=t���÷�O�َ�S�����pmJ����1���kY>���\Ѷo���e�5�R��? ��Sv���M��D��5){�d�i����X��CF��1q�T7����*���򜉧"���X]q�t-�W�?���6\X#���9oAXbU|�Y\�aʾ�s��+�W�	�ܕ��4�ثə���� �\
�}����ж��M%��^Q�-B����u�y,L���\��	�m!�ܜ�����YU,(���k���gF��X�IR�JG������]ݡ��Օw��.�aI[d�"|u;����.�����3f�(6� ɚQODg�m,LY��g�2�����.|3=��U�J�T��nt%���͂�w�hW���byiUU?� ���6[B�רɑ��e�s�3��f� ��(���L�lֿ]���l���*�"M�}Q6m�n�,��jYKo�I!,z�EgH�����Do��F���b���gv⽅��"� `���;'ɮ^Ÿ+��A�Y�e|VJ��{�g�	�.��Ka�bdw�"]a�˿
�
�m�?0m �u?�{W�p���S;�o��ܾ1�f����$�Ь��V�^}�:���-?c�23����J�k�;���C�TG�vG�ڂ��/��u����%j�ѯ�>[U�M�3�FC�=���`@Ճn����eY��{t�̤�4�B/	�r�
��
O�s*�d����k�=��'W4��5���o�!f���j {�!�+�l�_�]�
���gӻ3���6��fq��[���`-Tݟ�q8���5"cCC�߂)���Uߎ�Q!� @�s�c��F����L')�H��N��(�W;i
SR��0(�C��2	I�~@��e
�G3�Ɉ?����0�J��Q���\�Xv&���$Ft
y��d��û�:������~��/rp̹\J~%o4ff�]��8j淿.K�M�`�D��̮ x�-�YQ���z����C�;�5<�e$y��d"�<��5+��	^(��A)aΠ<�K>@0ubh��
	Q1(�fɂC��.L+�;h��ާ��20a�Z-~+렡����TN�|�5��M�C��Tg����=(�+4
6U/��ަ�&�5��^�Փ���V[0;��%L�֯{�U%X+�����&>��M�bꕦ������[Ikό@t��lk��������p=�h~���ȏl����wK/q�c�)�'�y1$N��Ȕ�W��-����n�]i�
ή�ģ��8F ��]���@���:q�>h�W?��(�u�Ąl`�õǓ�mZ��dq���]e�Ģ�W+�ij�����bA���S��à^����[k�= �o��H���
�G��+���G��6�=a�5T#d�|�c2�_�IѲ���DZ��/$�Y(�Xv�i'Pk�ޕ��"�u6���z�c�3��PR� G�����d8�Y�6]�0���/�bU/@���eC�������61Z
���~J4Kal� Dz�t>�a��_��?ڠ�f�r1��*Y��-�j1���=*����;+���\̰"e�r���c�WaCL��=|wD<#�%+$� �bVօ��jufS����ޒ����ۭ0�F(�-8o2 ��s�z	�z�X�f�#3 �t��F�6��sg����S��B� $K4�M�9Ӥ�q�\����|�)���������oe���ؾ�>�W�5�l�����@#�1x6ڋرlR��gFe*Ƒ���[Z�f� ĝT�T���T;62(ޖ�,I_��Psq��q�SY��s�1�F�@�f��'bG�E�0��v͕�����y��M[L�p��AF��|��r���FW���RF��V_�3�X�-&�]Z���zD��$�_Pì�wa 6��Wۊ6[U�O1-Y KQ����z��.$�JT�"{��;b�@���#��B�gBd2��([�Hf2W����Ê�mVQ����y���k���Pe�a�הX�-��"A�r�x��F,E�,��r��e�[�lGV���(�|�h��v�l1�I�X*\�C�Z�c�3ϋ��[[�i�{O֣�mwcj���"���٠���"�rJ�n=�JF����W��GPsִ*�T6w0v�nE���x=��rp��6�ź��#�]I�a���d���-{� ��fK
[K'bׇ�����H�y�U�N�A�@���E�0�����(o��aã��ͯ�s��E��w9Ϛ���T�Ur�}�m/x�����4�dgޛ��������̇�C��O�W�c��M=���m�OWKr/)����f��#���:�x5��W���K�h��w�\�U_�\�,鵋�*-��V�t�)Grު7���cz����aD�^zQ���n������v<�@=D�Cd41ȏ.ʱ%������ �rW��"��H��X�PM.��l�8� بs͏�b�.V����
�_TC�yo�8�G�A��I�db%�]Q[�I�"���9)��;OaTIɀj�./�:�����K���\����qa�M?>��H��x�������zY�q��>Bft�Ѡ�EU��Yj@�.���?M;4�@�+;���R�zSĊp*��$ct��^�;��pە��[ɏv�%!,�*��趹&�֪�v�vؖ���n��m���ʼ������^M��>����*�^�ܜEm0z�e�4��J��Vw����N�t�Z ͸�<�1]��k�X���ʅ׽%=Q �Ӊ1F��Xڏ�Kz���Pg�H9���&֮K��������K����q*h�I�.�Em'�^��"Ϋh��D�QZA�b:cT?@H6~�F-�A�9�2�K<�+��,ț�~�C������ҵ{���j���u@�^���d���=�����pqQO#�tF�v��ڢt�C`��r�g\A��}#Yn5X���P]��3�SW^R,i�F��O(7V'OktڋJ�#��+ ,�>��W+�"t֝� '{�3��<�V�_�?��V�-��?�����FM��l��Z&��ŏ�.tU� ]'���K����D��A�������bN%E������bqx�����쾳m�����G��x%�%�;6��
��^��D��ɑu��@KS2o��������h��=������c�:J}.ql�=+_Z}m*I�Gc��r+��/zى����yh���xa�Q��YV��#9m���<�Ql2[<Q>���tq���g�q"�y���Z��{dAFE��BL����D��-�^�2?^٨n��=���E1tG?@�S��ȕNB�5F�)Oԧ�a���0��"��	�yQ��|9+��Z��@���i�m��[Ä�q�Z��<��-vg��F� Q�R����@��vS�ꮻNEh&���`�*�2�(������	�T4�ʦA�#`�~�I�c���,����L�aI��Ht�f�Tn�����_�a-Q��0.{�#E6l��	ld8��|Y���e�(�pADm�t�$���l���{�֋� ��'a��R��i��L�k��g���c��;/�!g�.6��aM=�j��_��M��{̌�Foz�ړ,�b??�!d��]ex7�p�ܾ^�P�@��~�����=D���� ��_��*����+݈�@�����/PV�7��)�|9wL����;��Ӥl!�.����e��T�B�@��ݽQ!d~9�aվ�A��C�"*uk�^�"�����D([L����^�q�W��Ӓq�ꢻ>j䉀���{�[�o ����i����\6,�rU�7&�_'�ha�<ȧ�t*,	�5)�z�����"��r���}aZ��<��rR�� S��h�}�l��QY��w� ���R��)D��4���-V)�b� ��ܾ:'&E��^���!j���89~i��#�_�n3'[ ��jt�Oi�K=2�:L�ў�ݗfm3��nq�1ɫ�;�]�YB���C����lk�A��Z�
�m4ڠP�̉�&��a~ɒ#�{8��nH�`�h3]���Y[\r<%�����EM�?c�Ho?�aM�o��_>�*��xa�a��:GדcS��b�7%f�J�j⾖���Z��kܐ��`j�E�-` �Z�CN�Sr�E�\��7���4��C���|�!fɇ�
�L �%5tG[d��Z*�J9��2��6�16��1�id�w�Ax7>y�1t�ȥ>^��.����綕��W՞�x_�S�J�R�2��_|Y�bQ��%��G��D��R ��p�DH�ɂ��kvc�ؙ�����W�4�_�XE?�����R��E9F�*�/�̙�i�TA�����f�{;�(?.�TԂ���s����A9Iּ�Y��>~����hxyW�(�D&d�և:��lE�{Ta��%?]r�Y�Ùv���(-",��@�!�=	����֯=떟���h'�t�����t�sm$��Uo�i<7,�0I��� 4"A ��ՠ~��<��b+�O�zD�X,�c����(+p9�?�Mg^���F��G4C�rM�z��GO��?��:W�4��oo�6 ��`�7?J����7���ðx�WI��E��z��>���m@�^���`���\w����A�����E���	*�mK��UʌX����z�l@�R�.�d{qI����ULyqd�m�f�w�V�怅��HDI�tP��^
~����w� �z�u��^9�s�q��tp����V&��/�p�i\�~ۍ䬂���OI��`m���["m޺� +i�X�+��"o�5���(���{_���3����&	,�!����eLH���*ʍr��y�z�Uo�w*���|�ek��w���6�re{���%z_����,��̀(�h�yv7Ӟ|v�r��bB@�U]Q6s��P��"� �' ^�_Y�v��R�^D�ꎃ��F))lc�
���ɾ?�Y�h�rO;�|���b�����a��֦�^�o��76퍬ޟt���#b[�3_���%������	�[�>d���-0���5���o���ٖqg���U���<�l���+:�T\L���1�%,�����D��4}n�z�[���l0\�	���"S���ъ���תBT$,�k�Y��.9�)��:�v6�L���Y�0�j�}yz�M_�� g�&`��/g��"���"oj���R�<�K��@��;�h#�V�&|�!�O]C���;A��CQ���$-��wD#u �M���jd3��|0���Y"\o_��r�Ch���߆������M�z
�(-�K��w�S)8>�$a�[ߐr���5T�_.��N��C�_�%��q���֌,�~�.�P8 �ă<����K}V�r��3{(��p;��^�o���_�F
�����FyS �/��\f�.��S�Y׎�n�2�F,��
�����&�๣)�Ȯ�������ƟGF�\+�<�B�TsҐ�5��̇ǿm��L�)��y��JzZ[�t�0���������wG�<�R]	e^�W�U���̀��R{���ڂ��(_���;�w.U��G�,_�DQ��9
�2�ov���|�P�H-��*�%�ym���fF`�k'6��ΧJi�t3̡�"WϥV�D�`����s����I�8a��jH��Ն�D�cmw��uv�1�ums�}<v���E-�{WFL���1�JޘQӸ�g@M�ϩ-g�E{rϢ�L`��wZ<b8�}�khBa���o"a��J�r��t�9����ٲ0�vIb~V��}�I�M�[f)hjZq������Tdn^/CtR�8y�I5���G�}JE�G���[��<|��z70�ÇA��gɁમ�=����b
n�;���	\��q/�k[���9O��r����Az�xظO�`�h֋�\n��1�qR��4����gA;2*��VDZ�|��g����|�����tj���� �̹eƊ��A	p]P����u�F⋔�喴����fܱ����0́~��Kh�#	��u4����	�L�^{УB��Փn�� /PC�:���a)r�Q5�3~i�&]4�T�ȴ�o\znf�b-e���l�r�X�o;,�U�9[�b������N���t@^�Z�/[�����Bd��N���v��9Rw�!��=��� p�_�o.�����~M,>��D��U�$d�u��N��m}2U��ԟ�K��>C���A�&g�# �H��U�`�_o
��P;~HIO�����n��:�ؚ;w�<�!�ʔ:�w�ՙ����U`��	|�!=�g�BK�$Ɨ��8=l��K���ك�|�|����?n�Y�Ou��ܽG���l�#)[����L��A;�AVU���N6b�,ҙ~�}����o�<O.N`>B���x����o����'cI�0o�[���u�M�wS�b�B@5_��!������k9�ԁ��\�@��ض�~���g��J����%ڧ[�X!]Fa @^j��Ye��Ǝ�=dȆ�"!C9��?�?<$�S�h��o=[��@)�Kh�"��@A��#���}���'�f�c����	���H��ZC��6��rM<���]�w?A��I����w��84������t�5J'�e	��{I)̯H,���5l~�-��gI�j}Zw;*�F�^��W���}�4�P�x��0{��'��o����T��剒���(b���,�=�k��`���l�{�-���<䭦5�ْ^6A�A��ӘA��7K%�4L��������~�F�\���
\ސ�*�r
�I�������y��{���S(�{f�	��]86	:�T��e��ES�	���ӵ�Esk}}ܨ��|�Չ�4|�Е�D�R�$��-�`�P�<����آ�v����o����&$UȌ�n>�)�ԅ�2PKۛ��l���(s�j��<�	�� 8��ug=m��ۑ��C�n�P�� �h�v&�Xy%)�8���D� �c��duP!r��$0��t��<Vu
����Z���b֍c��pI8��fQ<J�5�9=y*˹���󯚟Lu/G�Y��I*ÉF��]�#	�	����g07�}$G�5�!\�F�I�I,'B���wҢ�I��ۏb��=�c�!\��q��2U�c$qG�	0�%5�R-�+��'�i���ݠ�Y���g����������6E���2�Lnkp_*ck���t%|�X?-	�h�`+��~~ړ6�-�.��:%PDޤ�`e���E�z�a�D�|���[��-����	߬J����h-���f'�JTP�ǿ�Y��*�/���v<�q��i�[�����6׸<��C��Q�L ?҇5G� ��IRN$�&{��^�[�7��1�r&?��˩w�A��)
��e�4i����H����X <o�}���=;02�]v�Y>B_���J}��ȸ��~l�k_�����pˎ�@��$Rw�h+�Y[�`R)�;���>�sF��9�u�mǼ��7:L`Շ3-焒q��܌g`i���B�몽���5B�-�12��X$0>s�b��=���5D6�aS�n]��\�:kΡ�Z�>�P������c�fls�r~\�͉ǅ44�V�&�ۼL��.��I���soO��srdx���	l5v��.�:��.@H�݊�����L%�Em�"�}z�^����6����-�78j�&;�t���=�����,�qAV0<�{O������(\o(����	>]�<�pӕW5�Ƹ���N��!R!6=P�\Q��E$�oѯ�Rn�S.r��!+u��?�i�X�
tjF�� K�z��\�g�Jk��
K�O���j̘�/�����4^��h*`�ZC��h{�So���f��.AE	�K�����NvMwG���_I�I7���`-���������D���XWCI�y����'�ށ���y��<��0��݋��S��rB�0���s�e&��N򸜜��a��3B*���=�2Q����l^���·u�ې��!N�U��]�k�8��w�j�"{�L|���A4�k{��wt��0|�э����y�XxB��eO�$ް��.�~=�w�A�	>s�e����n�w��{A@&�r���dY
>�*Tn��*S�%Xu�<��ʀ����OE��&i�f�Z�LdsՉNu��&[qT��h��Y�@d����.�i=P˰�&7Ҍ�nf���|_.oVwB:�!I`�%t3O�������\O�A$8cI��uV�S�R����,Y���ߣ�UU�DB���F��pI�^&�|l�]�5�o�[��̃�{'	n�h��X]�Ć�Z��ps� �Տt�5�~�Ҿ`����
�V8�K��3;�9�U�U���p���~Jf�m׵�-�q����ʾ��Ѝ�X�}V��|�<�;�<!�ߠ΂E�g:�1��յ&Ͼa�NU�Z'�j\J¬Yz^�nND̟�˚ER9��*���G�欫0R`���#�X����أ``oް��M?����y��B�:1WE]5Mc�?+�!�Y���� C�%�[ð����̘x;4�2�؋>�-�7��"ȹ��G���0>-�o��s��D4"p��6�M�aΏm[ *b�P�w����p��X"����E�NA��gk~�6�1l2��V�������q_Dȓ(QO⟍�Ql��֞14��;�Z�i�M"p"��1f��8q3�Pi�/;)�8�d�eo|��\��]��^pw:�X������BwGdINPb{���[��KoV]�p�ظaû��p��u���?6���:G,��<����љ�KvRE�{OC	@1�χ C�!lJ�G�D��|���+�~^�Ga�_˷�;��!'�I&��/�dYwM�YF����|\�U�N��]�2�@ۦ��Ӹq�]�h^w��b���⍤a���[l�Ƥ�H�e��9"Ưp�]|��|c2�::J��7pvkB�	���3��8mh�CJ�s٢�P�Ǳ�y��������FDT�n��]@E������ꌋ��2�iM�d�YED�c�6�,h.�X`��sGl��_����$y���5�:6���XĶ~��i���*��v��
w]����Q�����)0�ƗuQ�}�
��u7]W�Ĵ&��U�����)x�"S���/�\�]�X�0A1�7��� v�ny���)�9�A`�H�Ml.����,��J[�0�.�1&��6d�|��
��� �K�}|��s�6p���c�Q>ɡ�зrOn+���-Y�8Pr!ܽM?���Lt��f�^;�>2�S�( J�\�N�����oRע%�_Q8��C���m#��'2-���h޼F�	#s�av��&5,<�RY��ܤg!P�W\F�zc��VG(�g���2�dU#��?44��nGy�9�~ِ�彏3��_�;f�8�
� �"@�wA��
����\D�i?�$ɀ�l��u�E{���X��W��;\�)��n���M2�1���!�2Nm��i˗�S�2�(��@��6<�WѢ�}�\�/�K��pU�g��b�c�~v����7m�U`�UlO����+�&"sFJ�H,?r�I��c�al��==��I�B��|��+J��6O�g�yX>L�6����m���m��˩�W���������u|J����j��|y�Ù�v��k��5��zx���h~>�輫�q
��I�DO��^�΅��e�s1��LU����;���ߗ�k
���x�.O=��v2'q9Z��N�̠�Ð�>.\�>4*�3��
ǳ�{fqE�~�:��Mߘ�%��膪EV�2U�������Q>�����L�*^�@�m�5������h�E����o������%�w������:�@	AX,D���ڨC�Q>�h@Fʚ3&��:� lj�@>����캗�� ��d��@���l�J�&U0!�	`��p�U
��Tu��Pi���׷U����� �������u�]g(�hۂ�@�C�#ͧ_��UR+�<��Q^U��LK�5��U*��n��a�	�쓟�6.$��p���Cܪo���)ݶ�@��3�i�M���	]8����� �rE'�"4�8'�g��Ν����(�T���` ��@���V��K�d��=�]�E.��&u�/G���ARVW�!�N�X����*�<��j}�y��M�4�W�&%�Be�k�t.J�PX�$y�d��� �'�������L��V���X���II��u)��8�����I՚��b޶��+��#��������a��O��PR���u����Pa��r�-�xd��^9�$D������y� O��^C����Z`wnD�_�m�O����u���n#���-���I��N�w�ϛS������	����L�����z���L�ɠ�&A�xV��<�wF0~\j�m谑8�~H`Eg�X��Sx�/��:H���L��e��L�$���`ȷ����ʲ[ϠD�x?
)hv7�>:9Iв���9�.�?�avq�6�.)�s��я=D�<[�$��c_� ������z$d�SQ�vngsҖ�q6U�~R��\��?;�E�����R�@6<�d����L�g_!A�x�:G�ߞ���͇��.�ڟi��)�&>�C90C�����+���H�
�:��&�m-kP�M�-1�QX_��we�Y�p\�q�'�a<��!����:?�Ì/�`�T�H̪����O������sUA�똾�dK6�m�d�~����te�#]��0��\G�!�n�#y�E�G�3��lޔ2����!���L̏K��t�ܠ�,=p���F0�1u�5�40�s2SMZ9���X��9���3C�[�Q���K��~�_����}I˪ ߽����^�;����oj������k(����
^�zM�t�*qx��@8��!�/O���&_z�b���q)��
3�PyNڿ��î�,���0�>mAӹiSE�d^(T���m��`Ϩ�+�;��)��o����+.% ��Ny��8������G*5�����b�,��-Olbj��s�=�М�#���D��_�Vϣd�ŏiq��k�^^EZ�lI��y�	�r�Ʌ���]���~gFPE�|8�9\�7�wG��ق@���e�����;�����,,)�ܪ��,�!��@��R��{��MgF�9�N��]����8>V���Wϣvq��w�?���03�m��*�b+$|3&I9</�NjG�2KF!�,��Af��`��Bp՘�<�X�_�mDdk�E�C;Zg��E�.!Lp�۪A�Ssh�c�"į�uMTN�����E|���≴	����L�3�1���8�� l��@�s�������W)+��MO|Z������?�@I��{�ߥ�ah^��s���Dp4�_qU�/f.�z�<��e�].��ĉ��#��j5A<�6���c�z@�����_h��r��7��qǑ�̻]mޖ�~ �v�(�صJa@h٫��ae��{T[���3*&�ȹ���:��@V��x�s+��vs.VF_EY��mn�{R#-+_�DU��vF,�Hȉ:���8���g��ȩ#��׊�=*o��K��
�64�2��]DS|��T�j]׈(���:<$��^Y� ���%�Bo?j���ߤ�^(߿�����P�{��p�Ó��o�<�SE��%�-�>��n�\�0�޸�����s�,��H%��;1�h���j���ܼlم]1
�-�<$�ߟ
��p�Sah�G�BZ�[ۀ����T:�bQ����0�(�ED+�%PN�7�i�KK��G�ٽ ���y4OPS���7�32��4~6��}j�H	�_���
�Zb����y�u�U��V�(��3��F�=U2-N���*A�[&&�f{tL�_w��#���`�g@���Pے�B*;En^N����R�;��ȏ���+ӄ۠7|�e!-�wW���<2�o���4��֐[H�y"`�6n8	�D�OL��^�ԣ��E�⽠l8у5��q#�؉4�9�s�:�a������ՋQ�f�\��g�����w�F��c���\2R�����Q�	ǲ�b��|��t1�I��C��^	��w��p�6ߓ��Avv
��1|aL���BKA�\�SN� 7?�8\�J
4�Qlgb���U3�UÄ��g��̧K��:扲�z���sx )|�
��(�]�K�Ct�uE�jT����L�8y馪��
_��6��Ҏ����}z�(��P��Y�G��_�t.�����
�91)KX��(YK��K�myJ���鲯�W��f#j�lM�ᦲ@��[G��}��UΨB��I��sr��dK����賢5���r8a��`������7��m�B4�1�s�~�R�0�y����gx㊪UǦD��E���j#{��+ NǄ�hƧ��_�v|Tfb0��#)I��wB�*X��b*xʞ$�-�%�̝������U��)�q�w�R@�)��!v���F`
.�L�O��ԮN�6�ф)����L�����R���J8'gW>���y�+�9���TF�w�,�.���y�e��O�h�b���}(A�\S�g{��c����i�y����W��ڳ>P��|O|�Z�`�!m$�\�ZJ�+V� &�ظ���d,��#!�:�	,�7��/���u5Ċ{��K�� ��h6������8~���bW1�ڗ��p;Z$�h]�$d�o:_l���uz?$�D;&��~1�\S��M(e��FR&W���찮(�Ç�;<~(�MHS'}��Ң'^�h�Urh������<o���̇�p�~7W�ET]�@=%�&��!�A>9��#���_×b�C��V�����;��#Gs�V��D6��u(�=�����!�S%��B{���Paf�%V����3g��E�U�p�>s�2��
�v@$����2(S����H��\�h���&w2���j��z(B�y�!�=S�����H���붴��M�ܾ���x�1Q#F���Ѥ��ywo& ��"jvײpj��v�j^�[�=Y8ۀ�?��UA:���<b墖�e���J�z�gx���EL�#�7�°4n3� �_4��:�N�Q�O����X��!��ϭ�y�d�<!�/�5�C^1o>CrE"UÚM��P��)E�� {����^�MM+���y���weu�V�<|m��FL�>g%B�q�==�$�"��#�ҕ�[�'��_4�.�*X��4t_�S��� |7ff� ͋�c�¤��d��2�SP�ܻx���5/Y� ��};'��	�u|6�����*˦�W�~i��q�R<���?G����z�h��YD�>����cf��F�-�}*X2�x�c1�J�ݾ;�E�t�M�R���S��ڎeo��Vt��ht�Ŏ �t3T�i�j�X2��o��K�����>$�������i��2o�Gw3(UC�9��K�,5�Q��J`��r�W�Pڲ�R�b�y<f���!_�f;Lj��$:�*�*�;~�9Თ���D����|���Q�H�ft�ݝ���O���2��d�GK�ϐ�����䉎���"���������g��򸢦���v�Y�snnBxf�z@�h�^�R^#d�n-0"�����WEe�b���u�Y�B!�ٸu�~,w���Sc0�#]�o �%�8����\��5��V8���v���j���'Kow�2��ڐ����d٭�מ�A����g��Q��$5���4��Gz�k2���	ކl�-�G7�̓Nۼ��\�o A 'w�@[t���v/0�8g&hg>�(��(J�e�Mk���sB�K��g �R� �p��7F� ��bo���F3���|�wlկo��'y�1Ո�_���P����E�T^����f��QI�	/�a�X���mx�������m�!�
E�J%a��{*���=��+���f����dG7�T�%ImS��[b蝟�sK#|��V}�p��;g��͏Gl�x�wƑg�.�I#���I�`�
.����Í�x�Լ����D�6ؗ���"dW�r� ����u����lYy�u�m�h�g��5�'F��X���A�n4[��e��'>��,D��EW�9O��K�� M]��B�b$wF�*�o���FN��� ND8��)�!+U]
��4C,����[�J�dd����i��V���d�;]h�Ī�4�L~qٶ'�R��-���1�rL����"�@���)�uѲ.4��8ܱc���v�����M|�ͩ���+�֞p�Lm�&A�v~�����K.-h۷���n�/��j���c�_��clч��~Qo�]&ΦiG�m��!���'�l9�i\^����ss��]|���V,܅�����u9\xH2yF�9��LHB��IΣ�@ו��+��:��t�T��(gR�,(A�M����>�U{4���Y�-�b�j��_N.Zg�!d��YHq�zF�Fƨ�*_����d��	�ͦ��0�;�3!-�}��	t�3�l�ˀA
�.7#�14������P�8�Ub���1�]�-��~������CA�~x�6qa��_q2���m[��8|1I[ �N�Ŭ` �r#%+Q�>��2�L*�(��z|	�Ҫ�c,���������rE@�|�4�O0�6gǧ����'n���Q,��qrd��.��<�����"�R�Zl�Z)�sj>e�4�6��Ⅳ���-@GiI�U�?eJ5�[���J*��#�-d{ζ��u1G���b�ˍj �K��A=UH6�t	��%��������e	�5[J�S�U�:���;�f�˖�L�M#�tYfct���d4L�SB �`b�UV��⨃��K�	�j�ڞ}	��p���q��ւ;;���!�L�H��=^L�Qm]���M�]5��T��n��C{��<wLY��QU�I�͹�&�]_b��^�`�AB��l���v s�)�'�^[�Ђ�}�<%�]��YL�p��ML� �Э3���~�H~��$(����7J��J�s'����نzp��AXZ.�Q�h�ՐT�
"�`�KX����|Nb"�&��$Jм��;�d��T�mk�s�X0|��9w �Ϸ����Gw��j/kM����u�^��3�z�K��ӗ�+B1����-$�0��qP�^ \O/���F*��8at�JP�Z]����Z-m���f�ymie�)oX�@�#=#d�+Ļ/��C.�s#����$�Q_�q�r���n�� ���������'�[��z^��4�X�9^y�	2 �a��K�ߗn>�*i|�`d�f{�r"�zD�u�[ ���5���e���oBr7X	F� y�?[zFq��g{V.���fB�TG��~ξ��m��	�y��8Cf�Z�Ϯ�ꅑY��t����x:���wI�t(����^I�}� c�l4�Z��T� !��r
�q}8�j� ��Ẃ���\H��@+H��	��3i���KQ��>U�U`)�A +�?#���J'*T B���ҕ�>�ʡ����X�򋝟�e�VΒ�&l��O��1�xx������yt�C�+`�����-/Ϭ�C�T+X$X`H� o�X����hY-�ő�Կ�j=�u�M.o�p�	H-��"���� �|2 [���{�6V�g��":�-���b�9��}��������O���������~?��#���Z���GtP�2�p��p��g>����sH�=�0=���s��G�x$f<[����)�O�n��UD�a�~!h�z���՚���sX�h�&@�|n�b/��,U� Bc|}9�</[~\�'�}�cr���Xˤ�Ԣ+j=w�B�lD|rM�e��/R������Z��c�-x��#���j>��H�_Lh��)	��1�\C�2.ط��*�L#q�6�+�:��)��_�o���X�	&	���<Z�K<�u����y��6���|}m�*Ͷ�{��i��������'n�?=�ɘ+�jwDWC{�cG�Kl-[_�W��m�i������,6KwrAm�B��#O�b]D��9���CVv��`�X�	'�U<ƿ�W3���Tj�����G[/F�r�)0p�φ*QM��{��;6d�Pox��1�D����^���Ă�t'8� Vܐ����\���U�h���߉ ��]݂����^�������(��`���t~��'���+� ~�û�O������)�)�c��ORf�Qm��Zv�|��$pd5L$��Rϲ1�L�zC�eyS'�o 1m�'�o�FTѰq4�>Rv��E��ޙ�(L����V]���	(���P���Lߙz���gϷ�ޝ������Z��L�rE��ZO!��D�\�������]tӁk�o}�Ô�qf%����Rl��z���MR�U/�3��D�C�X�[W)��Gdף�#.YBA{;�GB�5 LT^)N�MZ0�H���C�nL��)��;H��N�yȾH��?}�,v�q�DPz�>\I�����Q0��ֻ�ؼ�����f!B=���W���_��T�<,	�1Z�b~�Sr,&Ĝ�Zu�>)�m���:	ɺ�_�Q�ZfK��N|'L����_�]#i����
�G&<��s��;S�M��7��C��X�C�^"|�J�M�U�~�On��I=!&����fC[92Mv�ѻ1mګc�1C��	[Fm��L�����g����� b
�~¶����m���&��@��w�Qp ��g��7����Max&4u��6�O'��/8��*/L�Z�1�n�K�>-�B�x�'dY�s4��߂FJc��]s�գ�_4��#W+�N,��b�-vK�֣����� o_�^�J��d�YC��J�}��S��#@�s�:�o��L����b2�U�7�#��U6b��2$�Wu��cRdZ�k#��	�vJ��|��ޘ��~7�ϳ��}���?�B
���c�Y0�����`
+l���'� -�e��E�2l���~�kH�߂��;:рiJ��ܿ�B��{Ѭ��yNa��0��Ը�q����mm7��ք��0��֏�}��9T|�IX�0a��ap����UӶ�.�j2{�6�v�a:{Bk��D?��֦�]�Ye�*��

e�>7�}�G�eȚ�� �TT�:���FL���t�8Z$��4_,�(x�/	38��S=BF>1*z^�<~3|6U<Cu��OjGgk�]��I��g� �Y��T�Q:����m����?W�N����zrFg��Gm�3�!��J�߂��c�����\�݊cU�$@Z����u"���dL�9���A<�G�c�(��m��H:k��Wp�\0V2���}��t������H�e�z��̯,��O����v4��7HX��4Ɲ�n�^Ţ���X2��T�I��l��M��M�ĉ¨Dz,���BK�� =��R^�I��ݥ��mf�!�f����A�?S�L?�z87,��qw�2m��ܢ�W�m([�7�T��+DW�n���IA\	�P�yQ>\�lz'�o�S�2"-+w�A`��d����j��Y��>��2��z|k�0��!b\F�����$8�L�y��Z���6G���c&��A�N�	�� ���TԏO��e��h�g����_��/���s�ۃ!�=���׈"WXm��,t���& ����"V��l����l�Z)?)4�M����<~�vo8��H�� �Q#1:�Z��[FI�uu�Q��j�����8p�+[w� "�D&�O9e(']�6��̈́�@�7�S�K&+��\��^r�V���Gl8�a加h�Խ�j֋l��P��f3�\OJ;yc��/�<�Iu���3;����Rm�eՀ(�o��v&��c�z�3�t�O!���_RD�ƾE Ӧ|b�8�D���f���P�M��_̻?t��P��S���a|�tZ!�V�%��
��rQb4��b�}�~n5R��'b�V�/ƛ���W{��n��G��O�1h(,"��Ҕ���'�SNPq����Q���[l�v�|O��9+�%	������&��rye��ͤxho
����3� `�2�@���4̿�����o�'�\g
m�H3b֧��4�]&��5�`)��I�&��Yܽ�ˀ�7<<r����]��­S�h�xuZ>1�36�����x8
��Mw�sl�� �ֻ=Q���p~�>=YӈȐGL����.�ŻI�zu�-�i���-�%h�����y�i�H�k����@���T��:���L�m��*�ŜuW�e6��x7mYs��� �����,m0ڗ��U��;9$3��v"tXP2����$E/����S�"-�i�ҷC��*F؍���� �xlbF�ލ	��.�{]��K���=����G� #2���$�\!�=C0��f/�`�6�˄-���f�c�l�%uƳ�l���N3'N�����4�f���5�o�<g�s� Q�Uk�Z�	�WS�c$Ba:���Զ�a�0��ca~����z���[b��L�h6A	�,y]��x�?jc��D�������Ѹ��o 7��q9�F��@>܃�Q�	�we�a�tm�%L��f����ܕ�c�*�S�-�F������u���qP�Č�ĝq�2�z�������5��D�Er�ௗ��de���y���CT�9���7Ӑ��t��G�G�E��ؿ�^��w���r�@u�j�����;e�����#@n�%�E��?2��[��}���G����p]���Z� �'q�r����z���o|OA2��!O<���[�VhN�����g��d���F:�VE������ό���0鳙��֯����)�xi���z���V���#G�5���3�9s���[H�C^&LC+�kY�ga���f���F�rH�1C�FZ�G����o�une�hS-~Dv�
dsv+BZK%�h��η���!�
�g�:u��P�Iӫi�O5�G�r�(HĀ �[8\��ń���'�NA�bjh���|s��G�C�4�!s�dj�(nh �_�(� �Hc�[��x��X��e>�G���d�pU��e�O;{�$%f�9 �1�����B?���b[]��1"���0���v��T����������!7���L�h�G;�?C�	l݁[�C�F-�[���=],2�+�P#�a��87��V��BUT�(z���r�j`�$�٘EZ�%"��5�p��>��a��	�W�͎)
�8 F,Q��$"�H5'�9���+���T�D���2��@!+m��ɱ(c�˙�z�8���Lp{ĳ�V~SDr��i�-�B�x�ӣپ�Em�&�@�:�pc\N����o������'P�Dp�^Tե^H������Y��FY0��M/y;ڛ=�\C�ǃ�Z�{/���p����o�k5:��~s`r&Bq�
K{Qvi�~3 G!'�"�_� �����\'7#1u�D� ���R�#���GN�f/�b��bظe��;��	~���l7#��KE`�Fҥ\�*�.�-M���F�Țz�X�ݱ\�d��#/�ӧl�bf"�2�ܿQ�Q�8;r*�=J4�(!_�2N_P���H�cd?��Z۷6��{�� ��������̛��p\���&д�5���R�suW�"���įqA6zh��e����8zG���jDm�)�\YU&8g�F��V�O4 :	=kV�|�RT���=n��C&�E1���g��v6�(/J�w-������i�2(V�Gu��P	��H�k=�Ɖ>��^�J[�Gn�m�Y��rb�����(�4���+[��BaRFL0�d�*v�ǶW#}��e=qhH�-�m@!c����+\����Մ�-�	�(:m�s�'����0�B:�pg�����Ɋ�d� �8r%�)���0�m[�>���Hg�O�v�{k�%o7+��r��R�6����c�h0�Y� � |^8hQ{��p����@;���[f9�33�{����\A�
��Z�d����2��8�{��B�>GXP�`atY�V�pm�tZ����|��Q�z#��;�� ����OG%�=Di�P��P�A��B�*c=��k��`�V���m.�����ȱNÚ��R|%��s�-d��S�V���$O�ةXV���Z.��is�� ��b'6�~�DGE��ni{n7�o~�ţ���Au������y�K��Ik�������y.�)ࡁ2h�6g����$�	�v�!���$J4Kp�h�j��(X���@�S��Ü?vӇ��V{.`b.����I�NB�Nw��y�l�g���N1cr=����l��}l&��y���Rs����D��/E�H�1�Yc������o�qM��L
;F5G�#F���
	g�6��۔J@Πɋwvt�Nא@7�y�M9����sYO�ccdgЍ��.�v�=���&��V8p��F�_g8핉����]�/���p��O����w/�n��E��������)�,[sy~4x�&��VO[��Ba�;���Xin����]�<$L5 ^9��FGUFr?~�� R�Ȱ�˔��;n�()\��CJ����b�=f(��(0����)���0�%3e
�GZX�M>�WC�8K�"?��� �Ƈ���v<�'���C#a4�*R�Gu<����D=�33�[Q�KJc��zc5�2K���_�\�f_�����=���w��r3���'�?*�@�k���?K9�X	�7�$	��n>a���{�2?3��3�4I�^*�(5q��O�}�,G3G�<���fe�3v��-~H��Q����jE��~�"�`j| ��r��Қ������-
�Dgb1���\�&i.�'�t\#Y�*{Y9�����e�y}'G�b�}�y0Z��[P��u
�␡P%�0d�R�Dy���ޤ�~�72��n_�\bA����Ƿ�7u��m�Mu@�R��ݯ}�!
�m���8�]�z�˖������������׼�t��+&X��[E��o7g�d���Vt�x�W�Ѱ���
�\ƭ����	r�"�\7���b�>�um���F7��=�2��#��F05��&�������֩"Aq?��T�� ^��=�� z��F ��Qȍ|�En�o|	�0/��9�V&
0G�	��%�� �L���=v5՜K��g��.�!�̓ &�A�p��u'����^B�vA�\P����Q3�V0�~d`NX�e�sl��H(�nA<�7_�_�A��jl�{Ě����/������l�|,m0����Z�<�5�9�,�H_�$2��')�%)��ͨ�:��¼$eU�3����]c�H��u%P/�D�����n�9�jL��a-hj�@϶�F�i\�X�R+C	�.آɤ�c����gz�<��@�`�R{�桨��sPv��n�K�@d#are�fb;5*�C}��cP�G�
�l���+��i�C_���[�;�x�����t��ގ~���U���� z�c���Z����؊�u�ވ��~9�ƕ%SRS�3L�P[�'	'�	Yp[�1��S0; �mcV~W�ңa�Vr]<�l~׌����+�y	�_l����_8�m�E�FW�TH����m�v%����HdN�'Y�������VU>g��w諚d�N���Z*��ֵ���i�>��Ѳ�1�7ѿ��z���+��1p������`	u�L��ǫ1�\278��8Dָ~�N�!�������� w'�47������)e'�eJ8]~/�����Q]�/�hD���`�@��F�x�|�W�e�@����MBy"b�,����F7�#^G��4O���\��Bń�» ,ܱ��c���� :#4~7�V9� L0!�!�$�?��8���Q��b6�o��	�s�YH�|vK<}��;J��Had\h²T�2k�c4�,��~x� �,q}>��x1�*�G�b&Y���X$�+�@��Uο���H�F���)v���i�_�#ėr|7}��Ӷ��q�t�M���H@�<%���&(��c�Ue���AOؘwT z��,���YMp�4.�pXŜ#�Z��?IE�~�f4��V����4=�e9��E%vQ=�O�R*��#}�*�u
}���=.�B�����}�N}�Ǳw���]�$�\��Ƀ�}+Γ�su�d����ϡ��\"�<Յ�~��m�7����D����
����������p�o�l���L*�:,�.��T��=�Ig�N�$�ZMV��|��c0{����W�JhI���n���#JNB�n�,�\�cF`[Y_nwcNH\l�����LE�ڟ�4��Lps������y8F㻰�Fj���bnu�R޼|��HY܊G�T�)�bG��_��K0=WW��c`!��cj�ǽ@�s޾V)��Dy�萦m>�B ۡ�A��3�>8�������d)�A�ȝL����sQoI��=0��t���i�f(�?ju��h#���=�(�Meg��7�-(n;��ݣ��W^_�O�����H߆�S\�ϊ�ؔ�Û��&��太��Z���Z���.WNs^��b�R�Rjp8�{�I췿|������IG��8hjH~c��&�k����zs���N�����-z ��t�;�����r�P�ΐ{�����e/K��C�z�nmdŸ���Ǣ[��w��������hWB�n��).E)�cB�%��$��&}�����L��~�s~�W�ukVȱ����W�s��S��Vs婘�������[;�ʦ�d+���@i�Ӡ3��R����<��>�Rwu��{�w�em�g�Y������V8fV�G�|+���(I��V4���!��V��ˎ��g�UJ�w��1�%��D:�(|"J����H))������������#�N�pUX�z�:r���bI3S������	�Q��S���)�o���A�e��N��@������#54�l;OyI�0�?Бި��-��Du`%G20\�&;I����n�*w��-fm��.���|�c���u�XR�M��v��;_����vC��ĭ����e��H�M:e�q�����]���RF/CeV�o�&��6�O���'Lmק�|���Bvq��/rG�Ao!m�>Ki�kv���-�C�zb������V�:  N^+��N8��3�Jm����,VV�끸��{ß(ц*C��Ȟ�%ܕ��� 1�Z`��O�Wh� $&9M�i:��8���з=ɔ�-���X V�q%�}u�q|:ND�$�]Я�j?���L��������H�V~���k����'d:���D�t�I̘��͞8P�O�h��[�M���ZnHì#�`:�63w,�����������r��2C��� G���eRP��=v.���]�L���7��d2�Ⱥ������G�� �l=÷���[#) �5�HH�$�֦xP
�u����7�m����W�!��* ;���ݳuS)i��8Q+��Pp<���p1;��ҒR^c�n�	�6;
V�������)�<�d_�2*N����v�ȁ?0�T�H���G�+�|���\��E1n"~�Tc�����\��2�����)Գ84����{�a��G��0.{���z�����6�����g�f3���p`��
��f���b$L�^Pl|���<]@�o�_���\����ɮ��h��������/r������M��~�/��o�!�C�j)��a�T��;d#kx�fk�'�Y�����Q����[*����L��r}ZF���E�`�X~�#����>��F�w6�N�n�T��fz�ީ��!�ީ��M���Yl�n�t���O+�"VL/�Zk<�P���OSœ�c�q^Yt.B�x\��Q�g����n�^�Rz�5eF��tت����9`�`O'�N�۾Z��q� �ъ�P�O=:�am�Ĩ����\-�X��r����w6�a��3r�Т��]�ӑ+5z"-�'�Ż���&������Ah\կ�P��kG,Ɵ	r����kꂷ�ө�ez��@Ѡ	k�ρ֕��Pt�?�Q��~�r v�]uZ���;#��a<�M)��8i#@�t�v��'y,� V���h��l؛t�����i���������r�c���{FR%8j���-(�/nı��3�Kl�x1����p�%KF���kD.���E��Du�@���C;�`n��3�I�C��eS��cp	}f�\OO�b�Fi�t��ǚo)h�Ň#?�#�hՉ�,�\BZ��y_���s�͓� ѲyQ@�}Gd>}(��[�6��"��Y1�^���A��>�\.�5
������F7��Z�@���k�������@�;����(����AK����a��}f��Q�*�N��8C���N�7��	���XE"��}�"�
O��*��i�KطM�,B��J�Z�L�ܮ�T���~��R��g���K��kU`��J��?����������Bc)�����H~����w���D��3��j7��Q*`XSUkuE>���U�y�u�w���Y�Y��U�Z��쇔�=҅�����Q9�����M��S^x6��_���4�j��'p��J'�4,�ω�Ӈ�P��\L��t������6*s^wv�i����Bv�&I0V���,�Q]|�G8��;�="P��R�W�3���J�v�Ӳ�Wc.�r:MCM�w�T-�,Q��/�̨�l����II�5yqs��,^[<@�Z�� D?�sh�=���>7�������v��/0�/�{��Z/���`z����i
�����KP�[I�kv�8�E�>��?�Wȯ��A3�R��	E�dj�V[�Jz���l?�v��/��"G�I���(����_Gq3�q����L�;�O���꜑h�I��O����*��'��S�c�x	E��xޏ����X\&t���j-�4����	�Ҵ�c��OvݯP����>��ؼ�t�%�Z9��e���C���[��.�&y���9>YP���J�y_{s�����>��Q\5��.�g��!SA.K���Er�s���J�t�]K��q7�����g.�)xE�o*��[��� ���7Q�G/�RS3��+�R�J�W=���'v܋X��Z�^��D	TZ��ڭ�N����-��~޲}�v��5(~�lC��]���a|r��O��K��M����>����v���m?2,�(c8����n�-w��[��19�9�î�>�x�>��^@Naz�h�(���B�,,�E�����!-�F/Ku�H�G��[J�����1�V�3��?|,;%YeO�Z@�4��Pp�k�B�W-�6v��_��~��K��q꼚c��f�0nk�W���u;�7���xy{'"���i99�d:N�^5H}��Y�b�r�܍�GQ՗��7��O�fՁ�c�QN�*���c\N�r`�G�n��:aO&G�|j�A��8�]$5�ǳƬf��e���W��d-@�g�21Gި2��ubǨ�뗀�zҬ̟<P�
����>)�2y��ҳKZ4���&���{UԂvh��b'�g�HWK �����B��`]�ȸN��ȧ9e���twWp�O��[n��>��g|v9�3�?��C�Ӂ��[����q��q��~ay]p@zFEp_�+�g�E7�(���~�d	�g���D���\E:o����0�njm�xh�e��u����2�~�℧��b%�yF�����_�|�*B�\p�w�baB҄4~�~m�u������l���r�@w -�b����AW���ϛ��jd�ٺP�&.����qv��k}�9���y���u:Κu8oH16��Ũ�eY%�ߔ�ح�&]n��UלC��m.H�>�:�W�;�h�ľ�@���6-{� �\\&4��ʦ��m��z��!n��C�n<�A+0Mm?U���_�~Q�4�Q�_�;w�&�-��Gg�X��{���"iˈ��4�b��k/8_(W�p��D���Vt��R��O�ň�6#�N��1���b�R*D2��r���`ua�d����xr�}`?��4�_O^!$+���r��q���c���K���=���C3������� �;��D%�c��B:bom������H�5��$�~l3�^/�/L�1��뗪`Rc��y�#G��t�r�TĳMfFP�/���I���7be�X���3g���ȧ���ݵ�)[��َy���:
��ˏ� O�����Z�ӽDT��W�7��x|nL��e)�j�^��֐*�c
�j����T�Ȏp2d�X:,���Z�J���!�1\g"��_ճRz�k՟�a,ֆC��Đ��|��,�'��ۍ1�0	��'|.U�\O���i2e� ��H�`n<��'Ǧ�X~ZK�W�;GMC��4�ߺ"i5/��Ӯ����L�V��\+c��Uv0_1m�[�5k�_F��J ^� d��*����Q>C-��^�7���T�2h�~�b��7��\,��p������
 0cfFz?΄�@��W�w~rX�����^�y�4��K���9�)�;�P�;�{���q?������a��xa�����$g�lc�"S�qt���~z>!�M��zծ�lx��:�6-.�V8�_`��|�*QV��Y�����
�����Vl\��*)hH?:bpLe!9G��>�^��Z�@�{S�B7��j#�tG��/,E�<�
ç!�ʻOHX�Ҋ��)b��U:���o��33X�F�@s�K� �� l� �:%�������o�Si�r�S�����$��T>���K_3?�
6P��X�o@�ƒ3��'�ۙ�zH�M�M��M�V5V4/�B ؕ֏��(=t�.�?�IfVt�	P�n.TI�ճp�HS��L$T�8-m`[�\��I#��E´�G5�1/_x���"�6��� I�u�~��0�c¯@s�.Vx�Jp�	��9qzΞ0Y�8!���Eu)�[����xB�z *�_�@��8����Ugv�&J�& ���C�$����hea�_���yS�J��2��u/�s��j��`wV!:̼!�:κ`U9�s\����\���~�=���}���xE�xOJ '�*��UL�g�~��'o�;�|=�:�����.���	��.��4��:�ǵ1���P g;�'����H�!U~�S�3�0�d���0\ ��W;���~7l3��N�*Iyf^ǌ]3з���f�1��n:��,��yɽ���d�p�*����;����%�٩?������VD�����$͠��66��w���$�"E�
���������������z���r~=���!dH�_>�fBk�݋����Z
SѠ+#vUpI'���&������)��!�Y���;jM'�QZ*�ܨy�m���]��⒦����� AB4j2VBrCȑf
cKW^���9�Rqux�T�"�	7h��M�v��g��e�����=P~��-��3����ק
x������H�%ND?��#��"��0q^�c�w�݃D̀�rM^p�E�Xg�r.2�n��`L�u�U8 
�=��3W��D�:9�Q�N��_>�8R��Y������]��Ǒ���y��>�.)��N�Ί !�^_y{)���\�}��au�a�X�V�g��5���Ъ� q�<�iAs�- H��'Q3��N��.��S��ӆ9��v,�oxZe�-�d���-������ؚ<���}]#n��V�'�p*�Ȫ�<3q��W�/=�2��LNy
�%�z~�'ޏ��aݙG#�E�9h#&�g��{'�vRB��DJl9��A!�(��)[��CG�8��Nsqh��܂2�����:<:F�'՗����٦ϐ1�A�n�՗oԮ�]?�S�������N���(^�`L�]�,~�\�Z�bd�S��tS��+A�;�a|��V?�`��-&V�4�?\1�S
���~�P�*�y��WD��K��(�T��CxN���,?��׶�+��[���C����(�����".��a���6��T�3O� P6.�J�C���Æ]�F?_%��*��BW��/[������5G�L�̢�_�RI UA[�@��\4����׈�O�<��)��yR�K�i�sG���FB�������"jHvg��HP=�ʧ/=�򖙕AbЋj �Da�R�w$�4l��G���(&�	x�BaU�b#d���8^��D��3y@��x�VH)
���_���N�I��_��y7��Ib�͸½�b?���1"�R	s���}��c����!�mI7fU1���qh��A�{phE}�L�(��a��h�L�.�o˿��s���ɿK,ô�c���b{l�ߏL�����)��)0�8�.6d�ķWe�PS+}��ek�3��;=W���>��"e���@��%��� u�����Qpa��z<G��Fvx<e@0e��{��@Ԛ�PFQ�Î��G%���f�4䬼�I���{kV����Ʉ�|[����͋�7�pAv��X] �yL7B����B7x�(
8�|����4:�dMP�`�+��9 �ᘽ����Ȩ��o$03m	��oVp��$tl�Q}�aT!M�C�mP�c�}����������{r�{F��֜(�[TZ³ټA�qN�g>����M��uG �@k.���!�\�8�a�8�yi����8� �(W����&�W0g��G|�6 ������	��R�������dl� L�t�h_mx���3�|�$X�ՙEdܜc�[>�ea�-$x|;tY�r���v4��V���'�����1��U�G�[�����`;�"@���_��㑈r�0����?u�D��{�oQ#�טrx~���,���}gQ���#+"���.�\H�Y������ME5�(�䱵��W�!�BX"���D���"ʵ�S�ՉVd�=�*�BB�Pb��Ap��ݗ
��&���ܴk�k����E�b����4VA�j�^L������vT�bL[rp
~���Ь�2e�i)+-�����t��O��S-���O�ܫ�_`�OB ��<������j�Jk՘/�)q�)�^��a�]A��r���
b�G��:��V���%�E����CV*Q�0nw`�2]�6���P1��|>gNI��moT��"Lc��7'f�'�
q��p2@0��.ud\ )\Ś=���r*Ad�u3'��>�ߩ�$�'�vW*��+���<���迍�e�l6�Gt��FȟN�I��Z���꠳�ڋOI��l:Qԛy�ɓC��>�֏Sb��vGR:7��DY݈�j�[�"?]q��?e�^���/ʼ�7�""�D#����_[�aw�$P ױ9�*���j%V$�dW� ��Kb�_�z�rV��vK���3��ɜf_�"�^�p��S�x���r�͉Q@8�@roc�-A�h�;���&�{:G�����l�R�Β�u�"�
�!�К*n�$�����W�1y��99K�^Bg?\f4�ɳ�>ۤ�,Z�"'0"�͋�m`WmO�/��P$QR�6�'8��5R>���߮�l�/�c�h�_e��,��n�8��c=�B(g*J��= �);�>�g���~�ʄ��g@�R����+r*ɭn���6_CU��!�?פo�2�rBI����Gz�����xm���;�_D��y���Lz2Uhp#��@�;��л�z�]��BBXu�yY�hk��n����X�0�`��m�-���c���vd,���H�t�B�0�5"O���f"=�X���gM +��P�{#6�XH�	����_b"��љ�}ɵ�����ֱ�����F��\ڝev����{�����\�,�y�2�8�����d��7J��OYR�$y+���9u����Y�S��(.z�VaV�{p��:U�Q͂=/���!�X�*�)���а�ٟ�c��R�#�Z�p_k�KS�%���ʯq\/�(Z���0ƃ�K|����,�k��Κ�(&~:ts��>�X�����Er<���
a����>u��V����K�g�����[y��Qm��2�Has{$�b�"ij�>�rq��xM���mb/�o^2E�1��MF�)�kq#��<-�8#�H3߁m$����K����_ �������k�o��l�C:�RR8�w
���O/�q�g7,ҭ�[�[s|7`���	��Tvj%���P¬8��T�.(=��fa�2�2�ə|�_��hg��ؒ�������oB��`u�
�h�3yr�����]s~�[�R�G4T�= '��:��H���Tf�TMb�)
��[�@�E ��Pi	��8�iW��"��sJ��~��E���1q��kQL��l��Ν�Z��Z䕿4�w�!ŵ�qÜ��:��X�^I���܃��? � {"�=�HG��4��F��F/	��KV�~E���ڕ#�
��B;��Ҕy�BK�:�J����k��>F.t�/l)ţ ��h�o�DHh��]P*��g�?�Z!=&���5Q ޝ��B/*���9���R �5XӞ�}��_�a5�5���e-+S��,��?fS~��:��5!��;���-3(���xE�:M�7OqHb@��������S ��b���u-��
�۞Sԝ`�� �6
Suga���x��{�f'_hU%~/ �V�,���H�E(rf~7+��,��R���R�?cvǎ��T"*(�9"���{����u���GNM��X��0��&�d<�%�N��J)��	z��/Y*S���N�7�Fȸ�r��~�#��7a����UD��3m	 ���Qb�IAh���q+���)�k�wS��������d��l���s���0�=y���?N((��C:z����2�}#����X���eҽ�dJ���u�v �G9��^��hnO�F���,��RL1����![�*���h�=�%���wL����ӝ����V>�L�)M���f���>�W�F���O�z�pg���A�H��ˉ�V�&��5�^��6�?U�Twá�a����Ѝ��Zc����T��f�N��|�����[�����C�jS����	�Y��<�p�u�0n���@��
l��I�Ш2`�o�OP� L�#u.Fzh��~Le,at�|~�s!����a���˔-��W�"G ��D9&�@�����-Av��'��U��$����{v܌��斩Z���h9�I߈�mK[o�����H%څ: ������f���F%���*��T��y���v�<*�:ʃn='fLT�v�9��\9���$T]6����;�.�꒱6�� l�8�U(�L��U�����/C�*HI.I�	�M�����IҕL�t���c�)�E	q�i%ȖX��R|.!�f�Ƅ�g�v�]i����,Y���S���kG\31Zi~���%�A&������n��Y�!Gc�Է�y �� �7*����w��t��t2X��x�s��Tr	�Ӑ�Hv;���:���ot���Xr'ݬ�W�zt	�����>�Yv(Q��Q�5O�N�&�!G��1���lsw��:*���[h^�����$d����-�Uה\QĿ��Oh뺷.)��I�<��s��NIUy��@�5(�5�|�῜eM>�j�Z�(]{�j��\��V��So�>��|��$Y�Mj����)�������\�Pt]QK�,$N��a�x�Ɯ���>����[0I.�*��F.�罚��i��y�.�e�̱0Р:�*\�7�J� si�ێ������1P��՗�q��3����}�	� J˰�q�BL(�<�?u>%�"��.Zv`���tt�uݏ��X��Kp�Cy>�����	��*��夃�$��Sl������5��R��I05�c��>���L*�Hc� ����ZAx^S9�a�ЛG��f̙"V��

6	>�\�޽�2z�J���L5�m��(*�v���>�E-:��	Z)�����M��Bc�[���X4�tA�Pb��_3�SX���d͟��:o�Xf�,P�@�m��v� ��	�v6�.�2Q����j��y�tP5����Z��ٕ�4q�A�, �,���� )�	����:Ǌ�AA,�)n�k��b�港[�Z��D��l��f��e�\�L����X��p��I�p�����gE���x����qzp��i�>���:@`V�r����S���7���vk��p���]�K����	u�_�"�'��W�zU�?����s�X�/O1�"|�+���~W���s��%Ұ�VI6���w�מDc�RΌ��K�R4�1�#��s��7�{��NNj�դ��~������Ͼܬj�k�������o"vy6�sM����� �/�A�hhZpRg�_냳���U�Ζ� ̙����Β��ؔx>�6k������F����){��9-��GBV��n�{��&*J�u�Z`��p,
���W&�N/���ecP|X�0CB��J������e�ѫ�r_�E�����>�*�C�u���Ԥ��R�7�=B�����z��P��; �Q�%�k���ՀEg
��Lr�6�W#�k�a��I�i6��UZ����9���o�����ZN��?��jҬݩ���)b���*7��,xcٰG튴	U��Ճ�)Q/S��t����u����U���s�����y�_s}<�8��/�ږ|��WN�i~	�sq<�y'~�"e��y/�>��c�
�{�B�q���}4�vLs��<u�i9Ñ����D�zo�H`e�ܵZ"Z��R*�>_ۿu�I��i���.y<I�ʡ�b�â�d��+?/<G��y6�� �������'�ȕ�4���+�<�oQM�ꨠ xPH{G�6Kf"*�W��eا7�>wË¼RT2J�S�lm�G�cX�`5�F��4��cX,j�|$���fd.�Vn�ŏ���ǭ�1U�E�1�'0���P�ȗ
rN���@	LW��W8�ATA[X�&!���& r F��8+�����2�D]����#�����;��~�+W&m�4M�d	�ď"�Q5w|����-���ǽ�O�u�3ε�êP�K��{��h�N��\b9����3wr!z%4n}S#g���mrV�C�CR(H|?��m����j0X��:k�?�hY�u���g�����>�MYP 
��z
+�|���9�+!j^�)��ם�Q��L֎:J��PM�LLL��*8s,�M*�+L�ÿ����~k�b5����A�)�D9��z���	��O��<�ǯ��HO�Ll�(|守m)#-��Zl�d]���ses"@+5��\(<�'��0�{u�J�9r�9������R#�;JViu�"V�ܥD�M�����zg���ǰ�����y��OsKG��z��$v:mX�C���>~D�	"��t��#�)�ݬ�jfӗ~y��<�*+�~�2s8��7޼F�Fu�Gl�c����vLF��ѣ�@X���y�`Xm��~��ҚҜȧ$��.^�(��&r���y���p�nZ�R�w&f�a ѐT,��a��"�$�j��~�jm�i�o��\�R�K���	��f���:��U��+ό_Z���;d�K��T�&o5�'8;X0�l4@�S�l��BgZ�@�q���v6�u�Z�'�?Ks��m
��@ْ0���o����y�a�@wc,�SHU��֬t� 5�q��d����I��t�d�
�g���mQ�mp���a�v�@�{iW�;n����"z:�K^C�Y���IB0<;d&�k���\�t�)�&j�F	���?Pn�d��	@Y�������x��i�F&�;cQ�?�(��X2o����;���[tKh
�+Q-�� ��{}c9nn~��Ly�؀���M�)A�㣍�#$��L3D���榉q�]+�\$-Qu�0�yws�-N,Q斡\
tS��5�>�*$d\�9@�+��Y33�u� +>b'h�p��������gR|
�/����b�i��7]j��e�F\�d���u�,�����q\�'������5Pa���T�����D��& =	�F^��A�l�[�k73�M#F�.���{W�/${9�56F^.�F�ϸ�&�\�oK�W�U��cOhyٝ�L�VW兹���Y~�ѣ�hP���N���iu�n��q ����l�L����4�G9��gBɜ���a�,�_�\=�ل�D��-`�H�M�I ��`ulv�h��
U�@j�U�(��r�đő��?��_�U�D�]i��s>SG�J�,ۦS����+3����$�T
�&�̎�"�q�fTB6�d��������?l�Ã��@R��f�	[D���0掲�C� c��	�7x��7��ë��	qt��17)���b� ��:b���ak0�׺�`&Q�ϖ��E�)���[>.�jW%�$��$�m��>������q�(p��L8e�|I7���c�Q}�����@���w�6H��w�a�0zF�Fs��� Z	��p"�� �!�i�I��G��K[T=�˸�A%��` +�~�����E����zߩ�6�?�K6&�����Nq�Ea:5�޾�mq��~�7��x�N�z��������:�\iW4G�n@2t��Hf�T�Wād2�F��3�T��a��,�>S�>��5)���N�躺w�u�Yc���^���eŪc�p.
��	e핐���m�u7$�{ʍKl���s�>�n���Nu��Ehȩ�.���^�нS�|��1���H<��2U�9s,r���Jn-7cw���xS���R�<�I�j�xi�|����Fܑ��&Bn���3�2b��Y�e�]R����zx���j8�H�7�� ���Ncؗ���/�F�3�W�s�O鋚�?�Q?I�0ߜA��Ukl�pK��FZvtr������6�����?\�|�r�{��˅[�>idď���x��^�]x�'\%����$���/�\��G�=,<)��P.Mn�����S-/���2��#�l�xb� �����V{�pa�(����3f��{m�=1̃H��dsEY�+>�4�.�/ѳ�#0�fy�{�VX�!$����m@�E�]s�Ԋ{$�0V�0������s����kae�gdֈ̗���F� �[M��Wy�D(U���BE��QK�CO+vɏ�095Id��&�t��G�N"9�E'�a�s�=�K%�R7�#3c��q~��,���~��t���?�ӭ������J>��lT�!�ؓ�`���ӫ�%)�Ax�����=;�}��sMz�ؗ�YX�l]4�����SK"�)L�~��$����\v�T]����p�a{_~��"��CR�R쳾z5p�=L "3��<�k�fX��52����yer��{��?R�H��������y�K�R���!�Yr6�9C�j�3�LU��	~��w����b�b����)ސ�Gg�j���edX�Q��9������ t�R��twRV��P�et�&�`�Ѱ�!��HLiw'^�"&����Yx��&(3��sdW͈"|z���zB9j��>-Y��_���[��jK'��)���+��l�d;N�ǎ�I�x9�h��C�5�Ai�j�都�aG���j$���N�K��|̪����7�A�X's�� ���m�};�_@��!cާ�2KAa��7K�/��#N,Y����θp�8��P������֑��܂�w\���c��4��q��1Zn�=OXq��ʝ?zjJ!�.�~<�r�
B��t�g�@�k��ZB�>�Eh[�4v�f�M�jG��"�{�0��UP�,������L�z7A�i��-B����NV��:o腾Fs_���;��q��$`��������򁠭s	N�0F������zdɸ9��PQ�����
H�9i���ՃJ&���>�� كY~(�1�m�x�C�-69� ���K��z��l�#�@��{����4�SpqВ1}ϝZ��_h�X�n��E�0�Pq�H����`N��]Έo|0�����O(�d��*�FNƙ�8��)�[#�<���I�+�,�pe?�>�89����WV�67cM��p3����hF�Ye5���d�j�יt��e�fj��c���G�ӣ_���&jC�KF�%(:�㑙�b4�3�8�[P�W�Q��bp��,�G�>dO��[� <��*����?���NwG�