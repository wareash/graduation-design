��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jåا{�\�u�?߷�dn@6�zf��r������;,��o+�[��C�����B�V��_��/xL��q$S��s�TV�����xc]��>��:��A֌6N�y���8������[eֶ%���p/���wPH����������e�u�t���uo�k�jZ�x?��Qi�/yـ`C=�sYW�S��"]�R�L��(xerd� ��@N�ꚳN��D��@��G7%��[2�$T�fm��;���V���ҭ�f��甆f��~��<L߰5��fvnw���-T���K��c^4\Ts�'��s!�&�|��a����S�zY��PH#\�-'{Ҷ�	������D�ʟ�� �W*�p���>zG�TIka�2m��E\���Ą�ŭt����m�����XLu��l��E�D��Fk�tU�xᔧ�:���\K�����ӡdv�ۉ�Ҽ�g82�� {��BR������
�ԽF[�2�
��ʌI2B�i��Gw+��q�<�:��6���z\>ū��u�?���L��_�`&�b��ȴȱ�ݒ���8���[rh�ך~S)�r��5�0;���G���!�G�_���i���Z��� ځ�œ췬�&��0�J��S��h����>�V&\8�JNk�����){u?"i�y]�eg!�HS������7y{��*���� ������W䛘�%7ʥ�wK��C��x4YԛS��Y�<�y����"qпҬh����Ĺt����G`RrK������GdM+����l��>�i��j�V'��J�6JS���Sn��I�ᎇf\�v����d,n���3���U�C�fD��"@2n����Kõ�g�H�[3�7�Q[:rGY�GcP����,.ۿ���QP�?A�D����K6�G����j�>���Q's"N���{sf!%�f)�h���'��j˹�¥]�0�ͮ2n}�^����[�+�Y��B�e�z� �-A�'3����� 4\z��y��0ݠ$�r�V�@Ni��U>�Rᡰ���X3����7*�>L�#q_�W43!�Zb�&*~��*M<��OMwt�71��H�����N��dG��US=�O٥'���4��G�tT��y'`�+�-+����)+��+���{��-��/~��%i���q�a��D5�bՊ���fua�e���^ʹW�,j���Q�R	.�>��.>p�hG�۞$!�u�U�d�z�s��˚�E ���ӕ�[�MBk�?�""�y������T"r|��1m�\vNq��>=����>j9�׫�҉���,S�����Oc��X/��?1b����)���SM ��f
y����!KN9p���'c�n���\�C@3J��wI�If$S�MPέ��i��闟��f�N�=�8��q��2:�r��cM��p �fC����QOfq�X���%����P*Z&D�U�C�L��%��/w��wb���A>�Y]Q�� R�|2M���oO����;�he�.��ŕ�汹W�F�.���ChC5،�5�����`���bL�PL/3��{���N��Y[`�5���]���b�z�K������zL����٨~�����A�8��z�e��?�#�ᐏ���[[>+�+O}�h�$6GGI%A?܁�	��U�d|'bh�pS�e�ۑ<�Ԫ�q�K`�Ԣ��q'Y�4�.���d^h�+�Ԙ�>�K��)�wS�+k��i���b �a��R�)<��˒������a��xQL��,|���:vI:�r�|�#��]��?%���(ӧ�����; �� ��՗/�'�ɀ�p��֖E���]�x��*�j[_w�k�]Ӛ�z������`������1ƃ�r�Ӯ�EV�� }�/M��v��.������>�V�Z���ʺ"L/*Y5Kc��<u:Er�!l�G|����waM|�k%���b��{��B����Wx��Eѭ���c}Q&��ZYM�3�0ya""]�G9<�,ӝ����m~�z�l]^,�c�6�J\�|e������):ۮ���]p�gIH)Ѡ;C2��M� �6i����ӎ�꾬�W-.W��̀P���q��"��ZL��M�QR�\��	2 q��j�J�i�
J+AP���7�V�~B�c���2��,j>���ufQ)~���P�S��x|E��0�,���`���wa=�q��%�j�l~�4�ِ��G=]]�N�Jk��5x�}����2�(�y@�4�V�N�8�:Du�z�.��'Ce�B�P����q��E\mzE�~&wv�΁�W���C���D�	�O��W~2簨uj֤}�����/�2�Re�j-����I�?�J꣍�Xxx)B�jf��{_�`�H��4�|��9��2I�LZҘԻ�DZJd��W��<�l8��2A�T8��=-��k$���I��L��5�D��l���aP�Ht�d�a��<�(��� .u���@��^�k�Ē��`%K��������-ߔ/�{URt�A�b
���)Q�M�,���M���F������u�͵�*��f��TGlc�v����O�tC�gWa��݈�Y(�^OXo]iEBS���Y~���a���- t�����l�T�<dsoi	Ƃ��{+S��uz4�6(�
O[���D��b"�݈^��H �l�>��D�|�q�Î/���v�f�p������<�U)Oex������ɸ<P\�	t���,O���%Ը(��VG��({����'��6~7�k��k.�n�<��j��~� 
��S�ӬCO��L�&ʯ���x�	ɣ�ͭJ����g��-!F>.��:��HaHS��-7_t�����ĉ��L����]cmC�tc���M��+�M�Yy}
(�6.\����F1�?�����6k�j�9�G��P�:qE�;&�$䮱`>A%x!�z���T@�W;���"�G�U�W� bd��
A����*���t���o����@G�6~0?![W��nt2г��%�U�>�s�����r��\�In�Ӛ!��+hRy�	Ax1k0݈��(Ԧ9_���`������{�y	���wt��<�X8�@�����}s|o�����e�s�=kHq����ѐ[zd$ Z&�wx��z��\�{(��Х*"�;zw��9l��
j��cs�[�ր������cҮ�35�X�G�n�D�~��;<$qҨUuߴ�C �%q�ր~UlU���\_k�d)�W�%2� �����+��v����B���2�a�JZ"���P5J���%wYk������@\���ج�C��Ң�!��'�A��(���	\ΐ����*��V�;�7�9�Ҡ�ս�Ã͜Gy�6��C��o)v��Y���|��H0�� ���1��F�8�Z��Z�������,Չ5��=뿞�1D�+n�n�q���<� ���=�mz�]�1Ю��X��Z��䣳�[��g��m}ū�	R�N[	���ta�)��U�	n{b�b���u�㱿����*U����}J���`����
E@��Q��cO�jdq>���u!+&�0Nj#�q���ӛ�V\�H�Az��RF�9
	Z2q5�ģ(������-���1�Jlj%D�&�#�a�`�ͥ����N�~��6��"���R|�&|��o�����sG��QKü���Sﭢ&@����c��cd��X�tvF@~�T���C��(>]m0c�ga�.��) o/��8�|�b1�����.$�:����K�1c�*��$�i���o��=މ.�(G�e֑�(5�c9�ݫ�`e�O
K�ôM�i���^[���ޙ{�s��It_7�@_©2�%������Q�u5��_�����B,&N\���	����xwM)�nQ��,^��y3m"Iޣb�=;���o�z��(�y�qb�{������)�/v&+d��(b��r����DOD=zrIޏA�8���j(�O~���Xi�w���ay�3>��V�j�ǈ� ��H��T�%G�+W>����ߒ�n�U�� S])�ZڝG��b�������9p�zaD��=# 2��?�4���vfZ��ç� �Es�t�/<Y�3�M�N���q�:�s!���������)��C�5g�uo� в�
�ݼ���T���>���Z��O���]��[�v��W�H,�{��Q�!cE0�w���9� ��P [��p��`i�����=`�pNa��R���f7|���g�7��ɚ�^�e���@�=�iA�'Q��ޮ����Un{��tc%����W�n�Y�q��S���i�15]�A���I��'��tqk��!����;
d��[�QyNGv�2�O���};��O��TY c���D�9P�)��9�%Պf�Uw�5	�45霜pl9��+������zS�s�I\����KUMM�+� &dH�y�\»���C����t�p>+IT�O�b�!eVp�9K��(�V����ϣ�?�J.��얢�e��j��?-J�TK����,�!H�T��O�b��`��o����6�	w���nbyJ��������0����k�"ǫ鵩��r�s�=/	)��+��o_[X�o�Ν:``}߼�~�Bҭ�G�`��;���,�kTYד~�2���z�6�t�	>�6����dш���Dz@���⹠oܬ9V9`��.S��n�8)*Jt��D�R���buN�g�Ϊv�S5x�S���1g��p����94O)�آޕ _��҅�a��e�~�
��y�����|���3-!����xI��	��߂Y>�wps6�W��5��et��^ ��ue�b��7����ȅ�9�S��LdՔE��gio���Y�u�Pl�{��M�M�T��M��,uڤo_���`��E[���	A�@��e�D[/i?L�����*�� f�;�|Ź!q(��y�e�6��>P�mKM����=���w�Y 7��PP5tC�������*6�|�@I"`�Mאf�ϻͶ�˞���ߩb���[fͦ��b��	���uf:c�F��&";.Xj��gں3-�� �ѝxmh\f��������o�3홀��겼Ӂ���LQ�.���GE(iƒ��6=���n6�9�+T�/&")�<���;������'}��Fچ�U;��\ɲ�����f���S�t�Ĕ���@��m���<�{!�~�\�������+� ���v�=���H����2o>Y1�FΧ���KNq��0��v'��I�a�����ks����T��F��
�{ﶒ����^q��~ub�<g�u�-ڷEܐ\���~�t���)n֗$iO#�~���٤2X^�73CƤW�N�͇��qY;$��o�uF�7�����k�b�˩ن��Ι�@�V����a��}����qO�F����w�\�ue��ۿd�W�W{��	�D��K��!�*���)�yER�_t�ʭ�w SÜ�s�KT<�7����2���S}!1��_W ��2���qҪ�}�h�La�R������ ��{;����O�
��ʦ��.u���p>#gt)Q2¿;8�|�J/`=��g�!ܯEb��Da��S��~o��9S����k�M�
c;ٲg��,TA�?ǎ�L���!�jM��1�"��WJ裌b.���O;<ֿ��[0
�m�y�[�tb+3����z��p��V��L�t�^_��Mi�ac�&�'
�Ӏ+����C�
qXXwaO�u����j#z���r��h����ww�y6Ӏ��@���~u�E�RlG!��#��Q�uŮ��|H���ort��(�bzߋ�8����]CkP PS�=�+A�[�̴.�����)�����gb��84G'u�xK~���3\lE��+\t������(j��Ju9�9pU����DC@�:j-h&�ݭ�YBUv}�?ҡ�]��Ĵ'��U\��@�x%RM[�J�.7U �H��ʬ��4��HPn>�A��	@c�.B^n�KX
�R�!Z�DM�%�d���[�a%%٘��C�9h����8�
��-d��>�mz��{h�X�|��8���Q�����y�Tr����a�U�ء��B�r}�s��1J���]$rc�M����̦eyq�I��gW�GF�ۧ�k��b@���>��큅뗟��p7�,��гԌ"��*5m��p���/��	.ҟ=���Q�IĔ��;���ˑ�Wt)�x�o�y�'3�>�C�_p�G�pf�W�b��7�.��kx��7����tf�1	,�������tP
�"��X ��-)�R�k,�U%w��._���F�P�f��r�����!Ϫq�S�����|n`�H�D�l���8�,�VK��d���i��鞤����߻�`F4@������z��{Bөq�����̺{��B��#�I���v���Lnih�f%�z_���Y|-�:�fý�w�?ZG"F��qى�2H��p'u:ܛ��� f�VP����2-���e
l�Y.��:���Pd���y�@c�OR
���)��T_�~�O'�[4T!%f�׿�+������E7K���T*�� +	�[_^���@��Hs"�[^(~�c'�Ex��!���(h�e~lw�c�y-A>�!��B,�8��z}�~8v��@��̲�Q�c�p	�8����vbU�E2̉iɺa>�:w�}IN	���@C:���D8�>�B�[	�S���)�C��9�a��Y�w�)@��ڏA8k&`���'�	��$�� �m��vnIE>=ͷ�l�LT��g�[s�HQ�GI��7�GO���M�P�m?��>(�� ���E9?�Jq��?$(�~�|��[�=s=Ĺ88�@���	���)nvmw����o����!��<���|Z� uP9��րsf�0V�^
��r�^^?�CLߡ0[��auckO�`"½i���+�����F�M����=�/3."�u2�9Fץ��/��>��,�J:>�����/<�AU
�������2�t4M+���R¦n����q��5{6�' 7���؄-w:t~�GQ_�ŝh��~�����O��Ϯ�6n�3����$6ɮ�UV�|`B<��4@E}75Ykc��;|Q�x��<~���/��}4�m�ڮ#��ב�.8qI�p1�gԔ�@4�N�Jf�B�������L�T<���S�0U��k�ǘ��1<��y��^�w�߉�*���&$��sEw���];da����uĬ���ճ�(K'�j�qƸ�a��lXdI���9�.�-0s漓��w���d�
k���x��z���Q�����W���0W?���ځ��{<���H��<˔�p�cr3�1f�����?EVC#��Vϙ���Lx���sk(������ N��>��|�a�zv2e�7$�K�)���M�/ȗ02d}*����������C��������u�b��&C�sL��*'��d.�dq��;�29`�67@yc:�#�	������AC�J��L��p�wE�����WZ�
�Ή�s��}��5v���πS�������Zs�� p�#�̆<�.E� �.��2o�*�9� W囇�H�'��~)�E�vQ�B���Kl ax2mhZ�P�H��O �n�(6�i�V��):)��:��>�;�Q��&���)���V�+'Kj�m�P��<�f��uk��-��vB!"\*�}󛪏c�47�{��r��+������ J-�����WV���2Pാ�[M�M���%ϭR�ނ����7�1�pz�G+��JDL��@�6�4����|�H�L�&�z���͎;U����KbC�塟�L�&U�il1!Īq�|�",)�E�ۉP"�*8s���^��*�t�C)& `c�B��W-4�0-gz&{P��I#3Ɗ-�hj��JzV�%��;1n4�4��N��*\��M�Ĕ�^g�W����zh�I_~Wl
� �z��߆�w8�~�%�3��&��|{3�j�v.��d`��,�K4e�@(�I�f��������c��@����$��N[��(QDIvq��!5�A����YZx�-l>�ђ�����ʆ��W��yL�O�-��#�d�ϰ���nq'��u���x�����,D>��Q�Z�@����UZ,�ח��v�!4ݷ�́��cӥL�y`r*�vu7o nZ"�"�T��48��g,��/��#��5�:���y��?Z7�-N��(�����˾�#��D����@	}�v��7x��4W����ĕY���9֊2( �'��f�x�M�*&_�%�N��hƎ��m�R�GX��Qm���;R{��� 偯������Va��c	I;o��#;�@�����	h�������~�� �d�Z�Z�wB���<afV��Ɔ��6���)����/l��oh ��=�
�\��o�*!I��!(�=RgL�����"���a Fv�8ˇ�0�q@���v��L�Q'��<���%�Շm��;�o	b�Y�-ٽ�� ��txX �:Ȅx�"���]��E���Zۖ+�����]$v�6ș"�`���,��CD(7�bſ��_��U&Z�,�i��o
�wD�c�ɌR��$�셐z�<�r.�?Ib�����W�jV��静̻l��C{_�rxK3CRF�u80IT�g$���a]��z1����=v��d\�Cޞ�&@���/�����T�PgF�&$�J����2r&šQ��k �1��E*O��W����*x;�T$K� �ȫ(�d�TʢcIJ�˽���O\�ߛM�T�FG�론�����Ű�0�5~�<�d��w��"��5(��lL$:��N��P������4�zP��(���n��U�%��X���9~��,�/��7=a�Ƿ1C��1��QN<Lh㒧84��чHq�}yu�Vbdw]�<gH�����7�M
bs�j�6��σ �rف�h,>/�hh���i�
B!&��w!��i�<��]�nƎu�1�|�+��bkmkec�h�྽�6Q��H��^�]����y�,��N�W�h�e��:)�ˇʿ�yN�s�@s�(Įx!2�ܧ��uI��)l��|��q� S�_KS�ts]̠�?9a����b^�҅¢���HM<UM�鈋� �i���>�e�7}�O�k�Vc�ܓ��P'�y��DÑ��݋"L`��%���Y4���M�����X�yG���&[�nz�Cr��]8��b�^y<��7$�uW�]m�ߍ�����+���V�bB!c�s���������=��j7%a��B��ԧ2��:�vg*k�o���m_�Ma�+"���jö��rVGS�n��VE���?p�11`��/�+��^Ro���:$Nz���A��0�P���i$E��F���	�IK��ڴ�"�n��~�1�T�K�C���T���N�K+��<a_�fqP��교.�̷�.{�`m�w������Tь.&"Z���I5�vRm���W�ik8��=9��x-$�;��hIS��z��ơ�(�� 	�Dj���-A3�$t��Uv+0�1�����x�X�"�dAN��A�^��,�oFZz,�z�w_��w�~�qub�_�D�Y� �Nh�-���S �@�1�n)�	��>
��P���C� �[�6f:��3�w��ϖۘ�n�
"��4}��Q�g�M�=R��I��3�����Ŗ��6�9�.?, 8+g���uC��"�>k<��uX�ZJ$}�Q�A�*�9���&��N�C݅���'N&�����v�]Kp ��S܌@*44�H\���7��9Y��)�>����ˋ����j�[��Fg��7��n�-,��2�W;O^��y�^�XX�\ �T��?����
J��c�Z�c0;e���ڒ �i�ο9���+�b]��%HA�x�m���x2���C���:yw��f�,U���z'��5��U�!謣�yi��c���Ra .)"2�!U/B'�	�e��S�xT|8�S�5Ɨ���ԟu�]��uCsp��Ʀ�I�/��ƭ���r葲����
P	�7�y� ���B�+b5\�INԦj�![Ke�����s�Ԃ�؝���e[y�r��_���Ehn�=eZb����T��~K�����tl�1�$Dq���]SrU#�����."���ӏ9=sE�����|���7��P:���N�ԃ�wB��)�\�~���#y!Ҷ.�%�Gj�¨6����@��!�|�#�5���R9r�̲o�N]��	�C�O���_/��~�;�&O�u�����H���mT�8pMP>�/[%hS4�!��D��d��͍WRSx	zƔ�3���4w��F��m���!OVȈ�Z�_u��/�\װ�VE�A���o���@*�p��2Ԑ���	����[��9K]��x�\�b�ݦ�^��}��X������`���5t�� ]Ґ�TS�"�9�ؗQN�>�eg�􊴂�=�NEt�*v`�?��Ȅ���՛�8�]�)����.���(�!��)���C@��y��t��	����c��m䞎���7����W.+�p��kQX*�=�Y�� �~v�j���l���ڇ�Bs�Ul����.��By-����	����αo�lQ+�%F{l��Ա�m����6Iq~kwO�M��*y����O�@[��O�q�W���6�.*#TP^u��5�D����s�B�\%���I��w����A[&���/؛o�>��j�m�P�5��$pb��$��~��Ѭ�J,>��K״�}73�'U����qD�듽 �̝��'�/�w@��-$�X��z���6q�ęE;�=E%B?��e�)����+����M kH|0��`���9t�sݡ��BOA��9G��Ds����������
���3�jK��o�xg+%����*�t6�*:�CX����
Y��
��I�w�O�L��ZH����LEC-�ລ&��td4�������"���i,��u<�����{;r͞��>}��ã�k^҃Cȸ9���hS�q���F݊�/8���7ޕ���{�,	�A���Y�vݦ.e�(O�����=}?h[�!~b������4�w�a�����[ V2�D�l]��h�����v����D[~�X�Ǥ�9����H9�d�kb���m�*�Qm�yVRJ��%���{j�C��h/Nֻn�I }��|a���ۤS����R�ad�@�����f��T��5ݎ��n�CP�ZO��~z��,yM����D uh&:�7�Ӟ���ۥ�!&{����9�g0&�(��zM��1�t�6R}E��	3������|�~��y�H�!�� R�����]���pz`T3p��>������2��B�;~z�mc�o���-�?"�4ݣ����u�8"������/~zq�;C]�Z�2��z�&�sE9��B%�4����x������r�z\`8�@�DZ��?H��F�(}l�9���Q�_q>�T��x;�A�4��}��:7y?Kk����5��0
m	��<����&�#$$�r?�!�@����pSJA����3͘sx��bH{������m��預�#Ϗ���ȥ�sAQ�Ϊ����ŉ���>JP��'ژ��j�S!G���i8f�$��pMF���ԕ���vqU�c]]o����`_#���d�;�S��,�CɃ���Vb�R�Q�=&p�r̖Z�ތ̦o&�������?�1����{`!��N���xt{��A��?t�m�?�
2r\6,=.��yim�h�\_]A!�\�/_���b0�����8�z�$*8�U�����b�\��{�����h�0^�n ��l��5��콁�A��j;�0��ւF2AuU�QT�E�����C��6#�<��1���#�]���Ņ�j�9ֲ�/��C(�J)�.SX۴��Ք�4p��.G�{��]k�Z&��󧵹�t�>�v��i bx	*Tv��{�j�!V{u�8D"mq#.)�"�Pf�ʶ�u�\ }Ә4$��h�����'gAN	��w&í�7���G�O·�KI/�M�8Q�}��^�#�B;��p��8����!P*{O](�M��P����Z�pT�C���Zo=��x���J��J,{~�P	k�ϖ����
��Y�ݞJ�!6O�vY���J�O�A����A����:(r��`u�z�౯_��U0�/i�_QT5z+��[l
C�K����9��k��4?�:BGώ����ؔ����;���\~���-�Ǳy�;���		&I��O=r�W�{�.�d�r��q���*��~a�nNT��)Y`�&�8j��G4@R��#Ը� �x����������^���2�#�^��8Z���xb�A�K�&{GoՐ�/��љ}�%mJ�k���];�^F�K���9�8���/�9�<�`J����@ʣ�R�g���=\���������D���6����Z�{EUʆ`�j�������OW�n���]��Q�h�pj,I��ͪ1B0��t�
LR��K�`,�0fbэ�g�f3��q0�e#��\����x���8��:Έ,�j��vֈַ��|������vxH����
/I+��}~=Y�~9nU�u���N*���lC�a��ҙ�*��)���b�R\<_(�|�H��7$Jo�BK���,�LF�eq�>ǞXi�V�={!�-<K�k����'��� �	4*���F��)���F=�� AgB���s҅8����m���׷C4Tt�lM�!���uT߂�+��iء&ݰp� �7�><�v�W�"H�Um	2W)F��Lbm�g�������?0�OU��a���8�d������rC����+8Ҟ���s��i�j�DB����^�ûe�v����;���U�kv��9��'h���n��bri�<����DF�B:�i��
�����QY%������O�Z�WsA���xS��9�l�M�<�u�շcb'���U�өS�c��y�5m����W��{,W̽�F]��k�M�h���E,�Gm�I��].M�/�rjL1@S�di���JB�9��"�:�o���b�`I��;��F���l�W�dBxSq�����B9��H�2h���g�}�V�ZG��YN���R�r��X_e����5�k��ol޿+Ēj�Q�(�E��$;3�&�3`=	���j�\ɮK��d	�V�q׿(g��
8~���.���(�6z-z^h���7[��)Iw�N�I�u냕}�L�xA�șJ�H��RG]>#a�L�s:/<�@>�����IÝY�O��%͑�>��J�6�i��{��r��A[�TIY6ɷ�(��?�����Q
��C��+�<i�v!�]֖��Cy��[3x����B��9dbsZ�Y����J	�t�;@�1�N���+bø 1R@�tM��Bʀk؞ �~����:?e���hp�بv������-+q1�ls�y�zxXZ1!{2�����5(wyV�ۻ5Az����}�<���
�.
�=u+��ibsߢ2��j'u��37�L]�/w����!����ME��ݯ�37_�GZO�2F��}ґ,���\���?�`��~$�3G�(Q�v�/~�D����P ,����A�/ѝ�`��=����gW�N��\��&3R��i�t�|�ԭZ|�t����๥���~U6a�Hx�[s�r��H9�D7+���zd�B�/ ��؆�g2Tj��N��:\t��gM#L�c�Ȗ֧봌����z�TȀ\L�g���W��^�M�}�,Qj��Zʲ.jR����|bb�>0F}	�*��*���M�d�#ǟ� ��9�V�q�su�};w�"@��PT"@��p�[��YTD�B&x?�p�<>����p\b��q�����Q�Ҥ1@'��]�*�lHR����5�!+���vH�s��T�k=!3@����;]��?�ye_�!>�/l��o�#u��8,�UN#,��܇
�~<=���v��e%�͛�>�X:(5<+h�������	��1)�
��-4JN	:5~���{㜔 2�}�x�]6מ��,��~�m"J�X��|;��y�yq�[�r�#h�?�M�yuc r�(�-�j�?fSF{��P��EHn�@gW'��e������*c��a$`�R��9N��
$J�-�b�3��-���@��FZ���z�,�j�V�CEdo������^�0�
bjS��a.����
�5�{	��݄1k��B���>� �>t'�$l9\�$�1ZR���s�=V[����*)�-Mv���wNI.r�d�3%e�t>嵐t��Ea�=k��U�.?s�cB��cӧ`@/I���p�-}��wo��.�W�L�d9u�9�)����HOa��]Zr��y�{%(K�W�#+�Z�|�&?���w]�(��N������3�U,��"�;��nbJ<�:ihpc8O�3#����������i�S����[ަ�-	�P��>/���^��oG�-�%��})h�AO;Sc��c6�Q���:�\��b_p�T8�0	�5�r#ğ�w�3/�����$l?SVՁ�H��_�m8�ΕP�K�}�\$�=��|\��I2Z-��M6(���3YF�xr�#���Q�L�����%͇~j�ӑ�o:��Z{BH���Y�,}kg1�M!%;)���ه��s��$�)L��4Z�M8�@��p�0��QQu�φ}xr�\ÌC
|�[�ֲ��c��%]�3_F��'3�hr�`�>�������^$��t�e>ͻ�
ߘE�[�#�9D$��	w���qq\��ʳE�����z��B~�Ef綰�r#<���}��4��a�*���<1Rr��Ϣ�G[��6!������eK���j��p�8u�:3��9���d�����$H�_쥃V%o򦒥P�E���C�fM�d>�El�i�xI��[m�HZ6�a]���̄��U�j�inDT����vQ��n,���$��)��5�R�5i�E*%J^��@�$Xb6���bG���d�ֱ��x¾�p�&AԵgs#c4���pA����-ⷔS>H�䮛`p�iWW�F��"�*�q
�+˙�"����qT3a�����O8��Y�'V-�M��5:i��<ft중�OK�,�|^��p(����zy�o\Xʮ��x���O��'�;�Za������/��*O}��^	��<������9�N��B퇝���\7o������V�qK��x�LI�o%gW��vw�,��gJ��"�=fQ�/��x�J���(��(�v2f��D�Qc���c�mpQ�^��V}�0~q_���Ԡ�V�Q	��f�:e|d6�$?��/�C�h�o��θ�1Ģg�%njŪLz�&I@9�
D�q7��1E2"4�Ͱy�G�r�QGl����h��)�MV���M��ɚdC(| B�NE�x�e�r�Sr�G-�y��pr [Cf%}s�/��9��vH}�aӄW�H<�kT5��A~�ݲ�+�^���ӿ:������T�j��+�B�CX���l�y~�隸}�e�9P9-�����N��l� �Ɔ������
"�ׁ���)6ڃ���8�:A�ֿd<�~��$=����r=֊�0F���w�"ۓ��o�.�=�x]k�Hp���(��r���В��XHf�Q�q��K/fQ�^m�T�l��~�Χ�@9���ȃ8
kN5��51_k\��~A>l�n��#u�h:�lˏ�)�).k�v4c�x�����zMs������z4=H^��A�Aa�)\��ȩbս�t���z'T0(H�E�N�U�.ǽg�X6�(U��`�:��Ƈ���6��&S33���/�zݓ�I*>�� <�3#���^l�@����*p��.K���H�\��:�( W܋D�Vaq"��/8ZT�P�P��s/��f�'y���,~~{���]�5@������Ut�:k�)���*Y�d;]���@e&\�w̓}RM����<(��*}���D$X��_� D6��Lw�QF?��Ip�M�*#���d�綪l(RI�+�G���T!u<<�/<|���Wc���'A�b,2=7ťؠ )���cOɐ�N<4?y;��*��ůR"��pNz��U)�&9��Erl��r���6nI4���塚�����`'.c�#0"���x�~kKc��9NB.=w�/��Z"�b倃����A|���Z�"�X�A�K��g7u7Vzj	�xFp�y�KZxG��#P|���cP�	yr�:Z�qb���lU�������ٴH���Q�~Ŏ���72���=�t�$�u@�ǔ�$����j����V�g��3����8Mˑ�!x��M1:Z�X<�ac5w�
��ck���0�H߅ǹ�������!�C�4х��&�;��/��^S����t�cQn� �b�cJ�~G�5b�}�3%X��9v&�|�KEp���RH]T%��Aj~#JZ��W�ّ���Ws	n[����])�ko,v�
ˣ]<8��X%�ʖ����+䯸�Cf��=�i���R*�Y�8���d@�FI�x=��ڐ��|�veWFۜ*���<��n/k�c�h�JH�3����C�T�'���+u��"ܢ�Ə���U˪�T4q�1	;���;�`1nc{�|�j���]E�G}�#{�����2ʖc6z���qf��c����g<�3g[�i�.5'���l:/$#f�S�O� ��vG�I/pYWY��b�sw�]��i=���f�/�egiA���Xٙ�b�mXFǹ������+�Y�#/��[��MF�[f��O��kEğ���V"��g�Gߓ4��t�z�M�f�ݝmf��p
�����L��+��JY�ϳ^#�G	cՋ�BWj��Q/Y� Y־�����ġC�2~��R���#;W����=:��`D}R�-�j����m��b�[��?B`�g��[Ӏ��"}mU=�+���ߊ(�P���z��ˡ������m�
'%40eKT��.P�EE%���{8e�N#����Z���������B�i��m<���͌�)1Y�v�5`Z�&$��'�ە�z�:;����0j�X
���Vh$��A��u;��E�)�����.���ZM6�
`����l�+Z^���&7�X����h�i�x�\����Sb�MG��i�k6��aL�l�	�����t;��,�k�?+���zi�
�hP�5� �FLN�x0fm��|"�٪xW��?���!B�Ý��r�T�BH�Sߋa� J�Ԓ���|��p�
�WD7�ZFq�ޗ�ws���UP�#4�9&��/��6�����IuH�"�	������5M(�+�D+�z�7cd-��~1��1�|\�g���փa�U���ގ�eۚ��aH)���=�/�C��+?�)��y��Ma����v*���Cq�HG�<�<3yy��M��.B��K�a2�0��J���وy�W�s�c\I10���O��e�����'���rՁ[�U�m>�lXD�&n�7Է��?�ۥgO2�KB�sY$Wg����k͛H�$ ӎ��`X�g���zvY��(�ƨ���N��B-����^�qy���<\���1��ؼ��^�k�C��	e��~Ul��i����8����J���1�$�n*>A:���K��un�ϳb�ZƏC��aOQo~��"���I,io���Q&X�o�-��1[=���iYtSlL I_����-�����t�W�z84h�9�8�A���%��於��o����?��\Ǻ���4��B��_#��V�������Sz6�,C�F@w}�KL�M�����@.R��:����y�U���
��ϝ�Ҽp�o��H���L�OXz|^��tV-*\[n<ߴ��)���h%�Fg�e�]��s�5�&�U���/���j�b�=�K��ȣ�A93�	@))���v��1�?Ź����-�Vul@��!W�����-� �9�-����Y�����NM*��aֽHmf?hkI���	��^ ���>P���=�#X2���H$hLG d�Y��z���`�	ga�!B3��@���=(���nm$Y�q�iD�a�$�#Q�Us9?�<O��WNs��0v�P�n�$Y��{D?�a��[+zQ	���g!g����HB��32g\*�Ji�[6ͷ#�k���.�>'�d��j�U�=�C-�S#��tO��9'Q�'�r��&qL��$+B�L�ҧ��b����?m��c��S�E[딡�i�~>N���y��!ZÇ�3��	��$����M���X�|__�
~�����su�$!�w�ky2��j�e���P�/�� "�0�DR�]Y�zq�&o2���F-*�y��]�������Qrby^�Q��R�U;�i�#Ǐ���ﺸ�(� �^�20�
�̋O@]{��Ys2fW��?����ŏ��|�~����^�����'��.��%�:�+��%�y���o�������d��ՁwX7/SP_·�zyY��V���0a/-��w���J�ʤ����\O��J'~�x�Wg9��W�U���y�$�N��{�z0oY��N����KK)p���l&�4֡X&�Y�j��r��?�\_k�.��hōS���<� yD0@�c�v���!�:&2���3~���OV���2��	S�4���+�}���<
�M��@	���Ym(g�cB(Y#�{�f�RЛ�2 �N{G��WQJ()��\aB�LD��O�������� �=
�aT�����%��!��}��k�[����[9�s�W�H�&�p����pǎ8��U�1���̝6	��j��5�u����L��c�\Gi�3��#���A�c���t/d�2�����+<��P��]��	Iq��Q��l��m����P}��A��ipl�H�l�C^�k]G/Y��0a�����#Z���Rq��KD��6f������j6��(���F���	.!�
�08�t�4m�׍٠6e�;!P�N�lq��V^�v�C���`��wVOkRn$ ��,�fP���k���4��.��u�k�^f�����R���~���i7��.B�ʈ}�J�d�_�J\�����$(��3�Qט�A���`�\�)C�3]W�zF�(�)�x䧬yIo!"A2G}Pt)d�䀻Tr������'�/���z=���~m�R|I��tKX�\�G�`�4�h�d}i��eIg �[/qjS3��^rl�j���7�("�yu��@�_�6"��s��P�x�H"��Л�K�}%���Y3��){9�X�B��CT)�t��� l�%U �kXbs���Z���k4���/Y�jp&���,�ޤ�&@�\�)���=ݹ xDL�	$4B�@��-�
��uY�8�8�� R�OC��3 i�D镵�R�8.޺�*����7E7����&
l�pw`����=�_h��N�ܹ��H���P��lãg�m�� "0�;	�9���i�[ᰲ��-=�I��P�7=�mǻ�c�)����� �}Am���B=��ў����Ǜ�>��A���A3�܎�t�
�-��tj��R��U"��FM�l���8o�r��L^��8޿����-��'ʱ�Hԧ�7@g&��D��ɬđ9�"U��uڻ�%��h�C운�?�o����b�~ FC
J�OXE1�M����6ܷwQ?|���\_�4*�85��pk�l-uս���?y�ѯ@N��E�t�bX ���~\A����}�����!��KWwT�����X ` _�F=��a�rl�b8L�w��Pt�h�u��Xo?��b0����������3��t~ڃ�O�a"�kZ�Ru�8�c���3�~D����Ñ�*�����{~�VAM��b��[�^��ҵJǿD���ynuN,����}�=A� ��2R/�i���%;'���
FC���h��y��S���؋&�����~!��xۓ�ԧ�96�M��G徨����&���j���ogly�����f��-L���H�`�{�����D(�tï�⽁�O����i$�%�ޔ��(�^��^�I�����\�]���#�q�K�Y�W���(ی�15���
v f��E��Ú,��sIS�F�}T;��{��ђ` ����4v�?-���b���B7�ʖ�����.A˸��}�v�ؕ���O�TS-9��)�6+4����ջ�����FZ�a�<�U5dKh��W��#U}ا���X��c51ځ�hKn4�`��^���� UI������ߢ1�x� {���\�9*A2� ���4�ʐ	���*k�P�{�ݖ^��D_"1�l@y/���w�Z�+4˼.j+K��J��D��kKy��ׂ�7s8~v�Ԉ��&V{��f(�_��2���"�^�x�v+!��Ԡ�@��T��X��K�o��9��*E[�sm����Q�zx��;X��4�K�������s]��:)$1�*N�L�k�[k��SI�AA���S���_���T�alB�h�ڕ�p����c�͋yV��K`?�d�vh>�$�d|,$�D�9w�'WT�;	o,o��D�U����zm�.peH]�q���O|�R�w^ȕ�ۗ^
��Z�Fy>FY�@�.�E�m�Ű��+�����$�0�J��"	�,���	dZэ)o���K6h���w�싉������sٻ#)l�y�W	N�|�?.�Q<_fU��pZ��)�p����Eexi�o}�ժm]~�3��N(�d9�]K�E�`r&�����y����\*9F �xڽp@����v&����㗀v���Y�,���O��Q���OH��X�s���͒:�H7l��b��'J��7���f)v����K��]#S4���B�j���[���sF�?����𔗼�b�.�Y�5�P1u������?=Y&& ���9�X'��R�2B&:JQqP��֌QF�xI �$��N�F���{L��F�I�/E�q�=�>H�g�l<`�o�m�?h��$`��Bm*�(-��^q�x��}]~��7��u�l{���q6RѮw�^x��{�Հ�kNbf�������ؚח�90��?	9�ۄ��Rim;�%��_}�^�~b�2��])! �z���ةRc0��H$�ڞT<P��G�b�gT���e���^���4��W�&K,�O�,?���o'��e�zĤ��k���?����y�U� 6��Ç����FK!4� ���8N��L�m�h"1�I4��2�&!��x�+��d���4.{`Q^��;
�x��H�v��vh��@���M�����֮���d�����*� ���!��(Md�کKXT����q�i��(?A���qo�[NA-0q��!Rǣm #���a���*j����Y(�@^�j91B�$��̔�����.L�{/�0�B=۰����*-L|��Ye��o
[ze-2Ϫ��?4P�^Pnq~~���KD�	����E�V�(����� g�rGuqI�Y�����1��ix8,���,�@;�	�TN����Os+�%\Es���C_������C$�n�3mb!��s��T�m�)��I�L���K�$X�)�˥=��o���|��t���5DBw� ~��H�m�Km�rh�Z��T�V�U�/G��TC�Ff���e!7��4�)�֨=<��Dm�G(���~v[ެ���B�3驵�Ѽ�P p�b~��Ui��\u�^���=�crp&s_#�h��G"�1�'$�{&Ns�
>��a��L����M��y��A�ygND�v��.��: /V2
��8:g���.�Fs袧&U��/�����wЊ*��%9�y �9*��y\�r�N�&�y��WԺ��{�`|��%F���$������^�Yh  �A0�P{����t����h܊��@�[�ʬ ��ST�r�����Ԝm�D�� ��.�����u��l=�$ ;ԥ�T�B?	�Gim��e#6#�g������ׇ[Flo�EsL��w�|傹n�����_��>�k��3s����$, ��b;K���E�����`�|	n�uhp�6�;� c���S��� 'ܬ!����-_ �C�4̧�\��ىȥQ�c�)��Bh���㢎s6���,$�0]!���*w'�<O�a���58ٓ篕Z��jS��x��J�ϔ�k����Nu�h�׈
�50t��ϡ�qq�cn'�[Z��6LK�y�x���~H��Ln��}2E�H�Eb�_�}���GW�44��=\GΪ��b�T_��P�w�vKi*�3{|��K���}�^��Wж��3�A<N>�L=���'���M��0� A
ݡ���8e��O�QVG���ѥ��:�_xS��B�-�u�����%���x�������Y�H�Q�ґ �/ή]���~��2WO'�Js�<`�v.deΕ=c�	����&�ɼQ����ф;c�1w`W�}P6B����b�X�*��q_#����[Ѡ���V>N޺)V&��&'29�ʐ���K�b��!��'XK�*%��޾E+����5Cg�*i|�ℹXy�ܞr?��E1"��XD��n�I}/'�c
�}Ճ���_�-�9�YB7�6~�-'FzQ�nֽ���-f@nv}r���]Z����Z�I�R=��ھ�FJ�w�� J�Xë��bГ+��f��J��g�wbD;����jU#�a���vX��Z>����`i~'G�J�U'�~u����-	��ws"|[�3�����;�������xO�o�8�l�2��C[��~�U�����+���7=���Ƥ��o����5w@�\u\�Sꒆ��B��޷�S�6���%�����V_����� ����y���rP���ѩ�
頃�����%� Q˩[S�e�B��栏 �C��K����y1��EԬN:�X����s�^���`�[�/��o��o��p��0
U������ɖ��%!a���1�A�5�;�q�YW�A�*�,Y�����L��w�j�X�����l�1���ǜms�3�RވeH&���/����K:�daĹ�?"�� �$��j!a7��㯋�ą㐬��a�$k��:�l�9�q�\���DBhPk�AT��]�[��m^g ���KȢ��yd�� Dı��$���Q5YL�j�	w젱f�Q�b�$o�Ĝ��Kt���B*S�<S���qԣ���u�vC'�76I����IѺ��SkЄ����Po�X&oklL��@?�
V�2`͹���>kttcGN���/�8B$n�$4w	���;/�[�w��͂�5���#:h�1\��XA��ez2����|��G{������~���Y�jбAx�RZj�-��u��"�x��Ik#��P����y͎׳���HA(g�aB�z|���^�����u���$��7Sq{��6���g 	� }���j�9L�eb���]0������?�����[1�N4���NU�C��k3�m�z��1_�X��GF�v|ʞ�}B�P�	k�`��w�/��������7��l�9>�͎5A�����p������|t�@3Ҭ�0����d�8k�λ0ک/&��*E����Q�t�Y|:��[�����H��/��c�4HX�9��=B��?���IG�쥌�Hŷ�S��"��!�o�ŏ�L~7�>g��<#���]���Ou)`|D�e�*ǯ�ڹo�t�5���vsd%�7���;��B���%��!H�io������B0��,�j����j���i�:+C�1��l1�?�ގ��PE�����f�t���La"�!?
����.�̶ra��%�e����H��98�n��Sk:A}貶g^
�ΟV�������c�g :ǀW�	�<�`�4y�p���M[�Ś�d�����|�WR�3����
�A&\{���	gzw��l�.�O�;�lmȥ������7�&#	�q�تΓ(�ҕ�%-U�d�̨����8��z|�;�9�Z�Xhh����'E�O-Y�8F�	#�\�'#�w�~h��b��H�PL�!��W���q��1�����s GՆ[t�Ñ��2L����Q��M�hM�=;l����D�c�j6�UlOŢ���Q�S��`���10��u�D#��3��w�����"m�B�#�x��
3M$�ރ��[�Q��=,�R�p9��d��d6>x��xRuea�F
VQ���9�ZU-��'�q<7��9,��_i��{�ݙ�^�d�s�"����9�e'�R��w��h��
B�?�N6�:h	Ѷ��A��ER��:i��[����1�t��
%�Z��~ �rV31E(����r�ކE����t�쩦T K�u-�)�o�������M�H�&��խ����h�o��s�Շ�� dg��
�5:(bB)� v�4)���McFKNL��B�xI�M=�7k���e�w����[0*��Q�F�C���_0�c�v!�N�]f�����m��C$�~��Y���;+�g@n�W�2�+����v���;r�M(׭!�9���]����bdES44x��b�O(��657u��Hm���d��7����q<��v͉`��Әe�݌@�Mb��A4{4ɒ��V�������T�ʜg���e]�0��X��'��Wҥ��x�jI?�MH����ۂ/b���xO�	���Q5F�R_&#��&AM�٩�X{�ɅqX�h@t���F��Ԥ>OL��Uf�|�e\�^����=0��?�A lV��se��v"a�"�3�UT9�����*�L�!��~XU=�˒��ؔ_˒׶�I�=܍�Y�G��D0*�u�,i�&���^�Lι��p���7'G�>E.�z^�W�3����@�E�����e�}ɾ���Mt��&�W�}b�z�l�5�s^[z��<ر�~=�@�*?Du�E]�C%��v�kvvʟ0��������^��Q�QDvq�����#U.��_d�a�r����
u�l�%�p	~ψE3_�|��xU�"���u���(d��iQ���U�-�
�l1}.ʞ�D�P�;�U���
)�
p+�G,91^&6'Ж�s�Vy�u��WFgƩ�mb���~pL%��o�$�����~|��� �$�P�+�Z�8~��k����&�����6V��0�Ήc)dXe�J��~�HQ`��_�Ѫ�9�^���}څj����DM�H��H�8���ڄ��
��oVNZ�E;��w[�p�ϗ1pF��j��GW�W�����~�Y���cx@��K)ަ�x�]C�'!|�������pث��^�U����wͨ�-gk�8����h�mY�*Г����3[�z~'8K+ȾR����>�>�֫��~
$��[��߬�)q����S��q�$�?�j,C�JB���{���ɰ	����B?�vI,�����  �@(���b@�3�)'��]%�G�.�!��(��3<�"�j����OI��/;Pn�V�Pt%�v�q(=:L9�$=[i��iD$w���l6(�n�VG������q��/]j�Ux�ؑ�w��RF�st���n�<�G�H��1$�qW�R��*�E�^Q'x�(4B�o�h��,��o1-)l�;�0dj =� \��H�73���]x7w?X`�iu��!�Y��Vf7���Ea/�˵$6`4E&9$X�@D�y@+�Y���J]�@�6��T	ή�w��hEZ��)�re�+���VZ.{5v��J�v]��m�PA�A��݆(+D��o��e�����=j���b!8,7 ��N��c4��5�T�<L&Z+�i�;�é$��j��_	��.g�:zY�1髇�}����74�(�z�5я��L��ݍ���4l�O ��A�T���1h,x�?֜t_2�}s��ў{���l����#Ο��"�:��~Ǌ�n�m7ˬu�
�۵�<b�z uj������o��oRì�?6媺+�^��a.�m+�G�j4�Q3_x����eg�w㴽W�ܹ3���:�ٻ��:sGiTbs۩N�ӟ���p �($ՖgV�R� �q";���X���[��LW3ji����ń��P�;�	��K)_�M��R�F��(y�W��S:-�����{Z��~��[�d�pӮ7;~�
)�#����_�,�T����8M��7n ~6�x����E����3�����55Œ�p�Z��|)+.��]�,��>	��7z��q�
v��S|nNÞo���u�Eb�u-�W�8��<ơ	c�熃���t �EG�z��#���MR\_���-��Z��S�̤��(:]�J��UL�_m���̴]'���Рq\t H�!�f'�����J2�A<b�U���V�٩��d�~�D(H��P��1�=��ȫ|]u�k��f��U��.�S���0"ŵj�	���n���ǡ����ω��Y<�N�Ѭ��_I�|�0�s��U���L	s��H�9b!� �bb&�S���ھ���Ԅ1��0Ș��C����ۃmY��6�ђ�ѝ|3�-׈�ȸ��ԛVQ��5�nƼ��r�,�|&��"�ȚMs���ZAGX�B*�S�R��~W�T��q�E�g�쯕�%��t�w�k��"r��w��l�^��Fk�'��jʾQ�p�}Y���.iq�YG�i�g)��AG������4�[xe��C�^2עU0 ����]�z'ct� �&�F�3�b%1w�4�B ����R��Zn�׶�v퇇�O�����d�j#�@9��+a��?OGg!4����͐�a�<�f�D�8G������gE����E��_N�xZN�m��+G��� ^țx~d��X�ޜC�Ğ#��q��o;!��t·3�Çkgc�j�bW�AM����ڷ��p�;�X
��v�0.o���F�s����V��as�{�:iH�>��଱jM���������k��U��gN�.b�:�>d�z�u������P_��$�1��a��e7�-�P��v�z$�P��&���%�TG!󯍧〮u�L�ϟ�B'�9c/��}DT�|HW!��MW�'�n|$v }�!3��.@���hbUz�]I����-�� �g��2�x��\0��7���!Q܈F��,=ل��jY���e��)�%��;U�ds������E�AVV9X�"�� �%���^�r�$ގ2
;Czy�Y�6*�#��&"��Y[F��)��<�k�}>A'�ڻ`V1�R٥���g���{���E 7j�y��?0,�|_�,��U�q��	��L�~�&�X�9��G%����ѣw~)2� y��Ö�0�lZ���g3b�<�'V�_���L�G�u%eX-��sFI̼��F�
(�8:���W�n����"��
�!�BAם��E�s��b+�伂�V���!>�*��H��Wu,���C�\hL�&c�|f1i��΢f��TE���H�\Ώܹc)��<�`��_���B�N��c�ʻ6�nǺ�y�q��a��kY��k�$k.�^f���P?���iv(H�&�]8u�r�r��/t*��*<%K�4���u�q�9��J����A�/'�)���i��A+��P?ӡ|�g��4��u��/fƕ��N��YI�3����訑�L��:�V
`O;D��og|�2���< [�#�$�p���D�FɨR��d�5��� �{��};�w��q���Z�}��_#����p���.+�M�R�漠D����b�ț�:m�p(6pSM��[&��b�Y���f�@Q��4�KI�h�!=-���O%��%�o!�	Z�^=�S���d7����|��g^h��r�r0���|P׍zA|׆�mǓ3�s��U\���E7���{7�詒J�]U�?�Y�H
'�eMQ<�7���v��煉�r��=�S��9[��x���%s���9�U���J ]��K� .U_[�|��:굨�ˊIyi��_�~�1��_iQ�k��P�23��f�|���C҉u �ǚ�kZ�i/g��_�o,�7h��˶D�{勰8W:�j��;�r������aX��]P��<�o�D�W��vMJ�)l^��vA���#,sm��K�]�O��jF�:--;����<|��t;�U�è{W��?I���,X}�#���ò@~:�/�'Ye!`�P�����f��)g
�d�09�X�۠���K+��z�C�8S�qUӤ�DH��n:�y�x0�1�����A����(zWW��/y� 1��^����e��:*����7b��p��.&����V���	e����}�̲�`�����:Skb��KU�a��ey/�#���#���U�AA��Ơg�L?���G��ndb��sRQ%)�5�;բ�`�y���V��lӽO��1T�	�$o��}
w"����_���z*2���S���!�/Z��]?�A�x]&a�\Y����}mlS瞶��v�xp"#{
;@����|-a����x>��h~?0�%Ŭ`�f�~+�S%^�6�M���oEDi"l(�U��8�x.[��#0�>6dAq�Px6'��X��Hݯ��8�[��M@7[��Y ���#�	�`�X�Df�Zx����AHG1kB`�_�l<���2�0ho�.yI�]w��H�wϣA�d�M��T�\.�%�-�kg��O�E*hʚ�*��e���Ʉ��Y+t���THV<�*R�O>Շ�6�~~�qV����e�͛���n{�c�y�Lı��wOtbUs?��� ��-G2���!����Ɉ��:��T�|�_��ND,"�h��,<6�2>���J�/�Oh�YQ� �&��sX���m���;K���G���	3�����i6b������ޱQ�8=L2d��� S�vabK�* ֔�� {���%K�X�#r\��f����C"�<?�����h�{���7"�L� �ۜ�+�n(�������û��
2�6�X�v���9���<�O���~������ˣ����~��eG������]!~�K\�w8:���E���ߟs��P`���?/������)L/;\K<DI�A{��nXV`���n�="��u�-C�$���<�g�Lv����J�S#�}��Hx���: �m�Hk�W�0_�{y��|� [ײ݆M��bQ`�<���6��C�RQ��~���,I��Df>�;Y�����Y�b|�Vd�#���{�a��NX6$�����5��'d��
G5$��,4�K���M���\
�&x����nб��ɴ,;oSn���� �J��M\a����/d�7-Z��Y�v`z�wO�Skg
�2�f(��/��y�n�$�v�c�C=����m(h����s�υNZN�l���7'\e8��,��:�
&#��Y��	�2��U�� 4(M��= "�'«Q�[�y��{i<=�J�;Xn����X��A17h��'A�Ci�jn���u�A�Ƙ���yp��.b��(�(��o�V��+��5�'3�ߦ=#�+-ASK�ئ���-*�����\Z�W�hъ�q���"�G��o2���H�|��|��`��.#������K��o��~��Ө�����"��WS�Q�,n��6S����y\����6�?,\��y�K��+����܃u��\P�4nq���sq.	"j�����O$^�\�w.��x-x9�Q�p�!cR��	�zv�^���!,�K].���`MЅ��Bdф|�l�9��H^��%�n�'��Ut�b�)�'e�FV�����$|��H���\O9g�]]n��Z�@�C�.���`���˚ظ�~Nt�6���(e�><+��s�JM�������$HF�~͢�J����9F|��p5�-rbn
�Ez�V���� 4�$��}KFZP�Jܩ'H?���69eL��?�B�u���DB���'��M Cd��2ϡ�N%-������	�����5���ǅ��r���7�Ř���Y�v���������a0�V�4}��A.���%k�8$� r���`B��P�$L��wB�Y���v��}�zPq���to�4�ME�ap�Il\����[C|��r�ۃ�\n���������E՘)Β٨�@8y�'�I
��~9�\��Yf�e��ÓH]���d��ޞ��`S�d��rd�������9Z0�,+�ZK��}��t��,���Ѻ�邲����MՕ�+�I�uhM/A_� !"���b�8kkT�@O���dXz���y�8ۘ
1�kت��QV&��t��8�fL�8C}ye$_��%Æ�i�q�<�w<�2����K	�SsVJ"nR���"�D�Y_=N�T`8���cq<b��/�\��0�1��O�(~A��Q��o0�����<L�#�|�LI�P��&4 7l��W� foDt�8"�=����I����7q�u���`rzi��;6�t�.��)!�����sazw{�� -�u��u��+���������d��ٰ���Ei ��ﰯ����Q�☥N�4߶�Axp��%4�/8��Ь�J?�Ȼ�x�8C��#�OD�z�|��C��%j~klȎOi%``�^[�;jI9�z��)B����&PBr
�����/'d=J�q��g$e�&=����f7���wݩrʁ^�Ww쭨hH��Ԝ�*�F��5��+���`�rͅͷ����Q;���V w?����za���\�wi~X�������Óu���j�֢���m�l�쒣NYe�r��QkW�	��_[>����xeEw�?��u�y�7�� ��@5�Gd'�O\7x� �lH����#���~�四��K��_;��C%Tt8��i�&�\�����>_��Ք��j/��_�������?#��f�)ZT������⁉�$��fv� 1c᫼b��	��� ��*�u#M��J�P��5t�JR (HPG_�Ol����Ï&�m�͍'uz�#ݱ�q�d@_�@��s�8�<j���-˴b�lPU[ᑹꃦ�Fe�C�7}~���3���|�X��+��Dm���4��Wu1�ʳ���D�֒��sؔ1�E~� j'!:�E*�Xg����M���ߋ?�6�,i�y"_�7I��!�+w���
;�@�ڎ[�tj��gɅ.��ɏ�@N�V��|�a��/��~v�j֋7~�� Mr>��5"}⟪n����׫�CY�t�Y)cA��)|D�t�MW�{���m$X�d�ە�$�p|Zn��GJa�Xl�XE"�$���x�HQ�̏��&���C`�d�}�O����
��c�^ ��n�4�%��|ʇ��p��	(
�f�eƵ�B8ц�*S���e�L�$���Ὢ�,�j:���͹���I�����xi4�!�S�������u����Vo�O-���^������K�H�e
6I�K��A�X�dj��6/�W�+��e�>�k�͍6@]�=-�#�S��2�$���@�X犀-8]7/r�:�kA�t�d�])c(�7>��ȢK"	�>�J�n�6���e�ZwLO�APQ�>��_�U�+/���Қ��D`t4ygӨ�G(V�邟gmQ���+¯ǈ��:�6�h��Ϙ��̻���"i��\��^�&��S�������w�JI��� 9��e^b�-���=|k4�ԛ���N�e>Y��H�5h -cT������)~P�"^����'�Tv���6�˪���Dʍ��P��K�]���3�	����z����nI��ԕCI��sk���I6M��tKrT��2�A�3ܚ˿(��K�k�L����s�@S�ej�����$4$�V��3O�Pˠ�~���kkDo[���7)H�����`a��1��@Mf��@F�B���;����I=oO��Eka�Oo��I���9D��ς�����$#%��f^.E�r;ᦋcP��(
iE҇������G�G܍�Ҝ�O�}�LͶ�������n�3��j��ht횒p���ʍ���r�9��L�,�se�s%���aC!Q(}%<�n���s�\>n��L�x��l52�|��6ww����r0�O*�6A���c+���m��k;��0���E��D���~�&"�{���eߵ2k�-4��)���V3w����?�e����<� ��N�#��LK�E���S���{���Y����a��{��!h@�{z�n��f�&����X�ޮ����Ы��J�[���S�]���a/B�uS7l_[h��:�С�E�=�E����	��lUs��2j������:#PXЃDO��A�٢�]���	ǎ�K�_D�
O�w��k��@�k�a��%�ӜN�F+F�_ ���B:�u_q��� �殕4����/��bߪ}-�h p�%$&{F���Yx��N���4��TF+�&��E�>�2<�y�%=��R��u�Q���0=���R�����.�T9\7����4-��A޼�?U �I�E�_�N�bC�ڀ#��|n46�1&ԠĦ�E���wV�A�R.c�f�+W�P�URWx�?����g/�s;���-1g��~���j�1�,���z{�.�I��\;&�ۮi����w,t΀]�]�� 5 M�/.�6wB���e�mH�MT�GW��bW���`>�{�ϵJνY�jVV�ۓ�P�����(�u;�:�ޮӔ�D��4@a$�� ��p��FG��y�l��J5�2� �wv��"!q�U�b0��F�|����Z%��Z��os����?#���I�)Gw�@z1ĕ��L�(�"���7��
̱��70R�X�	4�U����W��eGl�_ �`�@�s/pG�~ �+�t�"R��p0>�.��n���<�Gj~�M��ŋ�m&�4���H�����k��#_d�o%����ăi��E+�Y���)K�f�ٻ	�Y2z<o#*S^jz9(jx0�M��ŀ�Po
ptce�_�}��L������[�k"��Ԍ ���z`����u���
��hW��3�^ʄ��=�#
���m ����H�:�Ě�S��"K\a4�C�a?�{�e��)���bh��R/������1�c[ï
�}j8 ���$c����-ߢ��8(٣�)�%OpD��H)ڎ1�W��[eB�V�3Ȣ���~`K�A);����C�櫐d��Ħ��^{[��m�� j�3��qQ�����?��K+���cMQ@sCt�s����̨�C|CB���BLaq�Lu\~oW�	�7΀$F�� ��:>�-����]����)�\�j�Y�B������ �@qz��P�xYf~��K��\�k^t�U�Ⱈ�OvG�^��g1L@�K�g�9��쓙�e��.��=�%��L]k�J^�¼Րp*0�Ч^���]|^�5_�'��n�5	�u�U��9�?���Yj����wd�<c���8�E�,�2�=�y���(Fa��z�UV��.�ϙ�ve�-�o�%*wϟk�g�0�
�T���J�m��
�x�Y�:X�W�Q� L�ђsk���o�W[;��U�|r���v�v��3�v�-DM`�ߔ;V�a\�=��j�G�9�Z��a��@'�9?"����6���	;es�����2*,�����z���L�4(�#�ـ3���OPA������X(��`<������}�u��QLو�n��Z[�^�L�E��1��OH��i����7��H�A�9��ވ���R�~&��U�\9�0�c!x����N��"?YR6[��b�W藨���.�1��������\::�xX��k��i�'A&�O{ �����h2Gm�P�8h�i��t�����%�����5��r�-*#�ŵ����.FR��r���2r���v�r����<R�
6�~{[MLڀ9��U�z�T���G�ɘ�[���}7��	���C�z�F��=�"*{S�](@���1	d�S
4�VP��s��5-P��Eǵy�EP��EJ��.Z�\.(�`���`gx�z���R�eL��>_��$0epǯ9bx�
߃%�<�~>W��'f����HpW���0����2f��IE1��NI�*N��Y�*�|pf+�=y!GTtYP1�ڬ�k������̦�*�5]㎹�������%p�-��������c~v9ٻַf՞g�h�m"��v?(q�AzTAW��6���&�Yc��$���b��z��P��rd���JXi�r��+X�������h�j`J�E 5/�3�+ �<��������&'�e��x�t�>��L��S���	�J>�{gk�7XONX�t���맪�y�!�S��G��q��[]�+R��F=�C���� �vx����fy��=h����^�լ{��Ȓ��޿�/r���/�ᦕ�Į�$�a��4|���y](uԯߛd�O�[*���t8Q>��R�;�M�R�͒��޴��9XE���V� �L�խ���]������wQ�s.X�ť畏X( `������9����
��l9{�	^x��1$��q�����ZJ �2fCr#$���'���)��>���:0�QڇMcr�/�ԙUg=���q��d�� (�{8��r�M25��[�g��0G3p�p́�h��Y�̜�r�{��q��k�s`�$�L*�BIaХ �_)�AB�@p>T��SoF�
!��d�*,�TҵKٔxO��É���Zq�-�z�
�4�#�.�S��5��p�	����3ϕs��/#��`�{�ɖ� l&��H���"{�h��r���LR`2рq���V�y?E)Q9�{a� �G�K�6x<`��ȩ3r��#}
�U�Y�F� ��G%�q�/́q�KE�$��>%)�h3��2C<�[g�>ij�Y�'}2B�|��:ZAS�N��U~k�S���9$Au��h :����?��~�����>��9.���E@��V8��cA�AHC��U�<��w�:u�)¡����{�j�끞m7�8�B
H ����&���$��	��U�L1t�#٭��w��*u����Ce�0�Nh�Ce/�y"�:t��q�l5Q�q�z#����X4��,���~.�C�Y7�z@�<aI�б4,�m�{��s�H�:����=��n\�!A��2�x��829G�^o׎�ഞ3��0J�O���h� �����(��gE�5qݑ�;�*�G�q�B�^���p�g�P����af�_(�(��Ǻ��x\߸2l�_%��zUff��a��d*i�����C�Re!�%�9�-�NA٧�����%N�%	��dէD`����a�Gd��M�y��.�E3\�$1V�/�:����-Aa}�>~(w�m6��6I��#qa�斮�C�iNU���bֱ�^�ڦ�3ՊR�!�/vF�RT�J|_��sE�b7"l4�P��E�	�RC�QU�H�:0�R��w���~��{�;�1��n���L�m_ k�2=����|�JcH��)H$Z)��	�;2oS���9���&�Am�!�kj%O�ƏG-�p�����W�?"���`wݣ���G���k��7%T'�Z��t�C�������s��H	W!*D瓼K.S6�l���$d���U�sZ0�;AZ�����b��{��Z��X�uܛ�z��R�*�G|�Sh��QŸ���uK�G?�gۇ��0R��J��2����l�*x�X	6�0_����f!��H_�im��݂�P��ʋB�{�󲙇�A�¬�M�,��ų��w�5_R�}Ŀ�S����B�
�	��@��VR�u$\��࿻�<�\��O�-M��|�ϔ*��W��p�v��	����v�8��<A5�_	Z�}2����E��S��Ha�̕����)�ͽ^���+� F"!sh	(���l�)Ƈ*�8|Ƃ�߶笲 �j�?��b@"7�r4�i�,��吸��. ���s�$a��|,�N���8�ؖ����cޭ��,�f�tB�?s̏׫�L�<���.���&O_j7�Sm.���]�1m�b�
�2��!ts�כ�kk��2���p��Ol?�f%�g��o��kK��	�Ջ�Ola˞D1�6�����J�D�����b��ut��`봹X���P5��;�3�c8�$)��冾��!܆�� �eoX��h��h��ђ9��H�=#���G�/"��c6�f�vO�]g ��G������l�VS�P�)U�>H��?4n��
���}�귰7_Uf��\~��{���]�R���Ft7�tK1ɡ���a:�(afj���D�uH�����R{A>0�4ƥ�]�^�� )4�YՂC��3g�����R@"~��:S��Z\'Z�WK���UD�t��FF@���
+�&�#�z#��]"�&в��|Z�)D���9Xj�=�_;?���>�9O�%�����a��R�~i�@��{4d��dҍ�� �-�r������!�,1�D)�Kޢ�}��Z����L0R��#m4����AO���mX�>�M��c\������w|G�)cX�C��O6d��{.h@�I�}�{3����ՒP.rˊ� .��;��w�&�S�fۜ���|�*�#�QP��稚�N��}g������ـ�$���gbÍ��0kH�jE��ē*�& �O�u7Lg��Gz�}���[�[��4\�(w�5V� U>��U�~5}�0��πG�g)?�p��V�}A��Dyz�sF-�+_��D�<|^:pDї%@����BX�{10���W۟��yh�.��&hr��=�0]F����%�;���fU��w��p�h���/�)pk�������T�+g�X� �MWW9����I�,Ř��q�:Z�6A��b]|��ށ�z*@Y%U������l����s�&�R�X�߮	����u������k��9n;�Y��>_�v���/�5�d��f���G���/p,Q�$V�N�ۘ���C���sJ�四�?@iP-�^��M�e9c1�����u`�z�G��|�*�"�.i_����1�R��2�vv݃mC�0x�����Y�e���f��Ϯ�	�����P���z�'~&�"�z!g����K�MW��z��ʭ�&V9���z�l�HX�X��䙛:Xy�Q�([�j�����l͸J� ^�t���P�.7�٬,8z�v$�r]�r±$~��`r ��q�l�%k���?�D� �{�d���'�\N�j�.?X�*)9��(�@E���.Qj���-���z�}��9�`�ܘ<�e8Q�;�ʭ~���8�V�%�l��Q�Ƈ�����'��2pTj����'#y�F���a�@�P*�bA�U�