��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jåا{�\�u�?߷�dn@6�zf��r������;�amb��ݺ����.?F8mA�h�׍ڶ7S�ګ��x�Z�,�G�0����pJ�#���PM?)zY�� W�8n��.�?R�AC��Ĝbgl�(q�Y�W��r��uV+����}'�$��T7%F��"o�*�8Q���ul�IV��뻃oC~rD�]}���e�2�����{9���:�X� iK"i�篃sv��X�^� `����-�O!2D�O�	},�����5E���$d%4�pe�'�-���{���VFr,�9(�멏"t�MFrk^�ߵ_-�Ow@d.v�<
���|(e�,ͱ1�zW����^�K�3�A�E0�H^n��(Y�@7��&ӷq~�k�׶D�����ڵ��XӰn��)�&�kQ^��E�7H�B�tE���
�挡�l:JR����%�& ��c�8_���i?�V��E�������#.ZT[�[�I�f�約����בi#؏qt"��b�������BFR~��Cp�I:��Ljhv��}��������\�p<�릤	�8�^y��N�W�t�����G�!裠=�|T���V�q��K�8�#��7��/�4=������`�Z�'�|�y���mE1���eOsB��,\fC�X�uKU�= "P���E�g���ˠ�U�H	�d6�����۬5�O�!Z$�qD�"
��@�c�����=e��ҵ�M>�"���%� ��<����c����/������X�^z���g�h���р���W2�kNI���y�TЕ��ĦS�4��A��3չF(�p�!t)2y� E�pM��M����z�&5ܞ��|�%��y	��f`e+���VL"]%L�{�h1q�:�ʬ�A&v��5�����Z7#���=��`�Ѱ���"�ˏ�ލz���;n��c2xw�"
xQ(lQ܋̋�:��n&����[!��彗�&;˿�9��$8�f��r��� i���x�_ȗR�\� c��I$�Ƿp��b	`���T˚/}~߬��<Kspt���DQ�ϻC*P>��$�4Gꥁ	��(��Ӛ��{�k�����<��,�Pw$J"������J(�0��5=l����ci�i[Ff�&'h�)�U�?���*�bN�륥�.������|
CK�ˆb�A�=�N�
�O�G$/��Q ��&�_���V/
�c��1�A���<����!f+�r�w�a?�st���������Z��;Xz�v�k5�[D&\��%�z�ECSeա�^ֲ�[�u����Zt�Τc��[�\rU�G*^���o��kV���`�t�2�U�bZw��xl��&���ɬ^���B�vX��yO�w����G� ��kܮ���;�ft�絓p����,|"�c��iGv䇲�ٸBt�[$Ŋ��<fu�)� �$���)�򎹉���LJR�r
��Us��H%{�BJ�3�Z4��i�o�/ �z���@dNl�kpT	�[0�U�Y�����SS}�"�s"P0zl�I�O�������B'� ���`~��8�pt�V���E��-#����v�c���m/���ϟ}3k��u4�(����}��g�����H'�GiO�р~��Q�6T�R#���t��`�o���.�t^7����#bm�`�H7�{��F������I�n4(����~m;!9X
Áym����o�5*�N��O�"�j8[��W���V��ʛԜ�7K��+(,;
'�LG��6����W!^#�"&B��fU�������]�D�ZS[!��KRZ� �hԏ/+�V�C�4�'|S���y:?Rw���:�&z*��2��>k��-��-��k��fU
H*j����lPg?�=�pM+di��=i��ykZ��	���:Q��!^μk�-�Ğ���T�v�w��$"BNr���/v=�S��ڕqZ����jy}���ťج!3��ca�z�rB���i����Ƅbl	�A��#�Og=}v���D]�\���Ԉ9���ȢD؜W���ᩦ"�%�oߡ�<��g�]`���/Y~�����.��ı�M�I͗�lv�ݽ4�����>p�D��:ܵG����&����SFEKeL�;g��h-8K��r�/S52���w(U:� C�I�k]?����wٮ����qe��mo��S	_�Y�S��`Ee(�N�O��3��?�݁��_?���܂ }N��׌�x�M'h���$��iY�m'_N�V�r:�yG��>vo��� Vc�}m�����c�&7&�x�I2�j�%�g<HL��v�~�Nۏ��#Uz��5,����c }&βS�W��"��,��X�T��]8'�-��.�۬��H��ʜwL�qnL�`����47��u����@MS��ϖ�����`l���S7MY�$m�y�W�:��q���Q�G���๲!�987����d_��ܻK
A�]!u�p�
���k��5���������~�����Ԑ�8��糷F��^0Y�֏�Ǻ�6���/��DQΦ���\�
,ˬs�t"��~ёB��	���y�;U�W���v5H�!_;
f1eU�I�^�%u�Ia��K�������q�x��xG�q�k��A]�b5�4��嬒+7-�EB,P�P�J#v�v��o�!���lw���JɊ["?�=^։�@���hL`�}
 K4F�FH\+�$�ЭW܃� c�~Y�5�\�x��9)����,
��~�q�B��,!Kh�j�N���ٱ����]�o��F_�U�b����D��ͬ�h�}DjzD�J���U0E!�<c5^��|�Ž����V��0�9+g�1bK�c�(�ϳmk��f���p�{������ņ������/���T1������Pz�:y�bxu�s�� �n�8�5��!��T�o�t&�Z�8G]��<�4�"G����Ԟ���d�N����u�z�؟q�|��n�W|Vp��!����D2��=̱<.������eg<f�D$@w�y7�����(WM��=n�� �OV�b��"��
<c�M�g�#6��?r&t�P�[�:�`^}��k�,
R�rY��OArr1j���e��ݛ���@7Le�S��+^+Mou}����m5�B�I8G�/i:CX�t6�z�n���5jWUZ�)��&x����Q	9�Jrpϡ���_<��Ѿ��0�O>��&u{=1�R$KEF]8��	X��Ab�"��d�4p��,��&�^E3ٟ��?����jN�<�(u���n��{�#T��f&z4Ť�6��sm�C���IL�;�gmL��A2g������b���$�+���y��{̃����Z��N�s^����c QG��K2����>�\�늼��0�p�t��;(�3��c����	�t��v��0��q�Cu)��q�e�ӏ�����nGCD�E#8p���F��BT�H���Ͳp����\/Kw:u?�c�|����ra�I �Ⰼ=��Ņj?��A|��t�P��VzG��9M	�wU"X���Ʒ!�K~3h.g����zt.a�z4��b���_�BsR���:zl<<��7 N�������N]�hD���=Č,��n=�N瓕s�4϶�����B~]j��s��>mc�DW5�����l��G�
*e�#���L�J��8��<����>��QiO��#�����)�ݢ��ȔO٪̾�%���*��sb��g>���5\z-�v�)n� x.G��&{��%���F��g:�ATC]��řR���i!��p��l���E� lQ�W �;׬�U�\����E/.�v�#�ϧ`��[�< 
�g����u�&�є�>��@����m��a�nD'��/�ʋxճNJ���~�X.PtItN��AH��jKc��\ܶm��\�	�.�G��Xn_�&C�����;� t�
ӳ��B��KE��(j�e��^Br�`�4����R�豯D8zF1֫��,�d��z��;=>7 !eI�,�,�����9�Y�bF���C.LC���BC��M�Ө����!�Fwjȯ��5���	`�ׁh�� WLs=f@�6��A����v�
��[;7""����<�~Z�C�[lj��EPy�2�&��<��&�?a}��g���6m�>� >KM;���^�6��$���8�8���F��Z�~�& ��:/��s��m�~�.���E�N�JzQV�fC��L�	�c�ȧ�:+�^F�x�j t�iA�<~2TYd�:��."������m�_LNb����!���Ɲz\j�
���bwQt/�zympjD)�h,�g�E�׎f�@
T��S!;�&�|lat�s	OD������������x�.�L��p��ϑ��J��������A���w�Ow�����[�� ���&��30�.�B����,�^��I(��\���|��G�{�>���:��o-ߓ��l�T�s\>ށ��w��螃˹f 9ӪN1U��"�h��~FV.SzT�ηDC���L�M0ȹ���uik(�6CU�X5,r�֬�#�1�ۀm���F�M:n=�h]l���ɜ*�90�D&=����Ed�׾���ąqz��m.s�������.F��*.bDJkж�������⡔BPL�q9)e_3W	(��.�<�e��>�v��.��eϰKl#��6~w��	�.�r��g���[4U�Y���ZT�.�n�����V�B+��o������~���t�G��\�{��\�ij`�v�s�a�����f�Է���uy-���P�(7ߙ�񷼴�%��?7�Q<[?0����+	�_Z"4\��)Ky��zQA�t�F-S�вQa���JO��|�W�%/�ާ��v��P�<i��$]�͔�RxJ��	+�l6nq>���wG�ɠ����>-Z:���O�bڮ|�|,��_�7H��L$Ή�㎐\m�m�.,�a���Z�F�P��u�F�*f�~u+���B�otH�x�u2��y��N(2j���5�N��I{�ű�0�n�m����ɧB
�n�Ȓ��� ���s�OL,5��i@֜�C�Ap�͖�JT�⴯`لi���Nu$��8eh��8�z�?��8�' C�9��z�X�`Su0c�v�6vq�`.���?l�M��$i��vc"�"���A����lZ@8.jo��()왼P,���$�I�[�/��q�$���
v�O͞�����!�������x(�'���Y,�3�aS�:p����3�|�n����;[��K���#�lZgx���>�k�*��2&�W�����Mk�Lu�:���_�{�~~������g2'U�u��4VҐ���Dѿ�������x)c�dk��ߏW��2�;\�\��x�4�2�r��4Ǉ�'�uS��EK�1��DǼƜ�悆p�i�8i�]�V�O=C[���{��B����W<�\�����h~Gݹ�ܺ��7�g�	&�$��;��DV��١�Oɵf/���^�e7ԗ~yk~�S/  �c!��'�4Nk�j��ݎ�`'+\�H>q��=�h,�e�e��P[<J�VZ��L���]U�d�+J��Y�w�A��,��.{�D��6�k��8����>�!��ǂ}I.��a����gs>�_����!��ʿ�D��R�scvsKM4�s aG�Q���ֻ��n�.��B�,�3<^���O��4���q)��	ݹ@btL���t8ܠ�Ǫ���\��[��r����-������m+���@�CD��#�G�CcG��ݶr��+���W��B��8��Ogޜs�Տ����B��%��
Hp�&�N����T~Jy�=�|�!4޾��:�#�D�Bu�e������<K� E�:�x���&j���@V7��ݺ���X����H�-y�  �^�p��Qr��u����`���#כvR�=΂�fp��� �����V
��95+Ζ2Kp�fЖ��@��]>h+�Ǹ"L�m(��S���݉m�G���{�3'7hX��O����^�Cj�^��}o�=��{�s{�OE��국Wњ�RU����ji֓�����K��&A5���j�(��������&���"fn�WdX�N��1T��oc���;�`��ٗ��YM��5��TJ��t��'{�X�ο�
��GL�v�ЁL$�V�oּ�[G��4�I��$;���D�<cˠR���dŷ9QЊ�`ˀR��OODr=xoH�(��<Y`�c⩲�]^{�ߊx׊牀����A��Gk������L�tM�+�S���	Ht��$�vJ�8���4����:��nF��4{>��6zU���)���Mֈ�&P^������޾������-h��G�D����������;����؈L�u�Gv�x�M��"�^@�d� a>�)`tw�n����u@ǛF@�����zƶ�~	�G�!"b�ӛx�����ܷ�������Ӧ����e�$i�O�I%�(-T���T�^��ۓ0�z(�������>�����^|A8��t����w;�埭~���|��\̔�1�X��`�0�ᛆa:H��El�(�;��B� �E:�k n�����N+�F'����B��"}+H�d��e�e�vE��w�6��WC�(t�"�Gsm�/��c��ľ��N�ώ
TС���X�)�٢�ɺmER@���BG���@R1���j�N!����T�U���H=[�tǆ�D�;������^�	��P�݃9rh̥7f�Ul"��F��~���,���4
� ���M�g� Ô��P���e
��*�����G�ˤ3v�}�_�g�4fwXs��M'�����Ǘ/�.X�#9x�0N�g������K�^	��w�Nv-�J���ހ�q)5Ϊ�.j������X���������?$��@%8[D'Q�ssJ�Æ���\�X�Of�I��]|`H��N(�֋/Ўi@�X,�9J�E��{�ng�E�f������́��C�1q�9��!�_����bh�e8<3� ��D~Q1ϥ$ �:1p�* )��oa$�8c�M%���j���`�.������B_;�Oix�V�
�%PS��[H�c˘u(b�J&*U��`�M/��Z^����ЮtO�NN&�4N-r�6�����R�ye���wt,"��[�G�"i
l^H7�МxEW!־��gyc��0B�D�	�L��vb�C�l)����"���$8(ۏ$Gs��6�#��5C}/��Ԓ�+i��}ȭ�k��C-����"�� z�~��_�ʑ-Kʝ�����!���Q�V�'���>���Z��&jo_�.�Vy�>�����	�\D���F �������u2�a� ����}i9�C^*�Z.�/|���X�r�{2|q�x&���@�S�u��s�*�;�/��Z8Lw6>ė�5��YU�7b=�Է�#=�ř�yO�aL%}J*��<���͸��n����k��ȑ�~\;=�~n���U�8�B�ޫX�N?�qBǇ}z���%�j���-C���U�H���kX�[�+�xXZ�e�n>��V�o���V�p����<'�1���cK2�9��e�Ȣ[��{�/`~�@B���]�⾀�E/d��O��UBy�4�Xx�]���r'��O��N��䵅!+�xE�D
�����8��B ���^�p�	�$nE�>�H�	�i�;��.����!v���r% p��-#����;t��䖒)��~*�W�����Iާt]�Њ���s�b�%ff��N~VP�u�e\>�5��:���qf�v��>��� �]m��Y��	�N�N�/�Ғܟ������Z:i�q��e�{��
e1Ҳ58DIu���w�ūb1</)"��楙���ǹ�4=���6eg8���0y�\�}���u��Z����)�'�""6
~��ƿ�ڻ��F�I����5����&0�HG*��=}R�@r�R�ﴖEy�'�p��MI��ӻ��02�+.^M��kJb����)r��Ct��T���U>�nK�������E�����khMW:>�o6A��XPߕ�i��
�/{�lTc��l �vs��\~�XѲ���+ 䔽'B^l���ʀ�CP�_i�7��0�ۓ9�j�U`��1[{��/��7%�z�{ST*I�	l�1����_�a.�U�*�bF!��oέ���ѥ�1�%�O��y���4�M������LYEQ<�-%d#��w�r�-U��'�P8�v�ҳqZSֿ^��J{K��Y@�bbQ/��/�ғItD��pG�0|Ј�t���K��f�� w�N'�=(�'�j�&�4�o��9�{�2 <��0�E1��Ш�<M"��5�QB�	�Ǩ����r�ɽ�`��@���ǿ�af`�L����&A��t��m�B�3�8׊0�0�Q���c�i���RdxY�ۉ:ls�a�;�貳���U�:��I�u��If/G�0�O�8�Ą&�
���z��ȩ������y`Y�M�q���g5n�$�|���V�����*/~��oXv���ܥgQ���Ҧw�P=����̀c}.B.D7�\6����lh�)��"~Ą�6Nպθ��1d���M��ő�~J�:���������K��uPxƊ� �FC�󴡞�ɸi(��Y �]�\�︗#�6�9��)T��^���4c�!��|�|:m{�y �=�ǻ�?��l�H9�1�B����������
��0U:��@m$�T��w�I�.%7�_�1q����B�ɜ�C��H�2�2M`�.n"_��.�r��F�����)���^69�2��`:CKV���*5Y�b^K�x�l�x��q���7TM���ʮ��lL[в�z���{0d�O���ɺ+���QG3��V��2X�0�c,��z���{�^-G�I؀�t��(.�� �ɿ���o����M�t���H+"x��S�P�v i�Eޥ��%@�$�����O#���� ��P���_+G��#Dv"0�A���\f��q�fT�g7#��D�e~Ԕn>D.ʠ�u����?M�Umi{�^��t�uO�a}c�w�&���S�CAL�>�o	��L�J�٬z��^&|�4��Wd�F�V�����q8`�i��*z�s`�lOz�q'�{Q�E@g�<���ZG7�1�>.6��`��R��-���s����C\�0��b�PK.�`xF�x�8H����6�[�!�%I��p����O[��Vx���U&�����g��d����k�r�/���7��&I�����<��3�G6s�jI�Z~C�r�C0Z�$��X��]�pJ[o]E�4Yp2�+c���N+cx&�YP�t*9��06b>�T, [\\�ѺR&�ױ,#N���!0�oi��,(O]+	a��췫�r�I���8[М4O|�\���(5wK��S!�{x��w"��	�s�K���Rtb@�A�Qd�9Ko��1ἱn�6~۱���E!+�6Ci�]�
����*`���-X��Z"�<W7�B��=ㅸ�*.��c�v`~p	�5�Y�]ɩ�I	ؕ>kp�k�1�%`�Rɚ6ǯS:���Ϳ�Y@}~�TGJV��Z�c���38�����+�r��T��lu����+X��m&��OX-�g�D���{3:ShʒEM�[A|9����/6�(�w�:�F8<=N�|�z��@�����h��fw��t.���As!�R�$�P����=d�
M�]WX��T��I�y��ɺy�{�(�\`~E$fB°����P>�EFᲫQ�>]���>����}�7��lr�_x
{?l�Ϧ54�i-Y��s}��{��W2V���s
�I�Q�@�)�Lt![��.�*��=ra�f;a�d��]��Z�8r�<Q[aUG^Òp����*7��O���Z�E�ާ]Ś6l�4^=>�[��߅SFy��q�dN���a�꙲�U����t <�E�2shΌ#�.��`��>��+��=�x�_϶�տKcy	���]M��9�;?I%c���
�j z^ L@����#�[��;V)��1����6�H2������	�$�%�>q�N��0�!>3cY�UzzF-��Aq���`O?7�������@��ީ(^0��!�	i�g�E����h�}Ӊ_�n�>�i\8�突X(86m)c�?��{��}t��˗4�����>�>��}s�W#���XI�y��Hu<p�KL�x�������i���l,�P./xY(�j@�P`~{M�x��0-�iaݯ	�bvK�AA�}�Gms��ֵ��$�7��^�m�����T ���R�)��C5�$o�i�9�@�B�X��2�2 va�Ńz��(�::�͵�"����$zG�5@9{���+;�l\6NZ�?��^���(m�|P��(�joL����hfU��ޭ�r{�[�>�}���"[`cXҿg��̧��K���>8�ì���g3��\dj<�6���W�p����Th�E�[�F��P\���{�������x1��T�XZ���̘G���r�����:��{�&�L�P�g�����5t��Ӆ�p��CzN���u�i��0NN}�s!yb�Iى��E���grV�́��:��	��f{�֒FQ�,���:�gX�2�c���8jMEdi�:�*/#-g�W��M��c�h1=u�V��(a�vi�C�*��v��T���v9~D�W�(�N_ڊ�鲘�a:��.���U�M��t����Yln��Y�׹_9�U��a� ��߇���`��{pD/TQ�*DެnN�.&z!�@��Lg��{��[y�k�݇U��`V������������f��5�x���IW�ύ�UK��eW%�+�{U-�a.5��fXM�6X��;(O��,FC(4mfv^��\R��u�㊣�O���)`�p��kzٮ�G�,NT����M9������J~�����k\�UR��Q춘�ܔ�X7q	sJ�s�O�w��;��e
������y6��t��$�&�|+]B���Ê�����"�mQ�m�T��bҌ��Z,��`�o3��ׂ|�V+L%��00�"o��$�`W��=�N�&��n-8�ުѸ�T�<�T�:��qklR_r��}sa�]R�egf؈�17 Q��8=�S^ѣ��H`�2cNyd5	Ud�'�ـG�����~�U*���Y����)���y�2s4����\����ν�XE��\���]�:�������烦~�����~'�:i��SAν�l���,���#��������c���fĞ�&y����Q� 9g�<���um{MtN�"X��?��R�S��J>-�i�w��3�>�0�:f�O�?kF�)�	��q`Z��>�]M�����'��{��gāH�N6���=-Bٌ���秅�D�݊��"?t�������>�:�;	�1?�3�i!�o����G3r�%��۔�#�:9lT��moͭۘ����ƻ�«�������ۇǈ_mx|���~y)?&��M�c����Ek6��
���'��F�Z�׆�k&Iv��߭NQ8Gٱ����0T��b!���I�eڱ϶�A� �.B�(ȳz�+�����m�GIS Ä�R ��o��c�hq��;m�٫�a�r��/w%��ϕ��bB�$V�=
D�n'^����Q���6�l��ZL�A������6�F)��&W�pN�Xޤ�P�/P�����{7)4*��O�`,Th5�*���X��q"t��:�`� ��,R��%���i�[�+����s���6�K���U�Ȝ�)�[&o�ʹڌQg�6x'�. uSOy�L!��޵PbL�����i�W�n�hpl�<x�����|��X0���s��I������_la���Q�E�(Y@S{��w���9�Z�_]�L�-"��58A��$�����a*���P���mѺ�61s�����8'�>�����r�e���ꁪ�q�����QT��l���aQ�U"`�N���uQ*H�d�Nb�������5�B��/�����y5�0?_i}#�c�y�
{�0�3��B�����&�t�!�ܝ9�z;������yR����L���=�-�����FVoK��M���V��|�H�v���h8p���ptF|�n��9�\Sx�� �rӚ;Eq"Af�L��;Xa�RP�c��o����FJ��np�G����[v2��As�@*�I�Bſ=�+���ˢDg,	S�/Pl�닙�u T���4�Y�L��bt�g�Li
kJ�=`J-�7;�|?t��O�_t��d���`���6ڈ��qs�`��QV�\"��:E�;6��듯�Ny;�N�����l��z���V�A{_Uݎ}-���h�Ö�M��l��=|e�H61%�)ۨa�脥� �`Ç&�H�=+��8�<T7���#1iJ`��v��{;���8o&���"�2��:V&�L�1-!�f+�c`�V:m�JVs�4!��?�˪���Ԟ�҅�@��s��pw�[L�Sh��F��g����5�Qt���q���S����L��"���*!	�I�4�0o��9c�	 �-�?����4E+�H���Q7PB�������1��)���:�$Ph�V�}Rw(z�nՍ��Y)eg���Es�ň��<�) �1|QIX'��-B��R'wvS��(�1�z�A�_p�/1�50�O��{�L��\�j��8ݯ�e5w�޽?쒂@b�x�_��V�$ոX6Jp�4Ԍ�SeT�37r����[!�<�\�jt}G"��Kj;H^֝Ok�O��ӕ���/g�|��?j�C��~��e�g��M��۾�L�c����^Bg;���*D��U�1��C��5
��q3���R�zkFo
H��d�쪛j,)f�8O׷st��s��T��_�;r�$�7�p0oA����ӳ���H�$6�U�G��~k�1���v����t��,E�>���)���_��x�|H�>畬�(s� ��?��f,+���p�a^%u/��m�t��M��c��ۗƷ�vg4POJ��0U�y:�i����`���A&���y��#L�o�?�F����=r��d����01�	]�7���RGx��5�ٗ���N�6D�n��Y� ��9V*���5C"qN��"�n'�J��Yߙ�b�t�������ۜ����C�(+�ʳ����#tg�}t��U���l�����^�w� Z�4K��G.By��y1?�wǲ��!r��B��G6eբu�����(�IK�գtP���M�C�󬕻�ђC�[��<f��C<ǹ@{'1y����lέx��C��O�@U^sXH��>r?z��[��ҙQ�0�i�^�3�H��S�����~(kT&-��#�2��$���߲�xz�Wi æd,�3�h�E_�����RY�g���#�`�b�۪/�'�ۆ|`Y�j>Fe5+�>I�ť|�������#��w�l�t�"L���M�cQO�X���CH�mSB[-���(^�Ѡ·�Q������G�U�g�,oC��� S���2��������"If����|�Ɍ<%ޙ��h����l�I}�uc�yQ���!�2�J��:��06k�5~�P����o:p��P����>�M�d�{Ahil�`�2g��R���[*4��B�F���U�C9��T�.�yy��B���ߎZDo[�`��t&
�:�`
7EK�9�_<��>f��9��G�Īa���H.��DF�Ym��[������5�]b=8=]D�����嬣�[�+� I?��h��R�^��j��}uޑɧǇ��Bܸ6>��p�R��#���n�BKo�<)���t���MO�>�ۘ�@�pLv
��?^^[6+m<�}�q�j���/�	v��L�v}�v�L���$gmPǱ$S8p>�(@^UR3���Yq7u�%-��&�\�1[�ʹ�n��Gs�|�M��C"�L�&����f����QAyB��h��_Ԣ�q�_{?����KaZ3�pb�{jm��PP���Ή���{�9�kJ���J�%��k�1<��/7n�S-9}�\��1������Ās�E�F"��ь������OKbƖ�?�<j��	�k(��1a1y:�4F�{qn$-�R��Q�k���*d�4'�+~������|-��P!Cn�r/�������������'��}ԡ��[V���y�NMh�5�Ѯ���rDu�v��ы��W��u.0� �}ΝxTA�؛�]C
�)�G���n��%SG��_�n9�ۉ>V�:v����$qj��[������n����� �><����7�Dm����/�[�6�[�V����F�3��6$������!�~�R�6����p�;m�d؍�<ء��Y�d���T̕T�������\hf�����&k�6:��b�p'�${o~5��϶�����W!$��Z�Hc��'�q�&�xUu��3w#2�W��'`�J*�G@�h�q}i�r���}��(a���p��}ٺ���f����w����Cj�f�P��M�y�8lC�H��,���d�h��g$��Jh3Y�;`U}�%����*g���$f�Y�
S�۝5^��_L��΄I�u����������Kˮ���"�Y'����6�۵Μ�Y
�j���n�Hݿ���	��)/�B�Q�wR?�G�����,���laM Ծ�:���L��W?f�:^K�E�:��fdʢ��jy<�~ڃ(�/0�{P�>)�p���#�zy'�"*��l�4iq��%�]�:�ĥx��WnW� /0"�>�U�B�2@?��N>b���������F�Ƥ��b�\���Ѥz��h*�6��}���b��6���ciP��M��{�h(����0A8��i��j�9���D�fK� �d�9u�6|ױD"��2�Q�� ߯<��X�8z�*?42��'�;Q'B���s��Y&��� u���#>�o;A=��W�J�r��f?)��E�J�^�M���mZaA�f������%~ �|��OG:,ׁ�����V38ʾN���!=eJ��u`D����t�sa��b�}}��;�n�*N�ք¥����A\��a��
4�o�R G�5PH�p'�m��ZC:cRW��<v�Gѷ�cG��^��u~ ��%�ߦi���w�x��A���DL4�iH����w0Bm��c4�Ÿ��Z8��ۼ��ʖ�3�M�?�G�e3�����I����x���op�?�
K��)��� ���V������'ƯT;�ka��P�K�U=i��S�?P,��[�Ӆ|���˕졨�\߂J�'rg���RY�ҩǱ:D�yO<$�ԕ3������U�4�.�5b�K���N�{:�w���Y8�ٛ�7i��v
G�*�=J2b���2�C�݄���)��j4����=n�C���$�j��gH4dj�,��^m�%�eG$){ش:(��-&W���e/V���=�8K�h��.��r�9��̳G>drJ�/�˩�sq�&���b=->���� NP��YO���RJ�Et.�y-�?�O�p��00�}�O��[X��jyp�������˵�%�K�9�P���׬M���Ǉ������?�˩x+w�ٿs��%�8�	��&^0n��YU�504���\��ب���������zp�%��}6.}��-@FJ����/�U��.��������Cj��b���f��"�)���o��@1�6���a�����ߜQ�]�Z�΂q�y.�ـ�COL Q��ST��.���9�W����Xd,}��^��E�����-鴥98'������P���F(�^�kC�	O�|O$-ӭ��`z�6M�6]��#om���}p1��n�$� ��g/4hѶ�v���x�}��NY-G<Cl�[�3�^œ���auq{�쬷<�%0T�K�`���W�N~�^��� �Mӻ�u�<Y�q)�B|���a�@�Q�ܲ	��p4�W ��=yg��,�D�������vT�5�F�m��`�?n���"Ɔΐ�{�u��O��8��6�E#ּ��'b��s�6p2C$���Mڬ&9��V�����#�1Ø�L�CR��P�@K����k�v3u�15��b�a`�V�c�#1r���������9�S�r�m+*���o@���׭yí�>�Sd%Z��Y���M���HrWx�X	kZ��RH�Z�h�M�%�z���T���g�TW�(��,���r�F�פ^s�,�[U;��RG�DSM{��߅ � ���&�)DήIM{o�A�X����o��s�7�a!��v�̧���Ӡ����;��FT���j�`�K��w�P*:��JlD�'��l�L0�
�r�a���X�֩��dJ��U�W7�z�)�2'��6C�LzL��ޅ��`��Ag��-6��1Uͦ{�M�ϩXU����³:Q新���'�eF�R�������6B;H�OuF��7o~��ܴX�M5���,��`s����d����j��df�tv�������[���c�x��� �t9e�q��1�.������ܚOO�.���ٙ��~[����c��\��J~���m&�v[XW|{Iw�#"��8eZX��D�z���#4��Z�&�L�"�Ѽ�p���?:�s��u&��>{��� ���Od�KIuN+�ӇT'�^�kFV4�p��)(C�}��E�_6� ��g���$_��5��&8�:d*@�2!�F^�@��ƫ�a��+vc:��`����N�5;,U4}�#��s29�DE|7���W�ny�绯��P��*�@CގY��H0����K}t"���� 1Y<��϶�A��4=��D�ׂ\rژ�R4�b,��>�4�������r�d�o) �=δ�Y	��@9�	�=r($��[��
���=u�1M��� v&�9��!��(�z�-��C����&eD3HJygi��,��@�@;����0~*�k���<��z%�v�	�":�e���_����8
V����!1�f�dǊK����X���W��y[�$f`[7��H�U�'iB�1�KД�*�*K36��/�5����$&iY�/1�l��R�P�I�붿��fB�#/b���@����^M�_�	����?��!���>)A�K���ϩ��d��&�ʁ�}�x����\P��ۄj�I̘b�R�����t��Q]�TjV�"�Jp���==��u:Mc��l�T��$"�"��R9o��Y��������j��bm��!��G��Tj8����47(�P)�~{@i�F��t��:5�Tz�(���"�ѬP�2��W۫���P�[���.����D��șܛ�F�`9�rlۈ�G�(������a��Yy��:ltݔ�sQ���S_���Au:V�~����闌�5����?e=��6�'�|3��������`\�z:G�"~�*LC�1c�
�>���¤��'j �B�%z��?j�T�:�`	�%�j�d���N���.	6�t�4�Q�ou=�͖�CS��N�?-s���H*�����2�N��O/�F���oU�Z�"�^?k��p��-S_G�A��W�E�����*�bA��4O4\��"���-�g�/*A![	^N��*���Y|rO�� �|�Ty4�:��@Z?H�q�72��4�NCo�:r}��{�N(
�l� �z,7�}O�� ����tX�>!��\���f0��=�U�[:�}//'�s���עhJK�;�E]ڡ~e�<_�2�/k���%4L\�'�B���pl^ц�$9�#f
!#�X��Q��e�[r�D��&���)��3�&����Z7�5�l�^!�uE�pq)�/�$AD˾c�ΌlFه���;M�Vq�wS(�j)��ق��I�Ô��s����Rnr�'����\����Ӎ��%�^:H�ԁ����Y�P��Ya� �'�(���m?�j�H���4����G���������(�"�[�1;+T�E+��c��` �X�u��A��./��z�Y���\)�/�Wr���s�����%��x�e+Y�;��a0XӫX�d�ǔ�3��1�`A�B�~f.i L9l�-�I��G�Fk�u/f��cҒ��ڌ�XƺqZ�6ԈX��8r!G�c#FLÝFЋ�Y���<�[]��L�sa���֭ܙmv\jx#���Dq������zK��0�>�V{`7V��!���~>Z���ql��/AĮ���P�,d�Q�'�y�ڿ4�N��՗��ɦt�XTa�أ�.��W�DiX�Ff��$O�H�C�NIz�ndϓd��R�I~F'{p\�[D���G75A�_��|�{�Vҵ������0�c��>�p5 �xP�ځ���H~k�G�ܕ ��B/�:�`��@�E, |~�Eo�[��Owlٕ�ti��2�A1&��oڠ��_qh�z��T�K֏b�α��G
ԝ�����kRG���5գ��߫��R�7>��B��l���bM[��#�|��;,엔����-<��s�G�΁`%�I��5v�� 1^r�R=� ��0��d��.�[���p��K�[�Q��*曻�����lg	����C�׀�iߢsV|:�� h�a��)��zi`�ٗ��>6��{�������ن=9Yn�P�=�S!�~%j�T#S�4lɐ�i�mɓ�
��|IfGJ���M���c��h�%h)Pg��]m��ǒ�W���l���{�K!�u2����|����s7�FVV�W	'�v�&vaȠ�&��v�I�4�@�N7��ʶc���#�&�~v�-��n��u9���T�ȸ��0�mi���7����+���{{h5���������+���e)��\��[���MG�L��]�9��-gW�`f���}��0��}��M	LL��q�H�R�e%6U3��*p⭔ո�v����eV5C>S�t�i��q-���X�F�̓e㍹����7U��<�ց,�k�ȟ�:�Y�B��i�!�+=|�-�R��ʻ>�5�@���pL�@wF�n1}r�n��4��b\��U9�Ꟛ׊�����0	�˯�YƖ<?�s����-�Ƅ�f����P>�'����v�0��IN%�H_.Dʁ��OSpYȁx��e�.�q��HT$Q�NyjD6����I{<w����{BAޖ��p������[���N��vt����#�Pbd�ҵ��lc[�
�<�*��Jo�d���J4n^M[�@gOY�#{	OLF�?���`��,���ە�N����j�P8��TNӒ�����'b���"G�n�w�FI��� >�=�p��)����nn�b��;�k<5kt��w�S���e(�ڧ�����}v�>Ϫ��̬�h���/ŋ�--��i���Gɸ�P��y2g��e�y���{�fN��xx���B=/N�g�+6��L����;3��E2i����w���ky�ؼ�jJ,8���M�p�'� �$����d�_{��������sA^�A$m����<CQcO�1����+�I)%Zg � ~Yw�/��az���aRpc��r���Ґ��C��r�$�d>V�5���|�N�69�?/����DlR��;�
�HUC�& ��$/pj�H��R���'�x��G���c��P-Pp��$��8w��h"6�&%�#C�����̝F/���uo��{�X�5S���Ceg��2!ε��H���2��X���q���71�Ʒ�ې�)v���&|bSJ���	��9CfBO��1n1��n�Y��ɥQu7)��l�e�p>���O�w�{vt$4p���(usXZxw�5����}������=W˞�H�&fe�uh'j���r�a��4����H\���/����9��4Q�Q���N;�h6HRf{;��.{�Ki�����'8�ԎM�M�� ���������1���}�W��6�	)�+�����N�-~�뱨�;����F�^��F���\��5É���(u���[��Y*bg,%��8d����?����h��*˔G[�,e-.��s�3�Թ�<�;s��bK�w'�VqwJ�*������O�Ak]�<�{n:J�S�_/V��H�a<�A"��}lY��'����Eʽ^f\V��d�O�~�đ�m�EŠx�'��� ���[���h�l�E�B�a����)�~H�:A�A09N;^T7�^�M�������� �h�J�@����8T"쌛��M�,Z��/w� ���)ʜ�&���"	|B��r�5��4B*���tt���A�����߿��TNA�2���9��NvΈ!-�M��(�@q�R�t�%��{t�y����q� Y�b"����0�R���f�w�%+�w��$��֠m��*K�QxR�U�Hj1 쨇M��ϲf���N�8�H�j���bH)����0kҳ-<M9t�EN�7�1&����'���U�xK>ܾ{��'������&�1���-���|����}����Q��Dɻ��T*೎ʜ�t�0������.��t�ο�^E�{�$��~�[�����'<�G���%����<"��
�bB�䜠��X�T{���ǹO9�ڭЬ��r�1�7�a����	˘PP��1�;��]FI�5e��A��|L��� ��CR�������!�eI>�و�[��<��W_2��x�c,��ƹ�^�$��)���Ǖ1K�\�����8��%�Bx���+��?''o�b���CM���sYfU�P�dP��:\�=�x�ѳy�~"�<�&1VF�K>�}�H���0��ZA�|�3&p:�lN�Z�<)�>Vk�.�Ak���ԙo���m�WT��Ļgu�َ?��Ŭ��L"b��aޙV(@kp��4�BoM̕��̱Ř���rU����ϡk���#�S^?RG����6/�R�"ݯ<��ϼ'�b�4�Q�_��E����Hc�J�X�xS3����%���i�<)05N�^�.m|��� {M�`�|��l�R	@s���y���i �5�V_�4u�Y��|wo�͚�'f��R硹Di��4����'"L�!'f2�]�_J�̎g�^�f���r,��k���%Jd�V����V���֤�E5��y��Ξnz�?������~��*��X[� �1�R})���O�[HӔh��TK�c��'?	���J�U���ϖk��P��{���֎cSA��P��M{�~�bV���*�+�?VK�Ҳo/��Y�6���z��ݤ&+��г�>_�|�e�8���p�[O��L�԰��A�N�.�FЃr~���(��^C�bO���D3���p�޸�}�����"cݎ�G�v�M���6�bz�A����sI�7��B�Lm�@ʆt�|�y�� �9�����-�,���Z��N�0�"KQ��,4Ў�Q!��=�Tte�[�L '�o���Q]�&��&H��t|�3���{<���S'���oGkxa��h�(��C,v�`!��e�?m]sE��O��H�vCC�z��%��L)��A�G4RZe�"ՠ?����u��`��㯂N�a��s!Ύ1���U�f�J3g�q��@�p3ߍ��@n�6�^L���Ds��˸"b�`V��0Uh��t�+�[�G��dP���/����_Hi֙���?��Q{&�ڹ��{��Z�À�[���_��t�v:��\݇��2���Lݗc��YM!7��C�e8�;�*3��_c�#p;���d��3�(A>�e�K���H �:Wb���Vg�CUX�!��.�F����9^�=+A��$J�8��Q�N1"C�d��r�:E�gRU��������L|FC���OX=$�n�T�����Eq���&���]��	K"6Da���;�����8���q�~�b�%��6����c�t8�}f�&�OX�-�ҀbC�+J~�i�Pܟv�27�K���B� jA<����*�&���fT� uY>�{ٸ7	���9�-�I�-�^W`��g��/���z�p��V0$Pl
a(������`ǚDdy]���;�C�%?P�����|�j�&4�_wAؿn��갾��֏��h�QU��š8��ew�NW����e%�˟C/�-��I~�ZH���c��a���ㆬy�D�G(�7��a�5�H/���H��62,͓��g�_:޴Ij�>��uQ�Q ���ߊr������Ѵ	1_�#+��࣓|>N#��Pd���V4x��R4m,�=���Ȉy��-8s�"²tT0�mj�|KWF= -)��1:�`6�� [� Պ�N���@N n���'s]E���1G������Mؾ��c�9�f�'�7�Ư��������A
��;VI҈�%����1>(�0\�k�c@�H�Vkq����� fw���4���&Q���%Q���fy�	�x�G�����d�^Z/�OƑ]���(�vni/p��HAҚ oZ�v�/t����(�5�>_�,�GX�b�/�5ٿ��`��M�TBV6v�L�����@E��M=2�:&v�����F�7&�Ϻ��4;��h�9������w1�@�)'��Ee�c*�Fv�p�J��r�������T2��PiX!I�樤�D�J��zQ8��7�a)7K�{R�=��&>�WA��8����9��Fk��^R@��I���aCd��M���V���eF7OTJm�@����g�F��	��l`���(d��l�P�]�'�}�$����[,bz���S��u���D��][ܞ�66������VpWu��ļr(*��`�S���<�b#[�<n��)(|f��>��� a?���q�-^ȱg�J_"�����Ϣh �[&I��i�:
��d�V���GӇJjF7�VR.l�_'�xK��(Vq��բ�6d��@���I�);��/�V��g(��t��s���7qX�	�_٠�A�_PT[��<c��h�9 ����T�ڵ5[�#E�2�u���ϐť˞0��ڵ41�l`G���I�0$������M���p/�9�Ө��9�뜵�
�G�s�m7u|MK�D��T�T����n<�
�C��D���l�z�ƪ��\�yS'��ZyPd1�Ih*~�B�؟��ѝ���"�@x&zt<-fT��.~��8���~S�J5'd�n�|�IK�G�?Z�V�V�饵=m[�A	�7
FVi,�v9��M�B+>����CH�8<r�J_��us��)Z � ���U[���@ux9��Y3�Lx�(�����WKU��<b�qL�Uzi�9q���p��^��ף9�*��cU����{�Dd��ؖd���~�d��}ހ��f�ƕ���r������*L�14�r����܅�ɰA]�OþX
b��h!w�-�K ��w��4��Қ�Ha��Q:4/�
�����N�J�����	�H�e�#��
�i���}��n/��q�Y1�?�"�N�B]ة�,��W^u^;;>��ٷ�����	p��w�����4�USΛ��܁$%�%1D_�hO�{�e6�	��$�[�K@�

1wp/�&i
�n�7,����-�C��_����O��Z��0sU	�ޫP'%ĵ/�Bi��Z������и�ބ����̰C,�k<A'����^��q&�aX��w�/x�Lh�w�����o���j�#L�0E��7�8<[D���N�݂�q�ʏc}囻Vs#swE�2�C!�{�C���ӬM�[5e�G�PC��������$y�S]B����m��4i2 @F&��6��\̈́sڧ8+��J�A^�6�!ޅ���+����x�v��w���a�#Y˄���Lp�E���8؄���v߾ڂ�ɱ��(9��@ǌ����xn����h_�Cy=���oʀr��Sr5�K�MK�ʊ[��v��u<�+�=�����Yp���MX*�l'FW����(dT��0�`��ϥ�wYv�Zj��c��)C���Ns�v���М�+��yj�/�R/�J"��6��l:xct��5��St�<"��
@8��-����T���-C]��Q�C�yds������؛x1�\󌷄�I�hP�va]'�H
���Ｓ�<Fa�#PQ����*�Ag� ������w��`��R�%zG�,�X�\C���N�_���9�������#�w�,�-X�	MY��^ �l�����\����x��㴃i��J�L��8�w!�6*�	g~iW�\ ��'��9!���%�Z�� ���(�
�nM0�:F��MvG�#�ZS!7��.�(1��C��fj;M���_�XP���I�M �I�/�G.gezM�$^;)�VA�YJ�m�R��h �	yJ���J���xltY������kt���g��5��#E��5~^�Z���Q�+)!&/�\��czUh.��L�Df�1��:��`ٮ�^�}��`v#OQ�/�c�p��#���7	Խ�yn߭�<�� �K���'��m������iԀ� �V>��/�m�R�ΌM�-k�4��1�bZw�J����S��u=��*'��e���]��>q(� ����D��E�A*%N�I"���]f|����~��	Z��4)��"�OX�Ļ¿��A�ON��}���Y}��@2�_�^��i9>-�=gv��~K<�/a�2M9�ā�/��Dt0A֛���@0[!��f�t߽%V!|JƩ\�l�[X��2��~L.̈%nv/�г%���*~7�r��	����͠~��b(�M8�xw�i�6��\a��r젪sp	�`�ώs�.rUk:��z5bV9'BS������~da�c>�n��7�f2��ODg^���4��2��R�L	�@����R��K��벀u�<�r����֝�RW�O! �%���o�Ƶ�i�U;����|F�C�	�<Q�����=���n���x�{[~���3���ײ�F�>�^��r��8E��Z�z��A��/���C�����'m�x�,:�&�n,�u>�3h���hZ��1R�ȕl��Մ����z=���)Y�ȋ�mYu���{$�=��µ���c�7]}0Ś(A��`�|'�o���-c�Y���.�|����wwf2w ���(Z�^կ�hH{B�:Dr=�[�dku�i">�{��H�%Cz����QMpL�j3
���E�wq�i] 4f}oئT���E��G.^�2��V���9N_�B��v|r;��<|���NE੸�˨�^�xA9�B�a'�?��|�����U��b=]TR�{��;������Or�U<3����Y?���4/5$�ؖS=����_�!ѳ�e&����p���?7S��#<�~YrjS��>��NYK��i�k������{&��G#ԃ!����o:$���/zt��H��6��|;�Y1&��9'�X�E�;|�t=���轲0X��AڏG�����&!�凨���j?@la�g+��v54�ᰒ���[���#x�W�Q���?�d�ʛ�oi�D��
����̇G��KP��{�r��q�db='��ϋϒ�����N�2 ��ʡo[�Ø
��bN+�f^i�^�V��% �.�7.�ktQ ��k܇.�OM�K�B�Y��?BO���f���v���P�ۧ�h!�q�i2�w8��)��������Ũ�w����"��c���4��C�Y��H/�KX��o�񆟩�dc[�bI�S(��w�.z>��ڏqo�WQ�H��?���?J�t���(��o��zoj���1��V�3��3H����7��}�dj����bP�dyL����4�P4�p�7����g��͒�^^1���$۞��������ҫ�J3� #��3�s0��>7���Ѽ����|��\�^��Y�@&]��A�����&2s簰��cp�l	�$�L��؁���"L�f�c�=�WŻ[>Xe;���j�`4I��瞮���0ה����N���T� B���g�x��v�?Z�&���.ָ!A�vc���N�� �Z
��F��D7�%)j#�������'�c~A�v$<��,���aCF3�VPL>D��(@`��.V��c���3Z��e��S�Z%#��}A�L�<+e��j,sx���k��kO��h�#˥4C�{Lo���V�~MN�uW�r����a�!I��E5�	�Rd� uc�w\¢�U;ʌ*��.�w���b��n A��Ki����M�w W)	���d�Y#V����H������yAf`Ѧ�lE�$z/-�qP�#�7� 
��	�B���ʧ�^�����o�Ξ۷?�z�\ '��4h��{J��o~E��Iྉ�0P�M�͟�̭�|�b����	�0�$���8/F�M�N9X?}q#�ԩ�t1��z����3L�E����{��?o�������#�����M!�-�a3�mŒH&ڒ*�V��$�zrMBd�7]�����* ��$�әj��P<m��Sh�Jn��������a��?o��}��0�>���?�1	?l[�B���2���hh��_�{�g�n�Qҁ�}Q�;���3c��T�'����%��5E�- ���}\�|w�4i����m����f�b͔��O��4�>�j[+3�T.{�켤���F�gh+��Er�[�s��v/�3c�d��k<���p�F�w��N�!Ay�Xh�3��q��o��e:���L�M�Q�`���C���S��qd�ۉ
f��;�}JIlhy�ѿ���q�Ҟ@�+�:
��E/���*����N�E�xo�f��K�-Mً�@ǒ
�z��C��*cc��e��]��|�찹	�W��N���U�,��Eyj+�XE���h<^��80l��F�ܰ��a!�4u��n���a�b9<��BBj7�7q�x$:4c�����M�����?����Ŋ�ex�Z[�RY&�[�@�ZD��5�OD���D�}���1D�hL[�(�.	�V���n]���4~(��[��XkM�ͳ�f�N�%������2��0��3?J<7��@�8�����qދS>�@��K'5��[q|�+�Y � ߴy��Rώ���@"��6�wݕg"�o��c��ٖ����Fjfi`ܦ7����$6�A��E�Z00ӵ���\S��6�9JK��YJ�4�#����D+��C��I���Zh���my�HLe�#^$�\�z����ʼ띋��6˜�|ۧ�� 3*���"�)��Λ�OTEG6���'!��8u�f��6�V�_\��]����0Rj<)LeDܽk:қ)��4z�m���W���X-��"%�4��L����D+�q�B� ���?�)ee����`�����t�r� �镥��z���Dil9a���4"���b(Aa[E�'��6��7g$��R�����x�E��&}Ƃ�{�����dSe���+�����'��8h]: �5K]X��NbA���ʒ�*��v��i�;���	��11�l����3���n�bYb�.�h�g���y����X	1�tܹ1��,���o�9������n��'�*�q�X��D�~T*`#6�7���L腿iLU�2,�{��E�?��L����a�1��@�Z�ݲ���Q3N�jkۺ��tFC�� �PBr�HHVL/j��!°�y���"K��Sb��qW���1 ��jz}#��4��8*�J��0�t�Ȅ�����X�T/0g.·k��\�t�R _�LF�9vdp�M�w}<��ץ�fЦ��f��Aų�	GyF>;{�R^���]�{��(9���ᡆeǱ�����ኪ�#�.��=0��� %nb���۸3���v{���/J]8��n�A�/>��V'�^�EdM�-m��) ���D%���S�߼�)�.�,��n�����Qï�g������f�#w�F7�=�5���w2�?�5�ϥ���i���4�~�o94�>0�k	.�\�M�@c��\(D��-�53v+�oy-.��������d��!(�B~�LlS u���ҙn��l��u�x����~:~�`����2Ԗ��Ms�f̸�$��ޠ
}���6���Tu"Y`e�/�E�yG�✓����[�V�3�b�|�dz�^�I�i����]��*�:�ʓ�SLG�C�5�2�lY�� ��:�.;�N΅��凵��H�q�ε�2�%�����W/?7����9��{�u2�<!A����"�2��g �LF�~�ПH��BפDw>���AH��M�2�{�\Gi��1�-w�����K����p+���%�p1
�	]�;��d�e��	i'FM��重j�	e`Q��"vG��l��8s�g�4�'p�u�z)�����n?�x�	���M�3���L���v��E���34i2��D@����`���ǘq�Q�����YmMY���	�IB�0�����\���>��<� ��.cl�6�si��%y__�u�B���|i���@ﱭx]��� ��������� �W}{O�LK_vT�wʵOnR��L~=~@�lU�C���/B��2����+�f4� D�5"Z�SD�7�������48��Ah��Uc�wxs'R�����ӡi�*u��{��=w�ĳk�F:9���[�ɜ���A��2{K�QU�������+I9�{��\^uZ<�h/n6ɭ��� M���7�ib�#�^JU"�%�"�ࠫ�]�x��k� !�D�a�4��;n����?Nq��z�\g�dh}�8.5=���,��L�ym~*Fdpo�������O��[�bN�4I����h�ۤ���d����"�bM {�\L�F#�&�'�N�4EK�_8��G>�zT��u��?�����h���SkO�A��K�:��5��n+�x�Ð��++��jVшx������~���{�"	��r>����}u䜙�T�lL��$ ��ȥ������(��b5��]��d[ �@YqQ7�V������q#�8fS��px {lp����g>(��^ |\w���"i�j��kփ}Y��������D�R�G�hWQ,�U�P6��J��֒f6;Z���r�� �re�t�����O�<��ü!��}�2,�&��%hNrF*:؆ F���^x�k��h=���eG�Q!�[Ů��� ~D�a��:�����P6��C6uD��
0�����s�`�͹C�B�<�-�n�B����j`M ����]<��;�]#�#q���M��`��)W��Z2������i��&i(d���H`y"�Aq)�Rc�UY9���Gt�9�_k/Dud���?��^��*��'w�!Z���@ŭ͐��X:�"��d:��E��<^����#S�;���P:hÎ����+>j&��L�6��ID��j�^�Nа';=�b��g�sf�,�4J�����}
��_G�t$�>���T��^�ˎ�<)���+��T�th}>1���)�s������	��Iz�Lu��j��<���9!�B��TKu��Y��{bנ����� aq����Prx�P�~��'L�W³��(|����5�`,���f�dSY�e��Ԇ�B <{曟���|H�S��%V���П5�6.��Ζز�n�z��~B~ӷ@wW����]���❎NOL@xtΙ9�*U���v ��;�ʁT�"���s�S�o`�����S)�q�S0w��$�����m�`Ѧd�xYq����&4��h�J�qΟ��`^f�����~棋9��FV�2|�>�Ӝkb>,Ʋ`|�?�uQ@��w�o;��J#��No�����C�pԽ�zӄ u&*|.���o��ّ4�� ���N�_�S&��h^1������E�q*�\W�-|J��@�b�u��p�P�Ћ��:v��sk>5� �������2�:s���>���}��{��tCi��|�i�'�,G�T�:0���`i�µ�����`�b�g�Ėy+,x�e�dK�<�70)yg�͵�l���9�r���@} ?r�1�Q�G�_�f��	��������L��?�a���I�H����Fx��-���~Ht�	u����ލRV�S\���nj�|l�Ar� �gs^$uo3�&��.r��A8��߂����Q��S�Z�*�1Z�`N�}I���n/�����1�t���u�����<��4���>�GZv7%a��HFUq��♕�!���l��҂s�o�_n/}��D��χ�F�x�b�B�hڬ}����o����7�A���ʸ��6�'0�r/�6f�����/�ǐb��8O;pw��a`��m����F��!��
u:�5�d�ܙ2��/�s7�ݹ�|��l���D`P�(��?�2E'Z��(~�	��[�妥!�҆�چ�m�4���bo�69P��8���b��p����2��3�*�0m������睭A��5�dE�QW�x��*%�������ªm�?���cZ1�	��P��g���]S��	���ik�CE����)�*E}�}�pzv�}�_qc�D��ox1����5�_��p
)�.��������_�R���t���.$��u�z�HY��Ed��샆��m��k�ۛ�k��;���I:�YytU<b"�����AW���.�鳚 S3�,$&�K�x�.p�������k��@�.���3]�g��t� h�Dn�)���T$�6�c��ۋo����G�X��1��&�-�����E2u�w֓@���(f僀Z������/	^�2>��kU���3z����3�?l�^�X
��s4-oJR�a������\<�\-��Ѝ��#C$ $�&�
���(Z��/��}>������-��g���*wr�g��1���j�c����	P�7�"�\X�,�֠~��ـ�a0S�n�<O����T�Z���	G�T|�>���~9>�6�t����=�ˊ#��<��'^�l�Ĥw�^1�6g�\�t�Li8�L�E_\�e=$}��x��?qB|
ԕ+��@,��O�=	̏���j����ir<����O��lM�}��u�#��c�[�)\�lJݺe.J�4o�~��[���BT��ŤM���h�h��{uΥx���)�FV�*����^=?��0(T�S��ռ7�|�.*�f���?��������XY����b3Rx��+�f)��`b^<�4ا�ۗ�kƯ�<f�4X��J��*�0%����ݒ��	�~�'1�^�5�,�J�� �'��ȥ����{���!t�^լ�/'�uO�<s�,��?�`IW�FR��Gv�{:�蝶��_}���>[#:��t�;��T��r�K�C�Ah8�M����T�W��?��q({�"a�s?[twXԸ�UE�z3�9QGR��F3�A����9���J$�@(�&oMM�o	@e��P%�j���u(�Oҡ��e���?�q�F�EceAa�vD_��Q$�xs�q�Ԉғ#ꉉͨ��*{���so6<#_�`�@ھna�q�J��ջ(���s��u���.u��K���A�z�ju�Ys �ժZ�4 �=��S�j�a���h����

P�ky�l�w�n�r,ԯ!�m�E��-�T���v�x�SnJ����5Q�|!�b�q�;�N��6^y>��yҘ�z���p̉,�#�]�R�{���':�K�.�d wh.9��zJ�-�ȧwh��.�l�I��	$D����vG5�P�`D�&TY��jp6��s��?.|���� ���e�����J��ROFr���|Lu�y�(s�^O�d
�)f3�	�wd�8��kRI�ЩW��SL�w�3�����[�R�6,K�=��:�7��nJ@��	Ig����ֵZ�%��[�nEM��=�4��|V\%�y����O��^<��04��LqY.g� G�*��(���
I�EI5^DoW���k��MCQu�o)t��u�j���Gd}���]�&��O�Bd%9��fv���x�x)$�YxnM�6�R�Ad-��T]�?�P�Db~���I���c
[oF�<S?+.~���ی+�������o��g����Y0�bxr�X	�Tׄot��h"�a��p�pC�<�.�7^n��}W�O/����P_6��gYa=�8�z5<��@+'p��d��?�d�ʆ�v���m8���ؒ��~��2A�Ƶl%�c�F������+*�DB�ZVߵ�ܒ�/w8��,e2��[��^h�f8�棪NP6�^����|�t7i	��d��;bPC+�0��l~����aZ�*3O;�OҐBWR���������j�,,z���<6���9�Tw�����֯������4�����C�.�r�)�~�#��@�����BÍݺ��hҩ?r�`D�	~���2.Aa~h�|Ʉ��k��w��s�md��Ų䯸1t������B�Ag!�o'2'�����J@j�y7���5�n�A�ں<��^o�ǽ�.��G�+R&s�՜8��479�w,������&��8����Q�� Pĝ�9��~6�q�����$��h�;p���Y3�`�ݱ������l ��v�2	����B�ߍ�F�x��wWv�B
Rv!̏O�;5L6���xM���3�Ѭ�]���4�4k��}�e��{g���p���lF��u>}��~�Oi�́|��m3�،��	�G�V��������1���ᆙ"�*��Z�ջ�N�A�����3���ӑ�j�\�7�5����*pG{�>B|���*i�vځOMx�G��Y�Zհ���w��t��R��/X_98P��DW��c�x�m��Ԧ�y3���q ��n
�DkP+��g�� �E2�X���%�-pJɞDI6�rhi��T����-�-bo�ná�Ŀ���M�^"�!A�>�4���A��PV�0�Zإ��[ŷ�ң�������T�^�/Zq�%�ԫ���TD�1"˝��Z}���5��*L��S�~K�1,���q�IM��~L`f�~�B"_DҌE,3�߆v ��d4[ⷯ���Ȧ��BfoS7���|��P���/"/h�\��m�F����/�+���ů����u�2�Bl̓Yz%Jk�Z�z 0����=*�f� ��;�@?F��A�W������P�.��:�����$�MQ�t%�='r���n,N�(�3R���}�_���������Ҋ59�!�"H5��eNb�|�D�æh_�ZT�Ix@_�u��B� r��2�Ik����r䉖!�Z��Qxz�)[ Z��<$�ş�����,+n�	����뢼W����]�N�0��!=��Qk6��L���>��׀��ͷ�"�q�N�������Utyy��i�J��V��O���LL�C(鐌3fu�ٽi�⺐m`1�/r�K�p�ԝ������b^xڟ�-��^�yU<��Q�]]��6�mh��y��|��Or�k�Z ��Al�dfj�4N��Q.��l��Aϳ�MS��_�]�h�
v���>�c����T�����v�ͤ�������uЗ�8��!ݹ���:��UJAhZ[�6��F\����,����	�B4Y�>%�"�wh���f�x�`�W����L�ސ����Q~$��-�Y�_�I��(E\�W�`�
-�FW)���8��Eԓs)�K?��^��R$BD�Z�9\PAu����-k-I�.�<}y����󀱎Y�>ZN؛�h�_�`����
ã��GK��el�ڀ���z�I����ڃ�RIF�׍I����~�k~�wq(E�L��g�ߝ��ڝ�zY�/˰)��tbt�%#'n-4��'��H^�����(A���U:$S1�[nD2���T���ϣ�sI��!ȶ18<�g��'�!"x�V��|D�����S9CO�����ҁ�-16lX�����JQ�8�A��{���u�_����*0V���\���p� �{C��RY&(��)g�W�Pؖw���Y?�d�an�O=�����"��n���*��H�K	�~{0��q�N�Ϧ|�@�?B�����	UbA1��7�$ZT̨%Oh�V�CpY���J4�쭦�
��j�A��s�@�d���ɊIJ�f~��;�d �-1sKU;��](���qL%��s$�eؕ�	�(���O�x;|�CoW���Pis���Do]���Kd��h�ʌ����r����Qt@����3P��3�@�R�\D?Db\���|�JK^��_��f~x�=���w�<!z�"�^
ZzP��ws���q�&��X�_�Mk��K���ņ)�ٗ-���+�	e?���Lq������$���'}=�n�<�ٸ����C�'��y�"�l�LWn���j�[���lQ|~�>�-�*�s�r����auV�G0Ӫ�3�E__��������h�ϒ�/����k�Ab"���:�(X���^�[�U-�2K���Q�e����@HWb"৴�o�o��Ê�>��� 5�k{��:g�8u�i�n�&:%W�t����Z0�TA�E1�Y1���d�\��s�#���^s���a��h��f�J�a��B��I�vW�-p�L?�>�^��hm��`4�U�|����]f�WA>Ԓe�Q�^��X&k*ch�F�:��ſD����j*T���ßCJn{4�$)ޕ���<�2�j�Zo�� H,�W�~
�n�tr=<ѣl���O
cr���ỏ	!���fۊ/��3(6]1�����$��>fb�|�A������/�����o�!�%���r����34�J����_�)!S�UX �&:s���D����鑻�2�8e�^�����2��Aq���W\�ؾVe�!a�T� ;.^xŅ7PSyi��]��Lc��z�P����˘�m����%���V�����A[@2`�U	\�'�X[ia_����m�rB��ˉ��*��\q�ֈ�"���^r�Q�.�籛� /Զ���V<�����Kk-?:\Ð3����'��Q��bQ�?�#E��hV�Y����vE�-H4C�- �,˓��Wd�e��R]�ҕU����S���ַ����v7��wV�/=��m���B?��7��j���>���cK���`��I?"�n�Jjo���M�Z��À8�+}k �jx2@7 uKp oܢ;Ƿ�r,,��+fdl"z�u�է�����/Kd��e��>��"c�/���5s�E�G�B�%��'�T�ʦ�Y��e���g_�SN5�&���PM�X��d��`��}	���z|}���-�K���� ��Ih@%��m��P+����V?!\�}٨�+:�S����
�e@|)t I[i;�Y�$λ9G�}V��1�dX��p�tJ�n�t��Xg#1��R��IB�?(�o����a/���4��$��Fs����|��G�+N�esV�i)q���s�[Yܚ�n�]�?��궨鼾��"eb��m���rڙ"߆�,|�	+J���1��Ɉ1���ɻ#v-�v 4Ċ��
#�ٝ�J\ޣz�EBpG�>���8��*>�
�O#������q΍��o��>�םӞLn����AD�Q'��m��#ʷ���cl>��J_�+�_,�~�
�ߚ���`�� ��&@��5�L�G/fq�E�v�1�2���Qju"l�V�g����4�?�?U"�Ʈ��,�L�aF��>�����D�qѾX:��S���ؐ����W�pX$gIV����|.3��`1g��%F�g�3A�boe��S��~��4*��r&`8P,ܡb��5�$[�}n�e���"�}e������naE��y�d/0DފK��חQ��m?��[$�zR�,�ڋ�4�1r46����@{,\+e_d��)�A{����ێ��KT9V� Tݜ�~ۊ�鲅I"7l0�؂o��A%Ԍ� �ȁ�=qd�ȚR0��K� �vVi��D�1�3ԍ&tN�#�T��I<�)�0 ��@���O�����Jbȣ���ÑV�rQ���aW�uP���`��"��^����!�P�JD�:�ѫ���UfY�5��5��z���2�4�$^C�J �K�l�ċ����J���AXP�S�2��
[������ɺc�Ga)���s[i�����l����Gx�
��kԃ-ƅn9�b4�G�"iՔդ5��Uɝ�z����6�f�p�¤�c����b�t��w���C���<��Q���{t��'��"�*��G�E���g�ӯ9/�2/�%�W2���t4Ȣ7�����J�J��o��2��Z�+�T���ݻ �{����Z��T��k�_��;N�-�ʹ:ͩ��t5�F��D_�HM��mw��I� �d_��&����v�C*:
��׬��σ�����4�&ڬ��dz�e��� ���٢x(2FB��ͦq|��^;pՏ���8!��$�̃*���L^:�7�:B�8�O�~6k�Æ:�4l_k�Y .�����s͆/��iJ�GL
W�Kz%r�hGf�Kjr���n������"7���)З�^���)�]��J�1������6���52fL�h�h�M��Yh��w��|v�{v�P��U�ԣ���+����#�0���NU7���6�ϋ�/���d��L��d�{��;�J�nu��Ǯ
h�)��v*���K��5� ꅗҍ-<�/���|%��
��ꯛU�j�II�k���uϘ��B���Z��}�\Z�U	1yG���`'�C�	M3���c��k[7�}�u�E��Z#v��07���X��=�i��K�,V��1��q]���ԸS��5/��WzgL�8��1L$ �FBM��5ЯV�i�B�o�����h*�? �U��2�&2��L��0�#	�8i�򦴯1����� ��-�+�0�c�:#PZ���y�2�9FR�{����o�Bϯ����qX�`g|�_!�@5$�ԝ��D���d������u�3�]�刑�`�1�� �S�^W�_��R)��v!�Z��ϋ�wO"]���J���`��-O(�&��&u��;K?Z<HZ2 ���������úO8�����z5����3ϕ{�A��d<���)��Rñ_���Ipd��3�@���jɉ��s��zp,��6�h�"���P��1j�l۞�q_̒D�ߵ����[d���*� �.����F%�Η�Lc`i0���g&��]���MR�\�����]S�A���M�2(&���:9O�q�lꜞӌ+��)\A$�F��&�9���E�����=�̝�f]���f�]�NJ��9g*�Z�m �aa����8�����ܤK��Nz�5&'[�S�O�b�_�e<�C:��I(r�^v��dD��iƱ�8���vi��|p&���絠�';��\M^W�H&�o����9Xk?n0�Hy���k�������ſEBp�T���vN�:��&�}��L���+��^�`�D�fzڤ⟃�u� ������ߝv�Z�L��f���c7���	�qЧ>��ޕnP�64u���I�n�s�"}��y�`[�)���ϕS}�7GV�͔'��[�Lxǵȼ�Q������g�o@�Z��7yI��ɒ����H�1��K�H��M��K�ȋW*���ewɼ���O;���^���2�h�b��p�bx>/R����"��
���aJ4�P���ftt)�st�wI9]+!_���w4%=��4���l[��/Υ�/�M5ҜS,�gA��đ��Tq~IM�&o3�(?�2�4Ae�D$��?Y"���������p����oQ����f�B���$��5i�3Vv�-�	��W,�SP%*������聋!4_%����O�T�x,�ջ���%�62�Cr�l���.2���/C	�tn�K=��*>�H���s�q���0�d+�ӹT�g�q}l��SC�!�YKQ@��_zm���}�l�)&�$�)än��z}y9�(E�t�f���.���U\����d���K�&.�Ս�!�+�6/A��5ϝ�\Lǯ7�� ��Y�^v�]�H�`J����>#y�,"���bY��8��+��<�� ]�i��J���ձ��y�b��d먲9�߯�8��j#�Ύ3������r��h��r�&)�OÚ�Wy_����dV峋d��\���0��{ͻw`�#mj�v�t|�ofW] YT�Jfs��L�����
�����~B���~��� ���X��	��ص�k�d�19ʹ�?�P�=_&o$k�b���E�nV��9�C����Һ�ּ1' �{�N^���y�0p��a���p-3�[|#����I�����=��$����A�^����p�By����u|G|����w_�!
|@x��L
���� ��oXG��:g]���<�d���R�`F{2"m8����1���k��	��?g_�H��֮X�D ü.��<�1J�s,
U�@�����,����ہ��m��m=*:UA(������lg���.t����̕ u/�9��L��<��\ٷ��vx��$�Հ? �JG���(5�<��K�G�0J�a�8˛ŉVh`��.~��"ֈT��@Z�*_LU펊4�T�����&M������'|;,0=�r-�b �coV�R���Ղ��7t�UM�QV��g&n���焦n\K�йӦ`�N�Ô��c�1�I�|�7<*,�:��h[�H�Z��܅���/?���_�^�+�Ã�����h���!��:)I��h�#fi���rM�z�D�4�kJ�y�Q�xQX���-�$}Hϸ����U|��xau�J�m��q+=�G�i�g�f�SQ�=2��D�%�L�Q1���o����I{1�=���S�Z�r��#i#wE�����p_�n�� y�&,L5��F���q�\���UDn#7���%���J"�Jmܑ���U"v��|t��,{��N��������\T9mIE�����-Vؠ �afq����/8ap�|��碈�(����a��£w�ρo�6Ƕ�ǡze�ɴ���!{!�=т�B��nU�{�(���Y]v}��p�Y�@���ݾ_I�O+�H��ST���ؚ�-n{m����˼.��/�$z�u9716r$]�0Ðwl!�IEq*��-a�z���kLAV���I$n�/ʀ@*$eK}+}G����h���rΞ1�����/p7}������Ņu�u���{�U��W�G칏�A�PԚ��=6x��|=4�:u�˸^0]nM,CpuK?���Wb��>�L���ɯ���v<n�
A��dA��]��+�P����Z�
��f�n������A�U!Xg��ɂ*��)w��}�D��ژU�c6�߅��է�H=_�"4?������n�����F�>Eb
��i�����M�B6��*"�4]a>�y�8"��ϫ��15
��`�� M�%O�3��ö��W�E��Y�V\���GuFy�Y�>�p�d�G[�C���e��}U!o�*Q���!߅�dߝ�x��xݨ��sc�?0�+(H'\�z#@X�Bԭ�`�ذ5.f�Ͽ�1����+�cU��0���d�pabEM1x����r������Zp���ҡ0G��}I�3�D6�����Uى�����<��P Qq;��Mb:��?��7�5��&4a�dE���!���6����	��	�Vr��ko�M[����J�\戀 �g��
vc�@�B�-�(����"��j't���:�/�u6���S:����
ӈ o��ߢ��e���C�w��ac�uPW��h�R	T'j��Ŷ*�|��a���W�v�렣�0O0��Jx4d���F�J���W�`���!�h윧��U J����`fܟ
�!���R~"y=:"�����6���a��˥����`��%��ԝ�&�i�h��6��[�2�x2�����u�O��V´gv�*�P)�h��R��W�(+���C���.A��~��eo9D[�&��U>��6uL{ �P�L�Y&��%S�׃;��aA���b'�b�E���m����T��B��Oj��2����r��f��_�"�Z�B�8`��D?��.cȜ�z���
���L�q~7B�m_f%����U]�`F��c�mK��y��*�<$��C�ۡu�k�X�|~��yZT�,�>o]�DU����sJ[)��+�d�+{�Z;�JH�Qp��*{A"hI���=�%eŹ���O���v�Xn<v/91r>��w'~�[�F��t���E�ˀ�|��G*%R�3�U"$Z��E���f�^�gb�6��ڞFrF6ŭ��q�ح�^ӌ�pk��K�Ɲ�K-�m���- `�(�0�lW=]{�^~.�'�
e�����M���߭���!G�|u���9�����㪝w��������X�p�6�R|O�'��Q&��t�������;��׷$��ظci���J���]�D~��Y��'A����B;,i�j4�Z��_�5��5�	p�5�@�uI��}��9rbɴ�Sz��8ǥS,)������W۵`��� ���XElJ���`����>G���1TλF@OyIy��{��f��܉�d����9�CX���B3�$S�l�!�J-��d
e�=��M.�Eވ�\��}P�)@��Q��ɩ�C�z��A�V��Q�N�_'�E���S�pCk��p����E�Xf+�I�Mi����O�t{�K�_�Vi	�3H*�m�KJ3�#���z����4����ҧ�azk`��PʳX�����:�e�wdsѷ�Be�8�G2Q�:����l��:+�� {����#�����=W5�Z���-��1)��He����'������(�#cl��FN��F����Q��&h��G���ⱨ�q]M&���V&�&F�])��;0���0/�	[ZJ<��(R��&�R������ƥ�?�����.=�zq��M"�{ #wsc���w���)�G��Yh���8]G9Ō��L��ɰ���W>!'k�V��9
b������Y2�����,L��ۺc2��2�Ԓ�9D�v\f2�I��K�2����rpͪT��ƞ"����@BZ��O3E��I<����.�LP�8�<�`]X�+��?�7d�d���;&���!�5�@q8�"Q�������Z�dUr����\H��O�Ӈ��q8At����)$�{��83�i9�������OC�l���=�D���M���7i�չ��'�� �'��u�8֤�l�
Y�P�$�q�I�Al|d�;*iu�X��Qf�w`x��l|�`�ĩEA��|p"L�� �!�zqsh�#s��*S�$�H�|�3f2��ч2[l��z��k��KQ����v���~�75�0��Eh�fJp��#�л��Ė�E$�.\y5F��nR ־X��>}�+I��.{�4P��vɕ����fW1%u���Q�%�~ˊ_�MŰ�@yA����K",��Lu�gwg���q�h)�+�&�����l��  �op�X���4��#���s��6�}܆�0C��h0����]V}���@��u�,�~}5�0���dm�p�Q��,)��XO�Q/���;�~��P��iC�P8���N�0��_�@���]�D��3*���������h4����ᜨ�NgC� �7�9Q��;<�˷)/Wt7."�7�6�( �|5�G6P�� J��_<��s����.k2����	b5��v"<YD�>���ģ�7D��KFA{N9���**5��N*P���m�O�X~�}D�T;��i/�YҨ��C�������B�>��]/{�6���"��zA!����@w+&[��Ux����mI
�TU~�����dFB(6q���ʜQ�l�U_�:�0�`�����E^=)L��ށ���R���ϕ����W�����,���&K�u�۰X����ox�9�޾�?C@PT5XhϦ�:���˼�zʷ�y�[�E��ҰSL�
�+��9�o�PtӄF6�ۖ]�-�0l2��@��
�mm���֟Tp�Z��L�j�W�1��K�U��/MZ���Z��<8��G^
�\CT73&w~U/4�'���L2�eery�>��ȶ�=��-���߬i\L�޴����V�Cn�vS�c=k�n�C�X&�����a>,D�za
sC0�~�����=�kڸ�S��x8��*c�SN�9	��ٮ��=�W�q�!�L#u�3m��#�f��o2�������}�'��o�_��6�4(OO�@T�9mB&*��"�|	z[m�: J�9���c���i782Ә�`'m�-������2�<����<%����ő���<w���W�|�EW���;��"�j*fo��Y`M8��Hy=	,\�^]1"�ך$�@�>3��1�rr��&�'[�����b,q�h3Q�;r�mh9�r����E�Z����Q��͢Zbn�#wnu`����|��E��O�IZ��b��(�v7�a�YQZ��C�gf�{��;����u(�K/�h��B�g�*]�X�h]�Q	T)rӹ � J%|�Z��j���	���.Eg��7�jzF��Gp W*�:�e��·,Q�	���C�M�n�mY�vB��"zч���W����!�JpړY�_� ʀl����$a`���C
s��(UZ�^C��a��C�3�J �7v*rBVюh��#��t���nv�L�3����63t�A�gˠJ5�,��nS6�uǦ��,�B�9�,(q_��#�����X� G�!�q���C��D�n��.
Z����OG��i?�%�4'S'�
0ʁ3�a�[%k�"U ��n3�L5�DD_�&6
���`[ߧ��P��B�[?��8C?���\Wx�V��ᇸθ��9"��Q�'��6��S���r���ʧ�����c��拻l(�h�!�X��1d��F��upVv��j�z�Q�!���x�)�ub�۵�G^��nۅe���=u.��x,�0j�AH�j�?�� �~~�gc`��頻����-��֡dɂ>4�p�E� �(���?��K����lTO���ό?xt�y���&�z�����qZ㽋V&��v�������h�w�{����[(\+�)��q��֡J���,?�`衭A����#��Z��!�s�=�^L�pz�z�xa�W܍P��!j�j���h�W~`����s�y���=�Jp�V���K]��4a+e��w��}1xXr$3���@h���p�Or������^Є�,vt+��NH�����p����.C��8#�-y��7ဦ���5����/�u��q�@K����)a���V&s��!g�����+��0b5�c�������v6������]|��sRi�e"*Kn;�*�T���'��ۑ\��Ybc!��4��������N��W���ě���x�뜔�>�V�.z!F��N]֛�����Zm�Mw�ĥl?^j�J��l�������9p�D��~F
ڟp
O����v���h-�V�k�����I���q+� ��c���H�:�]�S�P�&��=�-�������5Á��P�6SQyD�U��0_�/ �5��aB�g.��ch:����:�b�1�B��."q<��"�=-�u��~�\�a꬟�+1���?�m<1�;�U�g�F��޿T@�/UTj����α�,(U/<�1�˨^����������dY�WA:�Qp�7薛<aY�BJ}� ��zic�¤���iB�ֹ����U](��0gv��o��fW�9q4��pE%�mm���W4����2Ӌʜ7��q�����e�Xt�B�|�H����^c�Mጷ�G���^�������}��ȱFn����'�����_m__�If�ǂ]�v2��g]1�m��`:��S%{�5y<� a��@���E�H8hӌ<��Ɖ�>��%�sG�Xb;=�@�X/Jέ���� S^���}d�5gR.��<��Ε�<�x��N����/��1�Gw]:8o30ͭ�SeQ�q-��op���Nr��n]y��=�"6p;K�h&	�����tɓ��0�B\�̮[�nsF�W�B��J��hCK�K�� ���aTB��nXc>&�C6���Z<}�\Q5�}Q�I��$hU�&��I�l�<my��d��l{�I����c^��`�o� �*8|R��3��g%��Y�a3���� +뉂ʔ(f���Q:�������a�ߪ%Ux�KVh!n���a�4G�m��_ǋA��kvu����~��f`����uuB!�w$�T�t;��v��'�Dh���v�7�_0c¯v�e����C���+קDB}i��}?g�~�m��5��=��O�ҿ�]��U�����t��$g`��K�|����<m$�1�7BFܒ�V��k���`sj��*':���FT��^�9�#�õ�O�o��f�<��]9&�a�<xdn}�����?���g����xǷmL�b�"�W��ͺ=��A�hO�!���b�bW��q������i1)
���Y�v��T�5c���8/���К�X��\1�'�@�§��d����A� ?\��ӓnj���� V�5L�\��/�ub2��S��
���hI�l11 _�����a(q�Ӄv��z�R:��
J{��h|�#~�����M��}�������]aO��,NNʴ1AM�%���*'���B[ �6E�%s���QF��)��"������A�)0E���%�����3K`N��	�dL$�ɰI�_�M<�%~�,�,��rv�Q��o�v����*�@�d&-��0���q����P\��D��� ?�zRp;1����QD���������$�qVB����R�B�6�ՙN���s�V���<��"*�����	���"ڃ_R�U���
�F%z�H�G����^�;��xZ�w��#�db�e,�l
��%{m��/�)[�k@LXK�a#�.�ޙ6P@m�:?��r3C[�u�M�G�'��B.s��`��qdW_���@:�t���i�E/��B1�AM	$��� ͵�1�w�6�z(_�q��s3O\�6nkBV����j:��p�#�~�jƌ��Ԍ�1z{\kE���1����`�S-��4��h�����"P��nS�qӘ~�Ǿ�i��>����b��X����h�F�5ѭe$�T��<!B�_p�^���H#��i����-~`�bb��&"6�G:���ĉ䈪���TzJrH��H:�����2���P�@����,�7V�T;�+�nK,P���y�����%-RE���'X��|<b��j��A�������﵏�^���߿Y=��q���:)Yc�ױr&��ڡB�ά�
�rh�~�H��.�E�"Ta��g�4x ���I��d����@$���П:�ӻ�^���{���b�pE����"v�(��������m�;B"��+���H��M��3+������曽�2孽�i�}�Z��O��[�M>/�&8osz�2�2%�+yP������U�SژҚ1L�Ƚ?a�E^�� vA���ۚs��0^�hV��C9���)d@��˲x��m�}2ݍ1�����:�h\⊅�e�C��^�W����܆�H=�,͗��G1��{�?ω�W�i>ɻY>Pǭ{�m-xb����ܪ�d��B2'7X�\n��k�U|�&�+Q��RQ��ټ>S��V�C�&�X�M���Tǥ��t������D�� ^ 
��FD�H׌*�!5�;ޞ����眢ĥn���s���x��;Hx�Ȥ�&�'���_.��V���Q����r��q���9eI��?�H@�KƩK�a��t�U��l�NI�տS^�%��H0{'�fnQ�Yǥ���2S��h�12�����J�Q1I��K�{��Q�z���T�I&cbl��>�F���N��p'����5��.�fFӜ���>]�|�� ����[�M�	Q�Y,�n��_(� ?"LI��c�v�I�w��pA�tɜ�����X,2lb-��ظ��fF���e��E)�SZ�.���ЌBW�ggA9��T�*��
t%��IGj��q�Us�ԣڹN�aUX����OǱ�m�{%@�NTf5����u[�L:-�E��@�����9��F����p\�Zi��@x�!�Qp)j��R�@R@�cb����^��u�&P�=�X���"KH�H����!Ă�^��[��v���5�[�;@̺�wL�,�T<8q���G�&Du�Z�=�G��)��b�bͧ��,�Q����l�AX�� t'�G>�5����D��4��?�&b��ap�z��n�U����a:�g�g�G�z�ӌXkE�t^f�0DU� Ԏҷt��B?>K�I�P�Eh�@�ż渟{�Zݩ����E8��J?�N�D���5�1�]3�;�����Z~���>��֙�H�Sx���:��D���,�sc�<�:�G1�Z�#͇F��\x�/>�T�k��W��ER�'�n����5Ռ�p�&V�PZZ�ʂnI�4^?�s��mo��I����� ��QdL �y�Rd��p�<��� �
�_�f���
>˚��$�cƀ;�42�'ZZ�4o�MR�KXt�H  �u�������\��Hg�rh譶w�Ϙ��k��F{�4�L<�7�h��:A��tE�<�絿c���#,9ۋ���@� �δ���H
w���!��r�.��=�o Gv��|��r�6�T%�8�
Ѕ� D��@�e~�����8l��w�c?et���Q���^5�|C���)	�g�\a%��܀��0]C���c 4��lo�����;Wp6�1g{=ƪЉ:���&=�%����&E�!pv�C�\f��Wź�p�r�,��~�O���p6qʵ���ל@��$�O��S����=��C��"�N�ueIS�R��L*���cwh0��"z�;{�w�d�F��I�s^E��zۖ�\F~�7k�`���t�AN��K/A��czg��;�b��ǵࢷf���J����n0��m�����L�Uc����⑳�����}���_������3dyE����T����AT+Xƛ�h���몜����z�$��?vmei����Z}��t-n���Q����d2(D�aP]�nWX?�EN���T�_��PC6mZ������s���cV�E�^p
�NZ�UTZ8�]{o�|pG�uTۍ�K��~��1��1�_��)��%�;��
�H��bޕ�o��3V�XҧXk��Y�x��ގ
`2XA���/K߲!�*�o1,��
���=/s3Pe�#X^@I>�$���QT�P��'v�_����q�ܞ��E��O�j���P�u-
4��.M�ц��^�"�%r /�!^���<6c�%�h"+�	�ud�9IS�mV�����=]�U�9����d����g��W����B��n�~Mn�z�b����k���E�r��� �罴���;WY���.�j��N*���+��*��ʹ�$K! �Ba~�XG�\V1��e;-U~����&?��-Sizh���On�㯢�!F��.C�J�M=�YEM�# �5=�D�%���>���.��(,�}�g�^d�pW���A���+�5mT�=-��R#���4]*��{x��./	x��ŋ�%W1'�v�UM�/9/;���f�j:�L��d�i�E,bL�:�w0�4���ȎY���e�~仱��%�2���A�+�:�������v*��ǣ���+!6��ٌ2J ;���J�J`����C��sdٵ�8�,�N ��TgC��`
�E71T���k�C@�[�����5�~j��>���kD���c��$�W���[��A9tM���bc�+T$��	z��_�#X��	b����m��e	������]��@��/���8H���(|�A+h|]cZ��+ܤ{����7����.�8=4�6�U��F���9����$�;� �J"ܠ�1���T��VX�M�%<��#��MT3�����&��o�(���3GD�4��{��WH�R��&k�k����Pw�ԽD;~���>�.�
����j����o��Iư�����V���7�Ґj������x��F/O���Z.J�S�ͯ�\��[G5�;
��f3DTק�c���-���<x�:�hb�Nha37�y���f�����cq�)�3�A҈����7o3l��	9Μ�o9<�5�%H�W��-v�=��n�a�&�j�{�2�l ���l��y��v#!������T80qx��(�@������_��cḌ%��{���ߖj�.D�FF�iYT������QU� Z�j{%ש����V�⿯Ɗ�Qz ��<=�k$��"�5}�.�#)����e.�k��|�� ��W[�������(p�/��\Sl(��vvɅ=\45J��P-�p#�r�-��#�rn��jz�~Ƃ��M�h~�w/{�ݿk;�Z&�lP-�s.���z���4m��XFZ�	>�odPE����� -�[A����) �E��z[B=4�H��@���>��aY�*m�`�����>=x���ܙj7�1%��o	?͒t��%v��uT�·"%Qn`d���M�5���Ոǐ�����t���m���7��Gv�X
����]�Z�IȦv�{pT컝4P�����
��~|e��B��'!�ϥ4i���l�Z� ��Sq�����d!�YB�|�N�;q ���WLq�k�G���^�f��X��x��
�<+B�|��T�Ԋ��n�6
NΞ���*t��#~��.7R���nPF�)dOݣ��2�����O�V���Il�T�|�>��c=[�T��W��#o���N�,�^0�T0s洲\����@"�9�P�7��B׷�m(����M@hod�PUN�7�V%n]�
���YH�SF�_y�n���c�ϳي�#�D=�P�ص��<g�+�HsL�9�ή��ћ΍b��^_>���-�u'GwBbN܅��ߡ�G��*j�D�Rd�H�}�I\MP�Z��Tnv����Dk"}�ゕe��NL��J��Ԓ���+� :\C�zڬ4@:�i�pM�bg�U:�!����0���kNxY�H�V���RU��5��Yi�ltK+�����A����䥙��}[�nc8]�3TyppjX�5*~���Ǉ�x����
��?0ʉ��(Xm��>.��SY��3�O�#�稥O��s��N��},D�6D�
Jx������\�e�ٳ���BL]�۪7�-5����7�4��g^�sW��{I��a6� �J_*���z�>[�5��;�0v&^�Uҧ+�ܔ�)LZ������m�,��&uF q,�]��MD��� }ӿ��Z�k*�2�C�O:����FX�oR�*��� M�>���d�|�JM��+㰳7b����Ŝ	��3����8=Oe>(n#v���g��c�(�S���~��׿�R2ԙ@G��I�B���U�{�R�+��(٧#)9��sG���h=�FIkr%���+�#K�-�֔]��XB�x�s}�k�&��y<o��*J�\�E��.�,�<�BVs��]�b�T���"�	�12v�h��"L�4\+&G�)�6�j��G?�hU��������!��� T�Hl+��{D�@�v��������Q|��j�5"��=xC�T�u *NT��L�*ɩҤ��턨_+���xFg/@�(M��.b�b������p��(�%�F!- y�"�0�q�Usn ������s5�	^����ՠ!�Sƶ�.���%Վ	g�Lb��yMnKps�;��V�����I.��w�G(B�K�wLWu�7��w�|Ӗ��Ni��by!�9w�s�� ����r2"[^�`�G���PJ�8s���u
��s�p�ƛ��3�z9���C7�	��t3S����2�ۅg��h3XeѢ܄u}�~�����3�aW^ow����x�|�͹�'6�����a�OA>˛	1q��C0k��8�5��T�vz~:c�4E���Q�(��3ߜ_�*y̠o9�+>�T�{��Q����̩=8Kٳ/I��Dd����LK��]����S�D��h�����$;Ni>�/��0��������c��a��m�FW�� ��ƶĚZi�܊���J�u��:&Q�Zl���6��&���㛠~��i���禩�km�����Ϻ�b`���So4m̞�$��{��<�tU�M_�S����3_�Un�z%%��f�3�^V�+m�T�߉�����q��|�~� �T<����mV�{���0sX��x��m}󾷻h��6fjD��)��C�FT�?�n��1�+xgW�l.�<�ಕh<�.��!ZԞ�B�9��f��޲��d�9�K^���Ь�lc�f�tmV
��|��GAS��#N�Iߦ����r��5�7�Ř����c� g
��h"��
��Tc�՛̉��)�`�ԻU��������2�s*nJ�?�X	�E�˜5���,b�BV��QӦ��(b�g�������	��T���v٩mB�wK�$��duO����;-r�����%�א�Ş۳���b~ٶ�n6�L��0�A@��|��J���J��!aXݟ��{rK.?w�=��֠�ǿ(��o��嚴��j���ة��X���"��J-�K��fcKV߮�Y_�aj�6�%�"��#|ٺm8V�����$}A�$1쪨��&��	����k�v���c�Mo�-�����+��a�v$�ܵ��X��:�,c����r�ywb�V����˞�4�b|1�Yh�;���e@��*�_n�x�0��G(�-��%A�8сy��O{/��l_�裨u4���!�A�^��/	a�G��]�T� �:cA�n�qtb������������~�-z吏�;~V�>5��-c�/aCR�װٴ��R��Vȱ��{�m��`Rb��+tߓ�����x��օ���q�Q��?��l��O�{��3�M�_,��#FJ ���`��e�l:���aL��(�1�ﻕu�v�����FNjU4#�X�<�0?�n|<fdM�~1���?&JFD��������Nnq��5N����an�v;j�G#��M�Ry��b�Y��3b�oN4ԒA%_c������௯Zڭ���o�CV�t���؝;��L_
�c�L����q�7rX�1��0� ;nêQhy߻}��""�_h�B����Z��C1Ԉ���[��,,�Kڛ� �VLt��#x�
�W��^�S�)�̮�P���>���t#b^���~Y�^��_���`�1Y"�S�ը~��zX}p�k�,��oeA�%U����N��ц��Ѷ3���=�	˼&�2��-@xt�1��K��U,ѯ��+�K+�}_��UQ�̹
�<�;]��8,�́�8U�B�B���W�r��V�B�+,H�	�A;Ɲ��x��L��!���X��?�|���Jڈ�9Q<)[�>��zb�u�XZ�Y�烏��i���-ib��xWïڨ�9%#w���9���{���P�".���.`�m��~4� ����ܛ�ά�׉ʶ�) H-��O-�E�eݝc�}W6M�ԑ��d�(��ე'�� �U�2�~K��?3fՄ���1���T�m�x���t)衔-e���wL7OY{:�EU�C�z��&��)��G��|���F-ha�����\���IJ���{�j���w�N�X2�v��j��k����a^ڇ��	?lj;�妔����N�TRF%�h�-M����B��zm��w'�|#o�9J1q���5��: 2Z��)�ؖ5MRT^�&]�y�7�D�E4my/S����C��'��)���͠J�i]+M8��@э�IJ�|1d�1O��;�V�;�ְIfxz0���������J듏���)-ܭ��z��W"	y{XN&���J
^�1;�����3`������Q��5�ѱ�{���5s�N^���|:��۽�g끬I�J�ĕRU �7}j��b�{*��O@�����2N������0� =�~+����C+Ng�3�&�i���жsɯ�~�`t���2C���e&��k7����@��=�M�|��Gƣ����/@à�YV�+��
�M=W�th�T�!.�^�#��t�s��[�p�k�*�.vՑ�i�f<��
�8�=Ƞ�G���.�M��;�e��P<s�ݪr���¢1�f#�'�,z2ϏU�.�&?�C�t�T��t�eq��üik4��baģ��K���^���m�)I��ܺ�	���$�J���_��5x�rtB���7�?t���(i��I=���Lk��B�|Xr�Zϧb9>�_-��P~wD-�x�h���c|��}}'.���N�]�Z<m����� ��-uV����A]���i4���N���( 1�:�S:]\J�vւp�xe�k{���Y�8Ƙ�ϒ��V0DC���N�L�Q~����#
�2+?MG�MYF�z��.�f���s��8����0���F͹����%�i����1�]�����f}j��54��k.���r��(��Yg��c��S+3[C�[5�]hG_~K�&\�Ex��ДΘogeXnc��Z@ϗ��9(�
H�q�-�m{����P���?ۤH�)��R���`�F���|�Y���-߳G5��ڥ��Avh�W*���%�l��0�x�S�
�yR�a:W#�ʵ� ���FC�A�iW�B,>X0�}���y�(A~F2w������[�� ?Wlk;%at�)��=Fq��m�~*_��<VP�hZ�$���;L��zt�^+'�&�k�9~�ɹ�LV���PXݵ3�𷲝g�iTm����e"r�Gs��і�}�.Y��'���)Z������IzTn��/�~��E9�t��?�;�7}���%c���?�ARt�������n����'� ��9G�����L�,�[�P��9��5z�n��t3|e��B��Ra�>YNiM �Bu��=���!O�q�lkx�o�0��s��Yl��4�YN6�EDY���ym*Dq�Ӱ�N
��&<���Q�5��6T?�ۑ�?���&��iIdn�4�>���	Cj�N�Џ[�̸�H�Ys��g��c��R)AFq�𹰜���=��� L��mot�8�p������7�*����ֶ;�޳��F�#�er5@*�j��\!��,VO�qW���cXN0�B�h�^u�O'�y�z�y-��em���p��(cK.�1��#��mI7���n�}�h�_�ˌ��$��.�z2�J
�O�߅6��L� /� 8٭�Ͻ�l1k���@�����:k�1��}�f�<z��G-=���X����,��x�� �v�O2&���&���e����=��b��?39^�T��s�k�`�t�m�Ƿ(�a��
��ZˆMx�WaW3��NxM��$��ݐ�)��E�9t����R׾�&M�9oMH��M�1ǹY4�{}�Y��{�PZ3
菃��͡�E粿t�t=�W��+���~��@OR��Ň��`�Z���m1t�Q��cR��{J�
FSD
�%�W�ɹ�ZK�'u�ܵ�w��w����!�H#¬��+}�H��^�aߑ�`}c��t�H���'��sx������������_";v��δJ�������Z�63��GtfGt�K�["�##%C�w�+�@��S�:��d���\���F��Ϝ����9GƷ+��o���R���O�<#�W���}�㭀MX�]���V_���׬�G/�>yx�P�M�7�(,4�!��uL�lU�> Y%g���a|��i�9g����8R�1�ਵp
�}��;�TS4��X�{���0���:�m��H���Ǩ��|N�B�œ����L����3�b�&��C Pd�������D$��a��R0�@|��8��P%k�^��Ot�X �ɺq�-Ƕ�d��!/1�J�s�?o�o� ��u��4թ%,��q4Vg�Un��IH��@�'�	[��񸽈��$�A80��*uUP��hA䵩��B�o]��/�����fc�_J̎�e�N��b(�G��[.n@���l�Ɵ��I��3�1��MU�/�"�/�c�󣧎ǵ��k>mh�|� D�؝W VIM��%���k��=5Yߴnf�0��^��% ����P���3!��I�w�XZ�'�{��.�c*� �(qd�rW��������g���N`X�K	��˲�B���F�v-\
��n!��w����ݶ�ɮ�Z_pHx�;}�\����*�sB��yI��r�`�C��r�anW(.��5�=j���Г=�##pnMě��5U�6,a�1��1\��g��'S3�J	f=r"ǵ����D�����{YpX��w�c�32��VY��d�a�&�X�ꓩs�u��H��C�Lt �Pq���7r[���ļ���mN�u-B�IO:���'�A�?�?/x�gJ5��>���G�P�&���,�Ѝ��m�r+��e5���������"E�����z ��ʫz�8�N��g�M�D{�)u3��P�{eU�Tr�;sJ1|=�䓻=��)������3�CLC^��������İ^F��Dz{��=��A�%6�=`F�<W�=�0��jtXc�4��������֠�;2EF���?�qQQ+o�Y%D����7"�)\����t�~TU��v�ن�|]�����p�ufW }Sl��ss��w��, � /�� ��~��{�~{�K�"�-77��
���m%��^�)��l;�_�G�����ԏWd�:ۻ#4���>[��i�LVy�v��w~�!tT��nǋۂ����.]�l�<hBVURw� O�W<��]��Z���ʧ��q��2����e���{�
������w�"@ bv2�'E泔���gQ���̠���kPK����P }=1y �!�� ��7�j� ��u~�)0����]r!��� �SЯ���I 'J��A5d\�Y�Zoε[��S{k)�+���i�������O&�崔�Q@`3\��t&x���W�*�}�6��`vpL|��+�C�ð�S���{>^]�O�۴^�
.��z<�]�G���M�E���h�>��V1�nҙnp{�T��J	�+�2v��O�3*6=����0��=&֊꠩�'9�嶎�3�7G}��C4!䝋����L�4�������:��~\�l�U1k���/v��^�-���O��R�H�A�F�-����t7��>�l��#����w ���%jc��*�`�/�d��h �	P�z��@XZ� ��yGD/ٞ6�bn���	�bƶ�8���;���HR�U ��=6�`mṖ�B9��7@E�U�����vMO��-7MW7�|'���\E'�4k�(Rq
��tY�=�pPb��khʣ��W��:-�_m��ӿ������%��&���,� #��Q����u�|&���շ��"{2XW'�IL�����sBR6�_�/�s�uh�@�B}�#%��� ndQ7�p��v������S�{q@�މ,�8]��{Fj�Vi\x�U��Wh��m������oҿ��۞9�Zy��>o�7�Ę&��\Ux������df���Jɡ��`���.�(A2��K�9H1
	f�6�Y�y�
fIg2P�����X���wN�5���5��[�A�[���x����R�������J!�2!H�)�5\D�6Z��kj�h'n�w�?ml��Nr��u5Ъ�/8��'u���QS/�dw����	.��bhDftaM�
kg�����O.���_�N�p�b�GX��6qa�R�]|]}�q�ϙu�ؤEݯ��"��<�/�pO�F��y�.���:C�ڦJ�ʒ��9��V_ī.L��|�^-��*���t_���!��?dK�� ���5ĭ��a���{��X�|��W�����?�KFw�͚&�K �<�d�k�)�����9ik�@��'cx��f
��/��-�0��C� ��ϰU����џ}���#v<��R�\��[R���2���fTc�r���H�V��ؕS�P/!��j"���)�G>��<�n�N</����}����c����SF�\�4�*��Chm�@���cJ�Ԣ�ʡ@�G6��௪�Ɠ���Ɛ�ź��1���>5��&��э�}D7�������m���O��/%��6���t�<�ȹT�U���2�>�{/�����skl�$���Z�P4;�b��Kw�G����[��+�	 ��L�:�:�����y�ȁ�=���5lU)���=7�����J�����:�/>�E���`��"ޝ�������pb)Ra��#���HJ2�@�+�]��lIc�܏��yE�,�@T�]�"@^cP�^���H�1�5�5s��գ�{�	bƵ�g���nR��#���:ze�%P�m��F	��Gt#���}���份a�`�RҢ�����|a��ѡ]p����$�J9�Mn=�`z���>a�E���hee�?}y*I�e�%iH+�5-a��o	b奺/i\:V)Ep툼�<�,��-��
�t϶�;:�z�%glCϺ�s�.��1ln�Q�{�C�&��$wQ�J5[��Z&�B�pwӼ�t�L�����Z���}���Ol���65wl�+�o'Y!)���+����A^\v�*1���R�Je�|�I�`����p�1�-$}<�).���%����Z����N�߸����.�4Nڔy�]Ds�k���X~�_ƒt�Y�Uлs���!!p���B���`�{<R+�[������n�
cA��P"�@�R�a`��6�m?s7&]J9b�a>�s��Y�Qӫuv���-u�0#	�iP���O|��{ˇm��M�{{��?��lUl��W�|��pY*:��3��>g����x����BB�σ'?n$)�K����#�o�n��}=�n+(Ve�%�}3�-G��Q�rS�!\�+���^��ٵ�Z��Y���FI6�*N��4��EGe)�R�t���L�Z:�$\4c������G���9��6����Q0�?@����ą�$���-��h$VL�4�eP��Vǁ�i�5<av_IԦ�zޢW�1���������4�F({$���s�������[1�AE1|��n�z���A7n�1��Y�]-sW����Q�������.Q�Y[�M�,4�_�4�@��Ս�[�n:�iDW�\�R��-������$�s�|�N�@Uv�E��b8I�i��rJ%av>�l��� o��n��L�.CW�.K_y2?װ�ѭ֨FK��^:��/�4�8~��Ѽ����y��ˁ�fFJ!�j��W|��P`':�)�٪�Di�|��4}������A� Y�Sa�p$a/;��u�����U׆�="�.��;�����$i�����:����J�|�k��P���1���^=T�U*M��	_���d<���}�|�du|L��5��.�PB���Z}���2�r;�r>Z�`I�{S1Q*>{�=2��I�*1EM�-�QM�Ly7lRJ�;\���CK%Ă�����0h >�%�F� {�:_ �I�`�F�S{hzD�ڼ�d]7�v�U�/8�R_��Bl�h����w��k�ZP8tf(ˉ��]-eF���cd^$O��B|�U��\������ŏ�Ӑ���Y�0#��_mU���k��'9���̨���Ke@%��p�U�U��A^���B���	v'�,�^�[�����k1˄N���汒I!6�v����I�U�b�? ܖݬ��#��0�~�xO���y����2�*m4W�sK�s�nQ�g?�Z-HS9�L�'xt�$>��J��,��N���f�!|�#����q�4��a��jrC��ɻ�����u��K��E�D&��S���8��hHH�4}����a���75�B^F�.��w{֏u����d�V,�������O��X��D��1�U�T2Ӟ
�Xu2[�Z8
y�P�h~l?XT�:��p��Mu���Y&�s���K;�/�~�N��]�=+69veBo �rM�ө7��axs9��!�^��Ñ ��B��� |gikXY�'p�N��sy%j�U҂E��y'���q�v�TC����uUL����u�U��֎��k�n$�v>��4�受����`ZY��i:�̟�l���ꇗWR(-������oU�+�z�z�8O�ZSC�\/�qth���ttp�����g�]�
m���7�ܴ/�G��)���\��w�e��v-�`��Iɞ�$>b2\۵:\9���F|-�L���@�C��F5���o$K<�q����M�_}��X=�����8� b�ȿ���wj���ib��oCՊ��w�����z&͵|4`Rc&{��CaC��5�Tk�c�L��5���]&>����|&��m@	m�l��J�n���5���m�tH;�f��G��RaRKsDJ�L��������k:>;�Qm�< J�9��ި�,H��C��8�z�/�&VВ�K��ѡT�tA�0)��1�C�FV}I��fiς�:µ�n�Q�L+��|�ۡ��7�~I W=�}/k�f9��^�-�����nS+��PbP�x�- ����s��>G��.6t�_Ж�g���X#BƜ�	~+&�A:kc3��#�w��~Rd@�Ȥ�9�J��ܬ���R��~^��{|J�m����+���'������	󨈤�v0���覂�����E��d5�Slň]�y�y�!����!x���C�]=w���_'�mi�/����ҩ�1�rxaS<�J�wy�=��9D�$��w4�LP�Ӕ`���VR����:r�c�X���S�4���@d��Ϳ\�!$i�5s{Q�)Ѥs����@`aP�|kd���c�gX����s�!+��8� �G���>��S��r�@U�v���#�r�
$����3�AYEݲp*�A�n����@Z@����(x��r�����6�PfV�����u�i f�|�'t+z[����g<�Q�6!��7��_��SÄ��È��܋W������B�.UH4�]5G(ۨ�x4��Hp�&��\Q�ϖH��6xbU�: (>�A" }�pLw6�JpV�HX���N���6^�#-�ɴ�!�k��l�'=m�p'�i!@(�,~L���+�{��!�/Q/`���{�@?�g7�Sf�]�:2��a��ݫ�c��UzY��>eft��}�{��w������1�_f������~�J�Ӈt��5�d}2dDk�i�����2'/2������k��Y�����~��.�~�L�m���}�ͫ^�v���5y�rEֽ;&=2�GL��B�ހ|+����缷�KB���<�������^���!�b���Հr�j����$	��;zH ���˄@�[e\�)�i��9X���DiTK�����oN���;`�K>C�N|�i�3z�e��;=�<m���@�S�K�$vE��a�j������`�e�p`�]���	kz0�lnm�[:A�4�Ř�Έh�����CaQۄ�kոī��4L޸ok�Qh�{�`#\E�R#i^��'^uml�x�M��>�Ǡ.qWT9>W���?�*B��>g�RV�$U|/��i��lrD�2Q��XnC6�
���, p���{��B!b�Z�������EI�j�ãp�M`\bh�@�*R|d�J��ûT[�n"�r��`B�&� �қQ��N�S�D���9Bʭ�t)�ҭcC�z(���3�����.�Y��� A�sОe3].��P� :�NR�ss
� C�*�@1\�?��qh`Gܚ�6O��lNt�E,��Կ#��پ��L����B"8PЍ��鞭�~��}�e�D�5������o[��ʙ�u�c�ɉ�m3U�_����Jk�&�_�n2m��V���k��vxd��m�.����uS��n��uT1�:Z�����I��EVE�e#�l�4����ӫ��{K�6���d"|@>��d��Z��^I�[��į�Mg����#��F:��n0���nd��x�����a�[X����"(�3�2bZ��
z� �Bp�ј�ei_'%AHz���^��ő��7E-Mސm�Ȫ���ϖah�c��_��$����N-���Ҡ���P�tC����n�J�����|�H�nw���%��`�'�����$� x�{�	-/�N�j�ja��#��I�R�����=x[��w�A�V�Z���_"�$�O#xN6�u[��3gR?AS��M��?�F������D��̿�C�rX�;�Ez�:F���n>3nF.f���\���������ʚ�&e�B��Ti���t��#�8� �z:�n���X��v��U��=´Ƕ�(�t��iv���;&�@���7�ʦ������y/I��{ŨH�z�����"�ӄ�5F�`Zeϔ�0+-�S��׈4�))8�½�� �@Wc�Mx�X摘b�/��⣖�X�&]:���k�);��.�W��i����G�-�Ut���ܾ�o���=�4�j��j~�o��.F�!�; i����?ۖ�z5�/\��{k͎r]�I}��:`/���l� �7���l޹�Ӳ�*���.�c���$=+�d9�~(M��AḮV���;�}t|��%wթ)�]}3@b��*ѓ��EH�b�y狙���q�T�����)���D�� d�e%<5��}R����eα[u�t��~ ��,�Cs�\�C��q�o�C��j˓D���y�pf�f�������|㥟��*�'�
��ψ��w\�Jh�`�a3�Ja��i�ѓ�$60�C��4R;�)77���������L�"���I���d����\9���l�����ڮ|��:u�#�3��~�߹1	���9���$�|�G덈�K2�z��6�]����l��x�pcU�T�b�8f�����N���25��!A��WXև��r�xl�^�5�X>^fkbA���i;~�:eM!�!�ft�eMa�����E�A�X�XKhu]9�֋C�{{d�Ǩ��$�����Z&��X*�[!�� ����e�tk*��f��^�i@O��7[�@A��h<"�ļr!��y?����v�]�6qi+��|۫��#�c�\l�G�'�(o���"�"6��Sh�  �(�5C%q��=����.�k�4�Oo�T���;����m��S�����WD���=p
(es����I���zU7rtt�{�5����AU�b�g�H����� �!���"�r�����0Q*�*b�r!��k�͙��|�܉���a%��ÍO���^l�2�;.�u;ލ;�
MUu�t;�Cͩ�*}�������3\~kO�
kT:��*�8�?�R9�d���t�o��~����<�a��|�}07�a�|�rKA�n����[�Z�%�G�^l�+7�I$w�A_�N�_;{�`�8w �f� ��d֖��c{����]޷%	R>����|���(I�,�|m4,VʸLu�V�%u���Kȋ�ҹ� �$�D)��c����ɑQiD���H՜��=T�)���p�����j� �\|����}��o��:�7cI2 �T��+F(��	'��7�ϼ{x�g�Jd���nf����h
e�+�Y��뭒�x����]G�q�(��9�P�3g,c}	�ls}Viq�>����D���d�D���Xd�,���k��Ճ��1���acQ�ζ�5i�yy[~۾6��@�mEi7����͵L=�r�r0��� ]�RR�$z��.!d>��R����U81;����a�|i�nq>a42\�^t!� �3)��W })ư("����Z�Z߰��
TeNp����Xс��b�B{��]��54X'�1�T�0l��p���n�,���c�[x_w�.���t��G1�y
+����ˬ3��>�A4�'�kb�m�G5�)�`�n݃s«�����n��bѲ����>c��YOv�]CK۟�Y�� �2��VA�U�c��S*�^�R�M?t��zq���#O�t��ͯ���;���Ō�q�\A����d��m�]1[^6V�������c}��|y�Д�RX������܉��фb���ǥd��":!��6z�t����쩥֤C]���8%Y?�uV��Bn��MpC�/>���Y�]�a���E�+�eeQ���$���Ǣ�E� ��x���*<,�+��tO�!GbV�~x#�ͥ���9��P��:#֮dÆ(ym�vV�x��,�-���
��� ���ũ�'W�z��i*3���� ��GT�\�t�$�j뎆Q��z+���7�`_嫩|���F���T��/��8$�P��B2y�1�gb�8 O�p������d����	7F@��� ��v�^?>��zx��I�����P��a4�2W��
�A�˥��	z`̴+6�t�)���� �y�!i*��<��CO�,�(F��ge�q-���EԹ�&����3��%6W�	�j�-�}��36uQU�74=d`��t�V�
݌E�F�'M�W��K��N�/<>���-!�T��9{�4��㫖.���>$���*m4���;>x`�2oHE�]!t~͙Of_���P�6�����SkP@#�&�h���gA�ĵ��.�WN�E6l���n��s�r��[����vm���) �<�g�V�Ϋ�b��5�jЪ�V�tM�0-]�^u[ɂ���cgٔ&q�a<������t��$`M���dɚ@p��u�(N�<�r������6�|���[y ݼ��Dl���'� NҠj�� h�����X���x��G[&�L=�"7)��Nl_��GX�͜Q�!İZ+J�0�c��$���]!h��5�| fMS�lQ��\Ur,|��a-&G�H]]��}�m�P@�uq����"���w��,�j^9s��Ԫ�2i?��g/.P����z�0�S��^X}(�T�����^�"�~�֣4��Ƙ�3k��c:[5oݾa�5���o0��
G@�fX<DH�;k++�o��A)�Ǟ��aF[B���g�L�;��\���7��ծ�?����y�5�E����tZ�����`�kA�7�G��(��ȝ�X=D�#���^�'��s�@���H��`�""r��;kO����L�8s~�=��Vc� y���<w�y��X�4�<��_��������_��� �l��)�3�W�6�9����7�#�]�b�K�x�GG}-�yǊ���L�)�'�����ji!X(���A�T5�~����I���OS4n#���� �`Q�T���D�+�-�N�t� ��b+h��H���V��B�>q4Һ�Gp�u�k��#�� Q��w�V�1�����z�! Cv�0�	�[~J[
�/�r,�{RdEh�i�(�7����q��wz��A#�z�4��O��)�-.�B�~|�=�^��.6q�.���݌�>��\�gބ} 1/{<�
lDm/�=
�j����\v���sB�ն F�� k�p,��hJ&\\���u_�4�+��)����A��#���j2��R���Au3v�x�(�n�E}�it�=� :�NyV��l؏PU�N�������������N�,Q`��g��g�Jz
%{�(���Ԧ�����Y�N�Q=̋O4�M|�d�Xi�b�f��i��*��t�*!���;�v�~O��
�2O�[�l�P��Ķ�T���p���Xp��'���+�@��+��0�nY�؄>�̩v�N�T�~������΃��G�M�ێ��eCZY� ��W�Ve�� '˵�RP�Z��֮`�Yt��Uɶ�u -��@�ȣ�i����R���U0&\b��9���}���ΞcK�����)��QlL�/��5��x�3��}d\6Ȣ 
$pR|��{�]OJ���}\�6���/�.�\~J��6a�(	�p66�Yi=X$<��NB4m�(Z_����h�/��V=�ԻT�ux�绛�@�+��&r��Hm��%�4�/KG������[M
�Dh����������?ҝ�«V\_愁2UJ��ssHn�s��(D;\;̾��)����_@�G6?'�E=��p4uk�;��+yS3m�3"����H�\��f��ȗjǄ�Z��'KoZ��FSl��!�fh��LPG��gV�ߊ!�xsT�z��7�lZG*�3�����7���8|q��r��5�H��&)f��&	(�UT�?f������jWBB���{s��x���si ���;iӈ�[�護D6�����6�.��J��I�qAfc:3&?WnGY����b��=�G��Eh���)Pr�{}g��t4��r�Ü�PR���Zws�;�Įd���,���]	����vo�ZtC����J7S�5x�>������Ds�XB���"V�qbx..}ݟ!OqD��<��
suTՀ)\�X�6WR���a�Z�O7�O�(�a�Cɭ����ގ��I��Oy��=�&>�ZFbɑ����@&��,�ٔ�(�\tN�.���u|[U��9�|��$H��#�����*�,�L��*�w�ۦ��u]����* /&�	�K|9��D��Fj�1]��ZS���O@��9����< }��u���XX�uYZ�C��Q�U�=��o�+病EWO��oe����:E@���,��H��Vf��ê��'��s�Ùb'	�G�@ ��r���t<�{�@�-*��j���L����6�\�W,Y�uU#(e.P�U�
bB)����H��� "�}YZ��DW��b�P?��f�w��yɜin�z�4N�����g�� 8#7\�?`y�W���O�"�;"�_�Cu�H�W%��NٲN�t����P����F_�VJ�	�1��d�~̗��I�����v��%7�"���?I`?�"'f;��~�|�2L�/j�9�W U	��Ȟ+6������а~�
�1+/�w=0kq�@��;�˝�	�����6�fB-��i*e��Q��͚8�������� ��=�Q�8A�|���Q¬����~f���^[��RN�fP���A�+�"8DqIl�6�Z���+u?Ҿ.��'li���B�W�qW�U2[�"IL��&
5��yVh��ou����v�!�џ�W yfdj�͜��������ZC��Ҁ �|�(��b�atyD>�:Qϭ���j�#�&y��[ʮ��vF�3��?�Ǥ:Cշn��Ia9a���D�{��b�ø�i��<Oؤ�_Z�.�̘^�yR	\n�D�ӵ�����_-U�Z�3`�����q��L���r*�d����~4h�B��-�8ꪶ��AK���j�z�V���N%��b�d�gNv�:+M��ЧzǱ��v���:!����\��ܟp%��f6�S�A)Ϗ�"��l��	�`�N=�0i�)f����������wƹ�uPT�O��Eס���{�p�Qe�����LA��`K�G�-��j���J}�2�o]��}7tb��գ��FB����reh�����6�,#U��"t=j���9��+��y��U�a�(ڹ:�Ow�u�ߐM�Lף�R�;��
{q�5���n,�Gm쒡R(�M��;�8)5�d��֔Y@r*<�7��VOS�0I��ߥD*���޽z�2
�~�az��'��S�g�f~���>G��}��C���=�«<�S�uک7�������X>�!��+A���G���o�B���f�e��ONUy|뽋��n����!��s��zi�̍)�d!j�O���7lV��<����&�N��ӹZLxI1ʊBZ�!�3N@�Xb#<E��c��-2���;!�������� ���j<�����buۛ����v8�F�(����'*������g4l���̓��X�͗LU�[� ������2��ݘ[WP�&�3��><��7�#U'�M�ي��*�E���f�t�8V�m������w#��^�	�ȵmKm�	�J׳B)4;���>1�q�1�Y���5������s������_��0�%2��
�8e�g}�
����[�g��R�s�8(��e�ܦ6ؘ���S�Fh �w��1.J;�G�jQ�9���O�[]nN�����Za�̿�<���ӛ2�7p�넇7ƥ��$��c����c"������--�XE�.��}��1��]U�`Э���S{W������[5���G���p~�y��lL	�>�JĞ�˥��o:�'�sr����zE�:B�E	��(=����b Sԗ�?������9���'�L�9ˠT5�[���	�?��"g>����uC�wLڤ� �J������`�+HO
~]��@���34>Gpr�� XNpj��y���7V�]�Ǌ�J�G\��qʞ�k�C@�XC�s!�Tm�c��G޹=S��v*k����eڵn������V�\B��|lo�]qr���EA7�Y����X�,�G�G�>;;q�G��$�P��ٛ�.�F�Ly��pڻ�?��i�E�P�W	������RwT���b�1C��T-TD̀��O�C8���	�����DQ�4�h���-Cw�3X������'@;�����&��`7*�>��XZ�w�坦�x�ϡ4(b��?�	�O��|I�����K�ځ�rŕ:�uݍ;@<�j:���YE_Z�ls��{��P,����l�n<;SB�N
�(�Ęq(�`��S�G��\�1xX���vc���=�kF^(�L�n��ٯK�!%�c��[0�El	�����.{��s:�Yo�ɒujWGr_8��$�*r�+��� ����͗�����Z��1�l��,�9����c �3�/�SȢ�)�v�)Mb6��<;nL'����+���k7n��u�d����*�I�y�tKݔ��+"c{.ha0ە)3��7�ᑶ2�D�J�S7*Z�e��4���b�[�:�kb�(��`��R�;"���.}>q�M7i�\�o1 #�'�{4r����K���!5`$5��������%�l��s�Fb�����w+�ĥ2���P�F�x�!�?�}�h�4�+��iF,k�>E�:8^��^�-	������,���j�_H��>�v��A8��+�Y��y �w�y���̊����F-���1V6bj�-Stg*^�@�B���9�箠-'�J���|z�o�g�UR��S��Q��ǵ�8*���|�I�=�W=�\}���p=�x��ͅ�#.Tp��:�t	�QSc>`�D3���ҳ8��9�RG:�� �pU��+;��������K�=�!�b�=�S�"����M�]���	X֑$$E�Wu-򁞰ES [�T�HM�.��=��#P��P�>f�-^ �Ih*\cf�<1W��I,���M�O������B�eZ�����K�V��U��c'���¦qGJG//��U��ֆd�G����:ȋ�Ƹh��u('*! *������T��/����/�Uҹ���BW���d���I�{���M)�xE��?:N m�e���-@���v�>�����z.p5I���8�M�6D
)�����pz��l<t���u�A�f�
��l�8�#�t|t��`��D�F��2�T����zY�??
�
��)�uE^��<K�On��n�H�+p�l�~ [��D�[8�Í���rX�C�DB#Z�u6s���lԹ�o�	{�uwWp�KM>n�V�|�V�4?���Q_������L���4���8�B����o+����=I~T�1u��e��UA %3Z�l�;���7b�ه�
�I=)���@KG&���K�(E&�/����4�F?m��NX��xn+��,��S���A�RXty?kڒ-M�y���UHò��D���_lQ/�:l��r D/x��R��X�~�%ׂa�� ��! ӳ���� ٪�F6?����I�<R�������Ӧ���9����~듑s���cڜHE�W/VD(�  Wx#�ܠ��:��½#><T�k����!ul�m��7�NXn@D�:�#��mYle:wv��Rh��'��5TD%r̮:2����n<?�N-l��^<FN��M=�UɄ�&���� in���.K	9Yht�����`3b1��H�3>����et��|�H���2	e��íѱ�3�9t�y��S�'D�Y��ME{��aISs���ת���^�<*�p��D�zS����s�5��~�W;U�1\�A�r�}�'��������Ge�3�_LT�}l͵'�Π���k���VY7�A�7����"�}&����_��P�@�&�F�0;	w��R��H�����0�䷣������#�7(��>?k\;ŕ�sopC#
^#��� uarL[���w�����B�	]l�T��.�Q�}RZ"�ֻ�n�N,���X����U��ʿs`�JF̄Y�������0PƼ�Q?N�\ߺ�5�QeF�Tђ�NCf����b5|z"\5�7I��p�n�T�$bt��:�Qq�F����p�:y�f��z�G������A�,��~��=�?&o/�ԡ�-8��b�wM��/�Yai����Wlh�r�TA���3Z�&�:�Tb�f�ZP��Z��G�nN&��%�x��wy0�<La���Y^:�+�Õ�2z �Y{�H �%�ҏʴ"��d��e)��,UdK0�æ2�z�nD����梓��gyC����Ke��q�a�84�9�g�R|^	���&� ¢��' �8��-�$:
嘸Ҿ�|���a�u��#>N�jT���"`z�%h��^8d ����x^��"�@ҷ
�O�v��;(�Bj�E/�br����oY!�Hv)1L���;8Y��V�m�E���O����l��N��^��T���x�(k�:p�m��q�RpkB���LJ)1]"��ʥ�3e�h�YQ�CO4����SFP֭+��Sy�����XQ6
 �1��+T]-�&������an�Jhh,�<ܬz� u�i�^xP\�*�0F�Z���DU�J�!~?	��R��o���"�N}cq� �.��Μ����<_!��/��	ة��X��;�i�P"�,�;�f&I�OTN{.���N9a��r�6{����^����q�!x�zؚ�4�Rq?j�y�dZ��W�BAN�r�ی:��&W~]��ޱ���}��7ϋ���Ԓzo�fT��ǃ�د�.�]���°@�;m���ťu	��Q������葐�~�٠������/�v��E�)�7�V�,���o��Q� Wn(V`�A�����q;�%,o(��l����~��c5L��P����fc���o�������=7�MFC�d�sS��R�P�Y��0`p�H1�E ��|7D�M޳V�J�Q]��A�i��Q?�*]8���8�_G<�ؙT�����,u���T1��Ӽ�:�V:���E��y'a��-z��U�WUn5<+��4{Jj
���
]���u:v�/ͤ�!�-�l��r@�z��������m_���(�o�����ѶS�>9�H`$���y�7�!lVQ�G{%�/�0e{�> I/�9/��<N
��F?���|.����AV	��Z]��px��� -??�rY�pg]�� �jw&��|)MF�+�� �h.�������`=�>V��`H�����$[�q`ό�)٭E!�u l��+�/���G�����ˏ���� �D-L��6-�A�cj�|����t&�����T��J؆���]a��a�����n��t^/`ڹ� 2b���A��%�n��$l�N���
9��h���zƐ��I��0K��	�(;IF4FP7aP	�l��TO#�k/��J���Td��E�$��> ��T�ڠh�����+�[2�mW�tʋ����J��)p�}���а�6�m�O�_縩.tf�� ��j4��=���=R��W�%�<=Vț(�M�S	HS���M�*9V{�*׹/��V6��28������#��z�.e�Q�\Yʄ�CXJ�:vOdQ���xZl�@0�%����TBҫy�KDy�h�y:�OM���]�e��X��d*�$B��ܢ�b/�Fv��n)P��rE�=�T֬�5��Z����[U=�/��\%a?�Q,x�3������g���cµ����?e��q�^���'@���d/*��_�_�9�fɐ��MaCa��>�i˕,���q��Od�i���-s��|I�*�h��u����M����}ث����,��J_�=	�c⛰���l$FE��{l1�|B�e׮rBѱǭO�5�����3��:iz��J�c�5�M�#`Y.���qU�L�/��P�=&�"�>N�҄��%/�5I�t�|��K}t�Z�[�[�����dt%G%�|�Zۤ1d7�I��Fiv���#1�M�'�^��Xȡi�x`i%Tc�ZA�d3m5��>`<t����L���cH^c/��f8d�%Y2U$'Z�6�iYci�'��I݃��c5��3���(�k�u}��umH���	�)O7��q�1� W������E��tC��<�@�y�V��d *4E>����z�b�0���k�#| -�\Ķ��Έ�xƪ��si�K�8U�߮���H�HO}ҕU��,��%I������ߛ��$w�xJD�W�i²�B��@�*�v�����}S�(���	t&�]�qM?�z���nъL0�#t{!:�\6j�δ���ڭǄ�xێ�$`ۗ�Y ���������t�]p���	+�Vu*�LΒ�6�~n:�!��9���=;x'�p+�8����#��C9Iv+���n�<����f�A��{��� �\���xi�~�}�?�07țm{t�h8�dK�4;Z�M����Ak����S�5��*XF�Y/�����P�e�
�[Y�K�uj��#|�:R��$���n=�[0�tP[�.�߹a���6�<;�s�r�����˵mϔal�'
:��~,Bx��m��\��w@L�ρ�Φ6��3�=J�8X�\Jދ�v��b#?��Ql����.bź��<K�d������Q�:�l�40gQ1�Za�sp-S�l�J��"���˺�k˸�+�ֿ6����,՝���C�/��4��2a���	��õ�f#�����x�z�m�M�0�F�:�G���&'0���ʎ��#N�g4����Vh�^�,)V��_ |��N�`\J'��_���Ԍ��!t{fW�U>�J��ܦ�.���\��ֆh2Vl�X�:g���W��7p���y�C���!^�@���fb�g��� �u�Cj���L���KI�p, �5�n���iN�������	��nYA^ґB�ɧ����h�!��F�>�X�$xT�T5rNƮ�0���`�K7>n~ge�;M(�Z[������a�Hp��ސe��2ϦQ9���c�ܛ~�3T�x�ό�%&�v�V�7��Q�w�K �|���>���
pZ8�����Z%��Y����Ab|���
vn�R��~��wy��c1�ޞ�|�X�F<�<A)�jHު�a�*���H �S�����3�������i��=��� F�Oy{i/!U���*��_焽�x^0��ym|�麛 w9b&�yB���F'����(ز��Hxi�)*t[O�S`��s�Ax��D㉌堆�\�݁��۫8*3	�s��u�s�v{�W�H�����u	]��>R����g�0�5%*�6m�n�x�0t� �Wi���E��LR!��3O�˘o� ��W��`�;�6,9�=�����
dS2^��gGu��E�H�\7�jh�V��*�,	c_�:'����sC���&g�������eʣ��\ [,z�qh�:'�<k���Kb2K�킆�(�(��u̶�#T2��w�1����;���%�.�n?�ݔy��tnH�u3��oȏ�$�,K�(�a�7���6|��M3	5�R��DW� ��T��DB���B0qD�״o��4�Q���O]Q�/B�yy�AR�j;t�XC(-g9w|7�QД�,-�j�����fڦ�H�a��s��� F�ޅ)ԑ��;�-�����9��݃j�FTro�R�P�PM�~I�Y���(��-t)�E	���lˌ/Nd���;�*�s�T�&��"��^��N,r�	�R?�vy�v!���V(։�sq���A��Ŷ�������O?+��s����0�9�o�׌���ҍ���m�:��Kt��5񴾍)�P#�4I��hN��D1r�t��H����k��%�A����*���ŧ��.O"� ���o8_g�E��YU�?�M�
k��o�\4�o`Z��*��H�j^i%3�\Э5�!4�0��}8;��T�^���޷�=}�ɧ��P��K�l x>��-����~�&A}q�	�g�oV�V�,5�,��Jژ�� �5�U^47�/!�*���~�}�Jwи����l4��
k-�"�ʋ�x�$����ʷ����7�D�kQQ����버�D�S�S���s�׳on�
�l�$)S/՞�S�L�(�ܑQ���4�c�}������NFl���7� �C�fF#����8С�����ŏ�
J��L��;X�t@��D
�:~⡞�*��/hD5l�j|JR���le)nx��\��+�㇪�((�H�`�!�+@�� �1�I�� N���7�̬h�d�i��-�`:��[��~jc﮽���=�̈��?���-fE±u/���1*z����'מ8̸h�יּ�α�Z�3��½<>�x8w���8w*��Hx�}!�J����_b����T������oQ�i�;U�3O:2�r�g̹�#@ڑY6��@�U�#�rG�Ndԝ�H�F=\'���C����]rK�����Z�g��'��-Pv���U<�H}�XNJ��Bz��%�����9�,�\�f=�o�?�{���χLg�O>����l!��������M*hW=����f�%�w�*�� �LTT	q��h�u��I9�][�"�VB�m�Τ�h�
H3�\��D��1q�{�o�_$���$�w�p��E���	#�<��X�3u�gV�X]]��]�@�W϶�B���$v�?����'+�n�J)�?�u���9n�����X�ica<vʺ��V5�t�3�z<Mπ��av�#��S�~J���J���se�z}�T76�c~l�^#�5.�;�AB��u��C�[}E�Wgf�宊�reN��=Ϊ���|�2��,�W�����	�|W�k�V�-4vaC�;��	�/�?)<�,O���b���]�O0���w��	�7S1��K�[�_ڈ���ꐖU)����UIA'�X�amq�n_�uNi�����R�i�JC;�m��@�Sa���0�X�f���� %?0J�7�}C�HR�fS_�1i? dh�[#�<B��p[���(�*Ji$�b�K��?@Ԁ"�~k�)�.�%o99�>p-:�ҟIӒ�K��*��)�9������<E3�)u�a�ʹ��C���B�׮��`��طڦ}�	[�w���)s��arV�R�Y4�.�`�I=��U�������Q̙��(�~W�k�����ʖ�*NwL��e�Rηv�z�J9�ޥ�<iy����o�2�N��y���cF�֚�.�#��y��v� ��^�>�s��a#s[��b���%�����ۆ�9Z�b�(��/r�����k��|����V�@���'e�̊����W��2�5m/ߟ^�~��ؠ�M�GJ���E��T�~�suw��T��]��y��C��6@�2�W~u����CT��C#e�_`��w|��)m�{�wq� n��o��1�a1���H�O�7��ksS�,��D(2��h��3��y�7RPDr�٪%w�)�(n2�<����r�E����͹���6XH���A���#0}�q0=
oh+�?[�L@��c��X|�VP�QMp{��]L�k�8�[�E{�ݴ`�3l �H��2;�A�Fݦ�lZ=�(��?��M8s1#���]{�/S
��']?��C��>�.��WkX�.¨��'�˸I~!Ok�U�$��K
ӓ�g8�+N�֚�`�j�9�����n�s�M�c�2�q�	UL��O/��"*��Fa�!���J�����G��2�Svc����ɝ�&���2�nG1]������~�vI��5�c$g���[�ǳ;�v��H��^��:.��tЈ�z������P���؎�+J�5_?'.�.'v��odҁ|����0�s�Q�L.?��󌦞� Û�yw$��4�u���:��	�	=)���͜����S!�H����Z��c2}��Ku}�c����|;�`�M�qb%6�)��].2���N��f���~`��0&�MA�ȥ����$�T@m8Z��������W@�j�̦�d�>���9�M|������s��r	zU��dph��B$iSz� ��Mu|l�+��7�� O|[)�'�TM�f�V �d؜� ���4�?�E~�]�k�Ϩ�����*ruV?�T��<'p�B���`Ӽ�~�O�NEHxoN���殝�o>�K�]\��W�&�������:��􏎇�C��~�Rkj�i����� &+�P�iT�Q��6.BW�^�6��a�p6����H���-ഝؗ��E�{�8`������,�~,��;U�8�Xd�c��.���'E�d�U�����V P}T�nT�$�=���H�p9� �!�Ŷ$&��it`� \���x8�h��tm�ēD;%YI��[�٣fy6��9����n����]\�7-����t$����˚�#��+�_��v�v�	�a�~�Hّ�7��J�8ro�p��*�]t>B��̴Ƿ��8{�^ ��/�̳��>�3ZWdo_أ ��|�4�wi�k�����<�RG'��g��
�Q.���weQ�l7��n���y��#��>2dg��ߣ��^Ĥ���U��?Z�Iƚ�LCH���0�j��3HAW)>��̴�D�j��z^1-�9�9r��|�'Ϡߖ���Ե=(����� ���$$�^�L.SN�f^�b�/��|��+3v����#���?t0���Y��w�Z���/%x�Q-ù���',�PB�'��w�ȟ�/d
h�	\�;�4�`LoNj�@#Sl�Bmڳb��2��D��ǝ�U�%O�,���ٱ4��a���o!]��7�1��]J@\5�aL_0 �i��L�s���ݑ�2i{�N���*�\�#�maϱk2ՠ5bPg��k4>�[�8zσ��Z�6}zC=\_�ʗ?Ƕx�G��s��Rot~���Ev8Z�d�Lh"��S�Y��rf���H�a����Sts���M%d�L�O��`
�	�7���X�Ԣ�	�ʗ�h�51T�;*v�І2J 3�:释!�2��A��rJ��`�;e����?��Aٔ�;�a)[��/m���2�I����r���9z4a��+YS�!���#*���\��48w�M��+�V�9��i9P�i;�1��UHh(Ɓ�@cl=Kl�0��I��J�P�Y\C��h�ϒ7�������"�(",,�ʾ���Mr5+�v�Ho�\>�5�7������� Ob|7<�Ϥ�a�
���H#��w��LǓZ���;L�����H����cV�(x�����I�~BZ1k�t���ĹLе'sY�]�G~�{�nz.h������Q$z� �1��������l�Tn���'	�{<v_!�/L�j��<p����؄�K���ά��M�e�:����Umf����D�G�ͱ%� f~��̬���?����;<�S��l��O�%n��G�U�)��i� �udM>���q]��Xg)d��ԙ����1	}M��[ �m�;�A�7 R|~WҹWshң+ܶ�c�Վ���H|(���Sp��q�ϡ*Gُ����d�ۜ���no��>!���u�ћo��>���sk/MY֖����mez3gոs�~K��ނ��ڹY���d7��RLOx�x6<�s��/#R���Z�y��ց�	2_KE�N���5��6���qa&4�Tv g��.Tl�h
۝�z�>�7������kSލ�Ï���r?rQ`s(.+�Ҿ� ���1<��>w<�^��X���(�M��岻��an��ا��C��L��V�w��>MM%lY��;�%)ds��Ǥ#����s�t��8��ZB����I�~af��B���WC���o�:��GP�ج,��$�`.n�Բ���'�]����v2.��Q��o3o� � �t�#�Ad�~| �4T+E��"&6��Jʤ��%�@������z��7,y�
F�z}I!OBi�������d�YF�a^��(�v1p��B*70c������mI�ٗޛ�ndD��8V����;����r� Ӛ�Zo$ɴu[p�iotʞ�ȣ��(���8�o����2��W���EX���|�9����椆`�Y���� �L�1�o��t�W1��5�BE��8�ih��q�=/��1㫙�kN�[(�x<�-�.`�VM�Ve3i�����9����`�\1��^�.�z�#�Br�}�d��b	˺g)8=a�S*U�՗Um��$��k˪�3ڥ8k�Z͑������'HfT+u���	b0�M���2$4E��C$�6����Q��j�+-��qt�4�1�M�; ��)�y�$�Ok�����