��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|ḱ	I*� @�[X�_[%uP,��r[��n�G�:���e��ի���2�\�.��[s)�>h�0�����,�Y�y��,�.�]������_�(H���h�Nts�_�e�L��A�!�K'97&3s�h@Z�xC�Ux}���y*��9���(ԅ�^Nᨽǆ�Ϊ/���=�ƶS�XjX,���l�8`���=$>=��d�6��G�o���̨)��N��jtDQ���C��h�;b�v�\\O;�^']UJw�L���J�<�>�f��E<��ӓ��Ɂ�UD;��	�_�96�-A��+�X�}{��*�"a��~�L�r���P��L˼2O9`a��k��0��1 49}�1N99:OʻԹY��uO퐜����JA56��A���$�D~<2 ˔���=�h�M��L4�	����?���yn0���{�~��?��j:)�wU"1GV��)p���,��o`�A�^x�|�Vu�=�i��'��K�Â�E�cÔp��⪙<��iO�1��t���v�s|��[�^���ŜQ�g&�J#i�/����A@E ���u$==Z��j�:\睷�}*|n8k1�U�$
鮴�
~ax�_��;5fsC>)j)��iFE η�<q2+�W̐�%�c��h[\���՜�{/�����p��,�.��
$�dM�a���Vp}\ࢸ��\5��5��.��&�|�/�>)k��|J�����J��ʭ;���נ��y8�6��J*N�<��-�����m�C�O[����*��C�AD���!�#}�Ѿ�p�۾�ЇyI�_�����(89B���KV���y�M�v�@���Sj2UT0�%���Q�(���z��,Nu��?�*vg?b���Xw�_��\6b�I5!����3,|�<�Y�r��Y�)X�X�&_�7�s�OI�M��͊�Ŋd�Zn�Ci̅.9����X=�ȴCŝ:��z?3����2�+���3�[���Dw���I`#�Km׸.Yd֤�s&^o��`���a1UW� �`<��a�$���	X!�mʧ����!�k�T�a	��g{���`~YcK�f�B3���^���f>�+�۬'�dgz#Yz�V�i��s@>o�n��`��>=�"�g;tY�B]���^P�fb�E@�&3�xW��#�G0?�MM��=m��z�r�y�ZZsğ���GK���`��R��3�J;��
Ŕ���:#�{�4T��O�9#�ژ��z�-���lP�:/\`�<��n4��"a�i����Е�|��ӟ��&����#c�  �+Po&�$}D#y]��L�0����A�3MgH�����y�si|X�Ӣí�R�L,%��fmzHV�e�4݆O�x�An;�w�֡b6��Z�����'j�Y�]�=Wܚ��A���FN?J���x��$��n�҉�O�G�����Ǥ���������I#�k��p�p���>�\Pb�6�tt��j�4}�%I�a�_�ڛ�A���(��M�C��.��A{)���8�� 0���*0e�r���e�=��Z�Pǉ�������e2 �Ż�wL��|�O�CF��ԝ�DD�P=��!�[�������J��ng�0eT=JTY��u���6�5K�`��ڼ6�+l&��mW�����m�Cf��햼��G�hs�:4��a�S�@!���(
H�[�\əR��Y��+�ME������W�2��@�f��d�a<��SE� �%D*�{`���=����:|�T�]�27�.�����l1��A���"���K���6��Uۋ�z���J/��.�JV�Q#���F��K����13P)��"��I�V)�
=z�z���u��Or���y��q!5���!�譍��.���
^�(� %�I�sI�j�_�!<z��R"�P��� -D��S�i�?��E�i�Ɲ=�?��O�3��ZgL���^�,��q�1	`�z�|2�����=��QVY�ܦ���;?\���9����Y,8&�Z:)�359�#[S5 N/"츾J�9�U�|�f����N�hG#}M�q8Vz�1�zC�H�i�XG�����z�%�.;����#?r0��%#]:
V��w��]8c�/E����BD�m����8FՎυ"=����R�:BHK�:�x)�Zh�q�~�e��`��2��w�
��9��WDX/p#QO �rf(D�����Ƒ��)69�#���	K2����@���!:jAD�bp"Hd���c��	�{�Mw���pm@�`�9��qK�(
8�×�M5r�P[�Ð��p3̧�:�.A��� �˯��B�/�Y�5DaH�cW��=(|�ҭ����0��ed���1�/�R�)w�k{{e�à1G�o�F�S��-KK��,���"TU0�o<Z����,Z'��US�"_�6��BO@y�[��F9NlE�?�{�F�IR��CK�w��]�f�xh�k�o����Q�
UCM�-�!o��zC�w�}�0_���j���v��J��^~K���:���sdF��f�=�Y6��s�(r�C�w{Y�+����;����,ۜ����°m��dt��P~ ���A��v�P)���!,���o���̸I�$��&z�q,��]����h�xDT���uEЭ�D��昊���`o�����\�V*�y&���p�u�K�"_��"H�S�
<c42*Z"���\�v��w��[I�fg������6 m\�MT�o���D��t�l4Cu�2S��F@���x�%�?!�/)�_Q �W9мf��9,���´�!�`�^Ak�3.�+�Q��z�F�<D�o6��Ǿ����}�H�[��������`�#RF�5�I�a�2o�3r�`ЁpS09�5��#�jdb��z��?�\y����B�'r{�e�� 3?\�
�j�sO�lp��r�G���3��)��ko<�p_ӫ����Y�(��*+sT'��1�\+�!�Im&�-�Y5����#�T�"��Nř,�gO�B����͟��yd�@!�=&�P�z��-a�Ⱊc?�f��V�fj�s�$��*�nO/���b#7���v�e�Vefy	ͥXg��[}�#�_���̕��g-4�Vg��O�]�5��`�|��d��Sl�ا�Z:�8'u� jF����١� H<�3�ECwHI��vfl,�u�$�&�4R��JN�R�_���fԜ<�����L����S4ÿ������{��.k��Ԫ��[�{�1����.�׵�ؿ�.P��Ss���3�R�Qwߔ`�����א��I�̸�V'%u)A�\�:����2�x&)w���x����AAX���e�"�Oo�d��Iu"��:Í�Y�}F���n��k#��!I��.�����Z�Pc���Z	����s�N��/|\���E1���i�g1�����B��,��A�Ljj1L��u��x��]w>��?6��^o����"�Ʀ+��5��]��� ��+��ki��JD"�m��y=:.����>�d.���z.&@'�3^p�SH���JbD�c�Eo��T�Rw{LW�h��3�9��Ű� L�kr|n�tm ;t
-q�cpmG9� )���F�Y�:�!��f�V�΍Qy�C[��� �߇��y�2�>��8��k�a���5Z�_����l� ����.Ff�qI��U����3������|e�O��D���$��%'L1B�r�3$L4��书�0�����9� �&m��� 1��4+f�Ix1�(�z�_K�w�0B'�>��~�Wm�<A�"�������n����{�4�.E3(�vd�O��JZ+����^���w��,�9�ƞ� /�O���0l��	hۼ>��G��b�P)jC�7=m���#z�( �r*^mŘ]��Z2�^�g:q7����aߨU~���޸[ ����W�v��:V~R�MƀI~��د6�#g���=���Ci�4 �`���r
E�%���������a��(�l#��*v���3B�����U�� �ʀ��j�s��o1Ө���H$��$,L�fZ���N���+]gj2Rƭz֭l�v�iD�IoLR��;�6�|�=�1x0�/�?ش
{��D&����R�ԯ�#��<(:�s�M O��.j���k'�M��9�!a�Yhg���!YT4&Z�"��^^ۧ�
;e6.w�i�r����hJFh#�.�*��
s�o<8���[ê�O�-LXh��	`�](|2�?yZ;�ra@_�~#Y�$�M�ъ��Xң1�>)�$V�o����v�M:�����2����"��4X��ڽ�	҆�Ɉp�ՠv|3'ǉT��f�GVUf�o ��g�08�n���$�P8*O�����RT2|�D�:����FQ!�k������<�y̱��c�������/�N��E��C〙���p<]���������S��PaQ׭j��8x��x`�8�6Wɜ��h?�7��u�Ǜg^$�գn�bEy�綿+s�iP�T�K,�TYO�.���LV��0��nC�� g��7���4���i󹐆4�����J��,�v?'U^x���m~��8�T��$��)�扠 X����"�D�0�Z���dV8��f	�FYnq̭H�݈�
nYS���^��S�	6��mD�,�5������5
ũ5�������u,�������m;�{�Z�n��ҩ�Є�X$�j�㥊~2��Tu��Y�t8g�ԫ{��!LaP���[�	5�.%{�#��vl�ۮ�i xW彷�e�����:Ea���5���j^)��anDXї�ƩL{���J(T=W�{auD0+�3�%i-J$��7JOܞ��!$

����m9�g���ۂ�ӸOg'?p���7-���a���#[��偭�yx�zk
Cj�N�[�:ۯxN^��T�L ��y����K� Z�;�Y��\���o�"�ަD�^�t��>�����;R�/�[�����#.�W�-���"��j����m�i�_(�hn�G-~�kC#%���7%.%e埲���h0Ҭ��3�I�p7˨���.��3<��lg��p͙��>9�$��bf�Z�r�Y�q��̶��E&���uS�������:Ps1�W{�{����}���ڨ�ĴZ$�C�/�;��ǖ�E�Tm0}�-N4��_��Y�KKl��1kBK�����zy�?T:cV�-[E��_�WT�?��4�!���m%���6"��0���Q 0�,�HF������Dx{@?�Mmy����b����ze��YRyp�~��L]�m��=���nlʀxjîj� �G��إm0q��Wr����2���(����Nب���RZ�QھOR?�'���s�Q�x�������S�EQ�s'���vޥ��q���V�xԹ�D�1��O��1T���|�ה%��0 x�q��=��.��mÕ|�� ���а[�*fd;x����S��w���{X��]F�"g���f�mO��ٸD0��JP
��`�������iq�c ��Z6����p��Nlц��e�`if
a��̥B�!�	zG��Y�ڤ9��_��C�
AD�33`�I��)�7	3
�U�oG�]����O�P�>캣1�& �'*o6VH���nC�(­��#q,u�C���O���*V����!�n�Q�&󝵌�;�������m�~ۣ�#fn`{��YB~.m��X�
������|W�W�0O��P��)��]Ek+�)�@��i���w���;U�Z�hb$����r-��ǁ3�׸پUX�.����i�4"�¡���L���z�J�;�I_��'�26P�,8�,� g`,�������J�%�֏U4j�E��+���;ɋ�#���充t��/�����G�y!���u�NwӪ�J ���� -���.E�ƞy(�#�m͞���vAac��c�=!-V�F�v�;E�M^&f�h��˜"�������\�����p�����fK�4�]���0�c,Ff�mJ��v7@D����v�����eB�g�{OnV;N���%���%"\&�"��zL@�r�]@�.n_ԗ�o��!J)�����P��+�j,�0c�q%T����mQ;*�ȡ}x u�[����1#9����?<k�̦ɶ� }�p�����+[W��:��N@h.,��K<��-sN��ש�lH,��?��
�c���On�e��&�;���#Y'| �v�D0%�GJ���G7yCc2���_;f��6�S�Z���58�j	7�jm�!���Q!};�����ҭ}��\(���t�_B
@\@Ks$[�ܳV�?��=<{��k��:P��v�l�*˂��P*z��܅��E�0J�.������K��2������jRuB�\���[9ԛ�NV'��l����,��q���&F��ڌӦ����8���5���LA���zJ*��R%阀��+�.u�B֫��#pO������ď`ɔ�)AY{i6ӣb�	��3���+���� ��1[*�̴q�+=��Y$��HK~�j�X�	g���46b�3�&��/���
U ���>�F��V]��o?�o#ǀ@F?�м}�c$���4:�nXF~��ۮ\��2"��J���g�;�.�����b��-$��=��o7��桐�>A��%$����P��l��%ֻFb����R���b&�������r��n�X��O�HH/u'�����l�����تyQME�c׎��L`YSUu]1���_�����!6�Z����+X��՝4
��$���v���sHl��;�\3"z���v�.�)�����
̦�\M��r����z+�&/�n떠دڳ�A�,/�/`����]�??Q�)�䒨��kf#2�V�,���+g<�>IvL�'�i���0sP4�N�bq�Xsji~;���|�#�]/9�y����_���m��j*(��$�U�b~��ꦠ�o]I]f����̓LW,�r�%|Ӎ ́V��,(e1n7_�@J�����c�'���U����U,��Ĝ�=4�Gd���u �y�!2a�+�����~7�)�ǪǱ��;հ4�G�U7y�ȥ����"E���Q���J9IX�Ou�-_�=���ѥ�ҍp�7�;�T�;y�$��^c*T��F����/�u��e�&;7�L��Ol{���D(�y�=4�$b��q�w���' �_�'6κJ��d`��$8T�~/<�t%����9���e��%����H^�O�T㷘`B�;-��>�i����Z
� ��o�ar�6�1��bKI�JZ\b���g�Nb��N�GYs�����w=�ָ��8\�uC��!nJ��W�,����P�{6�X�b,+.Zڊ�U�������O泅1�i��*��L��9� ���K���=���e J	��ـ�03�L���,KcS?�^�%uey�&�C:��ʝ�ZtjʘT/�\~$��(^���T�4�m�?p)e�pK��S������	�Ӯ'wM-�-��E�������k�VC�_܋����15�-ScN6 /hD�Ƶ�]���]�6�}�{e8���Q��G<G�!`�7y ��~�����|�3+�@��\'�jL��xW�t;�����Z�n�Vc����n�D��KVa͒��$#78H��Vv:���NF� �-rĖ{�ߛ�:�r���,�g��A����v>�1V0����Mv�|Q�#|�$�~�r�k�Y�/ ��P�-��s� _�d?s{�XD(�a����e���Im�.�c�=�#|<��S0.�<����y�&:r)M��l�����5>b��3�4Y�{�� "ik|��>�����*�T � �{��� G� �9j�����3�!gkgc}W;~�H8BČ�sdޡV��/sPwf�g���H^Ц{�Fx��)�DԸZ�}��Eפh_��J��'$:q���}uz�9�Ƽ�@M��Ѭ|K���Y�r��ĩ#D�wX�꺲�@�困�Av`�xC����)���e�5�^�"���+ч�:?�t�Tn��\���׾�gd�"D.-��췇��W�>32+u||��x����O5Q����c�m��v%�gk��J�ν#��p%D�h��g��i���z�x��ƛ�Ë�2���
U�Ɗ��:��L�ILKZ�?]`��	� R�G����#(Z�f�܊9;����/�Q�U��"@��W��'�e�}@K�j�?��U|t�>��׹X��(��:����SP�Fq�t�ئNY�������D�f��,���e��,�YPD���鐜u�[ p�:}ێ?�ߠ���嶠;��3�)�a������5�0�}Ѡ��BM#S�d�c �;4G%�F+0�A�o��	O���A���^j�515���j^1#�n���}�ї���`JN̿m)������Ok �Z����O)����8;�� 4?����(�M����{�Q��UԤY�bm���<����[��^8�1F��T��ɑ���ˠs@���� q!��&
e1���^J�G��Ar[*G
[�0m���U�ҥQ�TBu� ]έ证vE�	L�i�� ��Y��5R��X}w�{�L�������L���nPD���5��)4t�9���h�'WzCB :��T��ѕYn����(�ɉ�	k�:�c�)�
��@��x� y���ɍ�]�*�>�G[�Gʻ�m�oo�J�/�ݸ�~]�k4ޱ�W6��G&��|:
y�Z�E�������)C�� @���b t��G�@ڀu0�S7=*epوJ�	�Hl��*�3�,#`(A*ʋ7�u\n��g�R 4�Q��ũ���8����b#���Z���GN$/�s��U�?�%_l�,��h�>}҂�p��v��N�ӿDb�����t�9���;,xD���ͮ��_��b^`.�ɚ�0�1%@��X(8{>S����7,����76��[��M:�IYO.��P�E��Gr�t��,7�
�M��)|����P��P��h�gq��7j;m��)RJ��Ҁ��������d{���R�EB�5:d��_���Sw/�o~��ujy�&\ȯ,F�K�R��hԲ!ˁ9�1�,>m���\gç5آUx7�^j� uI��q�4Px��4$����_b�ukAk?7b^ [�'���Չ���0���CU�S�h�>�tf�D҂b���e�h 0m-9)8��눛��?l����>��*8?Z� ���-��� �P���k����{���Fz*��q�iF�q������u)�I~I#A$��h�"������:�Q�r!mu�G1b���IuY�������v6�E��P���s�����ư�<�����l��#f���~���7��xz`a1؎WV�L��|PN^/�'�8��KS�Es:,w�c���4�%Չx��ݑ[���g!��ֹCU��j�2?�~���l����P\2�M��1ܫ�"�K�(/P��Ɯ̃���\����3�p���ĕצ���(�o�h
��|��#�2hH��F��m��*`�]l�{X�<���)�f��U�8���D���Ul�`:�����o�ߣ�uQF����uUz")(D׬mP�>T���6l�h��zHA�����SԢ�_���M-�cA=V�퇓8����dn3���b��Z-YѠ�����i�B0���Q����h��ҁ[O>kE-���9%�!D��yco��8{����d,��C��m.�$P���{�Xѱ�f�I�<J��;wOZWp9H9�����}��ѭ,O'�����s���jM
=u�����M_7��;��x�d�u��q��	���P-1u}H�2�Da�C���3l7��L.jz2[����@�u��D��"�J(�s�[��!��Ru:�|�U�*o|���i!3"��{�2�f��b�:��32ژUi�bPs��ʋ�4�|q�nb�_�m/�_�P@qJ�(��;	p�o/�B�������MU����(�I�x+
��pꁕq(��?�:fd´�ϻ��8F������4`]�@�5�~�ܳ��<$��<��ki��<���1�;]���$ұ�!����7X�������3	Z����ٞ�Y;��B���A��Z�Y� ,HU�8��c D��(�c���_�[�&uqr'2�j�%=����O)*���|�D��e{�\/�Y??�J�[���E{�Vf�N���z�T�i�(i���Z�a���ZV]� �+ui���#��j��gq]=����	4Ry����@j6E��ٽ)nK����{n��P�� @m�q�Yk73�(��8U:��aJ#�W��S�C��{�X�w���<�\au]�Z�8fwO���#�'���IxO�"��q�Z�6�g�`��`q�9�(F�?#3�o
D 	�>��1�����0��V��>�bR����gy�͍θ̵�/�_���[Bu���,V�dA��vp�\��~�OG�	�ր��S�mw�
��s�p,ZL�@�Z� �����:~�X#��VdA�g�0h����T��䋫��6�s܂�����I��G�I9XA����*�����K�vR?�۟�� �[g�<��ZQ�����!��6�2�q���k����i2�s�hG'y��(�N���J}�K��sU�n��]'��Y��ManB	-����Vv�2M���m�T�:��]c6ԑ�*!�>$F��6�Y1����2	9t:��a�U���`����B�=?T�/^�-j�W�:[Oz�	*��5>p���_��!���q]�#k�S�XӋ>��h`�-��#�����.b;m�
i���%2��6O�4�9I.�H3�˸��+X{kB��c�~6Zy��|����r('h��i.Q(3�t�\�Z�zً}-�w�(��Z��
���
�;P���w<�,V��!�(���["��?X��r'uĴ�$;xg�Hr������q\�L�M���Y+fo%�1<��L�y��"��j*�����[�`$���8p����65'-ܡh��(���I���
m�w�隨/M����!��N� E ����2P�����D��a�gm��F������&��V0����|�� �i/i���wT\�����^��R�ٷ��wfaV>�[��\�#��<��,᯽�0��H�[/�R���7��&B����@oXϷ#�{حW;HF\C%��X�����d �&|���s!4�D�xT�v����������}�0d%涷"����Lc	�b��R�K(�m 23[Dし"�'e�G�.� ���a:�W�w�dl�T��U�e� ��7��-̻�c��'6�Â	�&��U���O]�B����(SR�;��XP��/b�7�RB�%���0����'Wv������U7�5�}q2$����I,>�EoU8 �=�IA4�c!(�N)ݫ�c�97\�.��/(a o\��z�D�$gktǯl�-��Z���_%gî������&�҇���d��$�(��줢��ۿn9;����v�o4TaNt���?ȹ��"'=P�)&��~�Έ�[po�gנlL���?�XV�b_�Y4*��J���K���Y<d@����WH�/f����n7CY���z!j_z�ze/W��R�_�y�M�=�[ ��w�C���_*A!72�kLR�W-��V�'���lR���%u�T��ۍd|8���\���u�g�>rb\��X�G)�T(����ᡣ����*���X�]j�������zcl�$_���9�i|e��CXC
z
M��ޞ��N�\�.m���4�@g��ns<�k�@��H�z{MlIc��S;�m���E��#���Ҫt�h�g߄�Ӥ�YV�(��"�}W���j�Տ����O͛��sf_��;�X��U$]L�ebU=�@EG6]z@D-<
9�F�וP>m���_hs��c+YU"�t��\�io��]���m�����\������~��/ϻ,�1[(4ӴcD*���>'�9���*�&Y=a����s�!��X0�f�|U��"%�$��Kl�f�ӎ"���ܤ�L�/]ʶ�ge*p�v�Ѹ4s;��G��.=���������P�n�869-� ��i��ڟr�ȧ/�_�qQ�&H��41"�[|@)=6�:��U��)&نfH��m���CЎ�IJ%���@�� �ey��QXV<���ޔ]�h�u��=>��S���<��~�=���V*�����w^���r a�߹���'p�z2���Ä*I���$GW�|����?�Ļo�]ų6	P���O��S�����iA�#*^nU9rj�_���h*5,�z.�=�n�n��F�1Yܛ��N�[ֶ!��P�+s�'�/������P�]�,v��sU&�-��^�9�/��`e�s��"ԯ#��W	Z�766�q�� >��	w�U��A����N 3�׼w����(��'Y$�?ho�J��[Xc��LU�R���:E~����?���#��	�{k��nb��4rk�1@���Z��p��s�[�@���&�>���)Tw�G�qDm��b���JbL7��q��=�A}�$UXP���F��8 't)��x`݋@��c�"�	��*�=Ʌc�C�����u��8봡�;M����^2�!������L�����1��ؾ�^'?�Huٳ5��QBQ�E��qR{�[,��*������a)% ��#e���2&�O���/Br��A�`�ˆ?��tad�p���>��0bc�\3mE���)��"u�y���0V�~�v�y�4�(���(�ז�j]k��5��b���-W�Wz��|�Ν&W��� ��@p�((G*�TFRq��A �'�H�����֕�ZÔNښ�
���m��y6IN�-�@>�x�:�[H ���ý�QL����¼W�@�� ��E����4j� Փԍe��
g�Nx��y֠�lN)�]��ݢ��}�V�:2���v�d��E���Y�w���^}%V;6ӄ�G�<�q��!/K���RE����������)��$'��W�1�����*�n�z� f���l`c��U��<�}��w�9F"���i�/�v�(��>�be���3��.��++zi����Z^F�Y~�
tS?@Pv+gF�5>�y)EEG�/'(ˋw<5�%R���7gN)��[6"~bvv���!c�y���U,�v[��*\�'.�� -,�]�ߜ������5�������LC16#�S���j���7�G��z��j:�n����W"
wEdU�R%�՘悮�]J���E2�z�h�=<�	��g𧫭�����CUV<�Z���A�S��y���f�T.��o,�l7	��k�,��6%
���zsqh��Y�y��si��	/tRn��b���"ɫ|�[b�y�S&k� H�����	��:F��9�,r�1)5/~����k�Ū�UK�Dy�� �f����o�(u���.�'��;�4��ZuJ��L��_$|��c�E�#]
t���:��	=#�t��'�f-���x�2�ߍ�\��_@V�5��Ts3�?νy��>y��j��?F��Q�?��q�1ŵ����Xô�5��j���n�P�H�MD���
��L����G�3��{9��d"��Θ0�Ax�M�D��~�����i{����{����"�-�O�+��AT�b��ffױ/�v�aoߺ<o��omպ�n�Ay� ��h�gc�\�܈-� �,@�!�ݒ����C�䟒|.�T�i���ư ��쌅�;�A��J�]?.�Rw!��#u5�,%jì
%�_n�B('u���&�<*�Xe2'��|uX���@��EGt���9\�ֶ��$|�|��JW��>G�u��^��y�?s�l^��U���ڇ�kZ�>!�,�w��Ӊ(���ㅆN��	�~�	w��$T>~���c�̴M��|6��=�ƻͣ�F��U�����,�	25�D�mLag��#: ��Oa�l˾km��h�Y VF�'4�?I�R�]:��q~���)���P��/�l�Z�!�g�X�bdb��~	÷|����S�T)��=,�;}(���]>��ą`�AD��D��zOX���V�)�7�������Z�m�i�*��0Ԡ���W��f�b *�-���vD;�5��Z��T�Ul]r�����o�/���x�Ix��z�U|����V��>�%�e�eR���> �:����ӧ���% ,��נ�q��v١�b�~����z���;Z�e嶶	�����r^��8Tܲ�)<�LUOV�D�_LOy�z��LY�s:���ˠ)R�u�]ӌ�&TDs�KN�;�;��"��=���7c��e(�O!�h�(�kgi����R��l�l6���f3$��u�g8G}pK?P�ݍ�����Yzk����OV�FO	#/�ݴ��n�SB������	�x&�'���\o�*ӛ���W�D�l�4��@>��jSQh�QrM'n汛��d�arH��V�M�m�y�X�4�9*91S`���t-5i�})@�<i-a{E(�5n� ���0L"�E���r�:M"��U�*/�o��h޸�B��dz]-�[�pIk#'ۈ����W)�;h>0����M0��]U>5h�?4\%!K�Qs�a h�	��2nq���T�Ʌs|�W��v��%�Y{,J���G�L�����^��Q5�z��������_6̦s��n�-�O�k����l��
'�~.m/�Xg�a��!>�55F�o����ݨ��t�#�;9
Ȣ.u2\��c_d@��<������� ��I%�y���-'�"�v��j�pa���'����[��V0�d�ەq4J7e{���i
�c����@퀡'�B�����x�w�qr�K��q��k�����Rǿ�pƩ�J��8�R�aF�%�9.�w<��|�N򢎴�|�Y'q0n��	J�aj' J�����tlV���޼3$ෲ��@*f�ˬ���b(D<���n+�9ҒuB��Z8��{9r$�hkSrg4T��I�!,��ۜ����Cse.������ ɬ^����s�����..�t�������o��B��n�����?{������vku�q�m�3����V��$�!�� !�hn����a���ݩԗ��(f�3��T���e�P���b�N�[F8[�x<��Y�����W�w��3��ǽ�s�2�!���aؽ��T��3�Ӗ��Wz�����p�+� fI�qGߘCqN4U3̼b[{M	"�������~���g] :��j/�&;�J`����Ӂ�d)�;�$|LG��V�abm�?sv6��ɵ��2�x��&{_z�T�a�+���5-d
[�/7��`��qW�𹣯%����#î-ԥ�\:`�� =M��
W�Jv-	71A��^���QA2�2�=�^�7��y]�#R�ӻ��d�+FWNҩ�	^�㌭�`�����&��7��)�v����P�<�UO�!��T�"<�s�{��n��6P���=���K%۫W�?����d�G��M�Iןb�O�AS�8�m+t��3v"��O��.��3b�<��	A p)�}k~���s2hT�ӤK �)7-0��ru��O��^��y@r�B�\ke8��,v���C)�/0úY���.�)J'�XW[�ƍ(�D�?�Ւ��|�����tx�[A��ġM�	8��r\�&'��P�#���~z��'`��g���� kw2�X�H⪛�PA�eM7 ���3�����6��TV/5��y3�aȡe�P)�-)B�o��!�����~{�<��h����PY��>�"���[�鸊tާK	�{�ʼ�
��^}8��?p����4��}5xb���N6�i��f�
:��#eS��t�a�|�����=F܄8:f�t�Sڋx�%ӽ�TG�̬�t�pTKWEƪ�%��9��[�vƔO>�b��T�1t���i��cp�w"�Z��M+�%��»iN o��@�84i�D/�{�R�\�чuWI��ͦ>`«AF_>}Ǔ3�jX�HǊ�~�N8+Ȅ��N^���N�*M%)���dW2���;�Ãs��ط�3��l�{�9�p	�)��.����]���f`��D����`U���g/\�����%@ˢvÖN+������2Ń+v&m*���:�b�,���B7��ävIٮ���Jk����{�����g�DD��k׈��R��T��g�q��_F��x+���(1�p�k�P���j�� �v��	���d�+dJ<�4v����֕>J��"h��/�N-έ������Ɖ���S*-��>����B�o�E�Lsp��t��.}VQ�2Qc�^M�w����ߗ�$����� gA�&|��[��BB��mδ��$�n7�dp/b���&jlS&�>Rf� ���Vv�73�Be���,�R{q(�����p��Ai�����ɖXUhl:9?ō/	W><x�������׆
Wm�^�{M+�N�iB����L��z�/[��4�-���ZR�hO�H��8P�;{��?�����I+O�s��tij.����_�$�a:�lCų쉻��,-xL�766��	>BoE�\��OU�!�hD�o���������"d��^��A&�nš�,a�+M����f�9�(��?�2����o�@˅�qT���6 h9e�Y��)�9z�0O4.5�<�5�lپS�>w��ξi�g�7�
�d%&���9�ro�E�*{F��/)�B����G��ڷ�{!f���D��Pd��1��<�]�,7��5�H��+\`TL���"k��$�n���ED  �
�`s�z��+��1%�⅖$t���P\�I�^�G\n_�,6]4��9f�(UpQ�r���:�'� ;e����ó�o�&y۝Bޟ�,�ϩ!ܰf�]�n5�yݠҾ<n$OJ��עWo��m��e�ZaK�u�I�1u��s����8;��wL�&�ף����VG����Lt�(,/T>a�w���uRB�,��pw#A��.���%�"�:�7E
KԭhKwj�4YW)�_�r��?�0���7��Dy�sp�O{�i[�菘ׇ�a@��r��i2��0�1[t��[�>?�Y�L�Y��R�Ec���T�D[Kz+��?A�mq
LE!�Y�eV!g�γ
������X�����w4�?_z �Q�z���}��k���5ʆu�SU��}�4x#�'u���.�e��=Z�������q�v+'���c�g�@�wM1�[��\<,6Xæ�m�/<�c1��������_e�G�b�\��ה%�"�̭��Q}j���?�����:�ﶢ�Ι2w�#{����GT��MG�&T�����=r.M]�D�nh^��q��gej1�%�� c$��m��I���SUl�����ߡ�!��,�Ak���l%)�!h��7�wq�й�A�]}#�EE�����X{�*�a�J�U	�`�)fc!�9V@Q;�>~y���u1���;Ƚ���r�un���<M���P��w�A	*2Q�h.D{rn��\~Kt����Q��l�?4��XE�" ��o��`.��隆��+~�Q	e����(�� ��Mo̴:{>�BݜE��h�v%��pt��Z�p+�jFt��`8/B���i����e��('I@����FfO��e6s��M���B�UG�7�K�.���J�Q��z�Q��y�aI�yx۟�8þQ<*�$Tw���>e�X��v�oh���qvM��d�G'��R-��x�h�$_�VqU�'�d��h��og�9}��F���ܧ�c'������t ������
����'7��`��pܡ�x�R�^"���9]7�y�Uy�L�/���Q"��1A�uV�8ڭ��,���p#`��Wlm>��X�趃�A_�'��F�\A�#W�L��_rF��0X��,��r�G��F\�fM�o�V�֢3�g>�a�7T9'��e�8��З�z-�H��JRV�-��E���#riB��:ٕ3"	
��>z��@F��%ӟ�n,��o)e�u!P��cO��2=�Vk�O��r�/�^��G�#�g�?~�m�	>��B�g�j��G����&��A��D��ᮨ��r �r�|z�L��� �:��g)Ґ�y�gGK#a6$>Jl�~{���.7E���BT��<�53��H���P2�_�gen�Y7BW|�l�=m5	ٍ��I�5��Q[	�bYQ_6(�v'����OBbTi�j�3��ے�)�i��R�s٭|Q)0\�xa��!�pn�X�=Nෟ��aD2��\.`�@���$�)H���J=']DVK��ʂ�1�;W�N5�R>���׾QV����a�?��l5\0���.7��W��I�o����35J�:ocd�U��`{{y#_���+h}�e� ��C��ΰ�	}���c��<yU`ɴ��{ҒE���Nz�3�(vj�0�&�v\?�����iQ��"g$�K��f��R ѝl��kv���5��i���X���$M;��fn�D/B�׌̌���Ji_F��
� gå�$����V�((�>�:�k\{8�� �<��pl��|w�1=�S���g����n��"K����#��Ҷ�I;]��8敓�:P"��hϩ4�p���y���	k����"Hc�>�������:��m���@�N���	iO��,|��wk��w�f*�u��hK��lw� ��b֏�AR=�D�ϮB�C 
�x^�?�«����<�e;���i�Md,$WF[a�R��d�'o�U�p#�l�@K��#k�#�`����:q����^o�kZZF����ڭn�����f��"���FӺ�5�l�-�̂�����0N�-W�G���+/L��9y�~l�`�#F$�,`��6;c�گ
#���7u6E�^���8�^d		VR	��f:ם��)��WF(�	�����Wg��1(wC{Ж�=$h��R���Z�v���6�ľ���-��.8��D��K3(ێN�w����[�X3��s��r����L�U�����kC6F4C��z;Yn\InX�a;�K"��0�+�oS���嵲��5B�
}��Dqs��`���љyBQ�ӭ0�ҡ�t�F�g8��c7��5��π-�;>�${�<��_5��'E��������������j5�4��1�u�����dZ�IN>���]RMp 5��Xn�J<zm�Bk�!�Ǣ|�q���0������;2��A��)U���^��I;�"��?��f<�5�fTS
�<��,q [����fCa�����79���x�@EM\�����˟ۃu��srb;�!@���$^�ByM�x��+��P:�p���yi"�M�B�ܚ,0�$�$�^���VE��1CK�*������O�?�0��ɫ��u���-�W*���2�K��]~�]Q`6�q����c�����eq�\#,_��ֵ�W����E�J,�[�6B�B<-�������%`���
�4������_bYRNM�7�Z�d�V�hŶc�B��">eo��a]����a�T������g��Wsr�\���l�{��R�?�3�$mJ=B���T���"ྏ2e�C�-
��݁y��V�Z�"�X�!ѭ+�8�0+Mv��fnin��V+ˀ�%䔍�j����]�g�3.Au}��.N#�܏W����1E� <����H��Ё:FIu�������'�R�g�%��0����8�G�ux�5V�>��=��m�D�yl���y��b�f��q$H��.��C��L�:a��|>�<��?U�z=��7;�z�jm� 0'��[g��e1$K�Цgl�f��S�@�@��e��ǑS1�9�8eC&��*Ç�;Ѩ�w�+�$�t��"��R��rk=4�8-��kK�F�g{������'p_>��$y���3*�n���^�j��.�8J0���l=!�19�ꞌ�����2FGBД��M������,-�G^�t����D��%]L�L��H��+J��ꌌ��AS�V���H/N-���
݄XY�5��u萓4���@ӑƹϔLI*<��m�D7����^�Z8`�tR�u�>��4�dx�O7=��`��6�A�,J_Mt��t`�;�+�\��p ՞X��$��B����
ܞ����V/�g��Y�JW�W�"^�m�&�h,��	�a��TA+6���{��bi�Ӷ�!��2;�xp�](͇S�l
�DD.�P=��T4��)j�@��tPڅ�o�����E� {�����7��8,M|d,ޥ��(�]�d���0 J�>�S�`Z��ӅH�Z-����ˮ�?:E�C)ҮѤJ����|�$[<��@q�;���J�s��J�A�l�Gw���;�V.HNR� :���$���bk����� X�(S�%�4�'׬Z�3�ݬ���j	;t�9�F�O+d�A�o����+CQmk�W�C��ېU�"�mN��|�N��yiISgmW�?1�pn��F8U�*�'  @0R�Ҋ��>��W�	9xߘWm�=գ�b�J���$Q$g�a�?8�̎�Z,F~-0s��i�t� ,�6��Z��pe�_���v��ظ�:����AU(�\E�8P*�ty�%�&�?���S)�3���\L	��rt�<����b�#!ظ����s"��䆳*?%{*�[�yp�����t>.j^�fv��3Z�dlJ��Ev��	�
�"�5z54~tֻ��3�k��"��PSv�y�@��ٱ�4�;�+f\�'<��Z���;��X.1u�c���h�����B��vTa�sa`��.��EćL�BN��W������f�J�$�Y��
���mT/>�*�7�ZX�	!CjIY�l���)�)�s�w�i�i!�<��顿R�s:�'��r��������㣵��h6�����q8�i����x��J(J(rCk���Ǝ�<=_�ˤ����٦�?\�A�F��+b>%���ݔ����MC^
����6��M"��7fZ��N%�	�U>�/��{<{�sK�;�d⻣G9��{�F��>����z�y<�s�}�a���ۜ�IU��wt���������1tܱ�� '��f����t�3'���y�j5�vT̷}mνN�x�Y��������7|1�A��0�lK�������{�D����]��Ft�ED�tD>BeP����\7�m��l7K���d�����h`Y�d~{(���� ���h2��� j;�Ry
�Pi���4� ����Ð�����´fF�XMj��-@j���[������������~F�Rsm�3�s< B��9�@�1��R"��/��r�^m���h�����(���h�Y�R���M$�&�O���!����:<;�W��/�O�[rYk]��1� �f� ��g�Xϱ���^�M��P�*��C�f]�0V)�iK��%k̥*�1��k���c����H�H�
�w��$=�Į�ȏ��H��J2�!O�:���z��kEx��اCfg�]"TU�{QVU"u9�ZrD�6˵U�jI cR,�;�4�W��17v�X!��Z��xK���%FP��[c�`Mv�r?G"�s����8��N1�e�fu�R��`ى���B� ���l�AQ�wj���[��N[���C�>��y���1��Er�6�H�0T�f�ƪ1�Q0���m������=�m�"����rK=;A3��;�֫�BF[�l��d�mX��t�7�Z+4Tf�/�@&���`,B�aP�*��+Ѻ[e.�ᖴOU�0��x�蕆��i:Q�/�-=I��%cH�X��NP�g�P|[b�i_Ru&5XOP$c�,�If5��d[��U2���H�⿋�RQƦ>�q!C��e3iV�Ñ���?wZ�I3�j���1������b�3 膣�v�K���2.�;���"x%�[R��1چ�
�K�|��v�"�T|!��)�9��.�PK}�Hq[�hy0���B�@C[�׹#����Ě��%<����JO8x&�8�ʅT[⻔��dw��s=�c��C2��#����EU���@d>���ʇZڱo]�{1�u{��܅IgD������XH1@