��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����Mڨ��˳0��`q�M�'���2&��Ȯ�W�4��д��|�6�K!b�'mY�`��L����T#�
��𑑂
��S���&Bp��ǺOޯl���i}$������ǽ���y��=p�i�̪�#p,($ds
��8j�7[5�1��z%�l�K_\)����h�V�v=�4|��cEMF��U����t�c�-�a'n,�n����y�gtO�?E/����4��K���u��`écc���
�E��]�5��`u��?`�q�f��㽄�kc�b�&���A�_��"!S�_IIZ>f�B��:lJ�櫇9ܶ|�e��%(4{�?y��.�Q��YQ�%-��bM(AK,�i��^3�I�cl�Z�4���d�\L�gc�g�E��{��d��6v5\��s�j��L���4���5�h0.gJ����q	P�ݨI�aT�bCv�4�e�V(��I`�_.P@
YՈ�&�L_K�}� =HQ_�&�3���B-K$u��q&�/�Ҁ&r-� w9�z���yV���hw����Q����#��
$�!Hp�C ��N����2��܇%�(R���
?st���1�K[C�[�@t+����wzF��)>"*���=@����7@T}�$�8�6H��8��z.4>�u�w]8��I�����4g��/q���7Aq��,z�Y_,Z>��S/bm�����{��۳�۸N��#c#��
)cM�c@��7�&K��/6�<r��K6
4����%7nIU��6見�Z܆�.�c�p"W ���P���y%�T��w܃�%h�Sk��]jX�,Q�� j��M!j5�i$���{ؕ��ώ~�8�sV�p�X�^��+|���Z�Ҧ����o����E�r�?���O��?�3�֓�GX��,P�2 �2 ��^'ͽ�ʃy�"蠛,�,͑)���,�����,w�4N����-���;���bC�||;O���"N�U�����A��� E�>��0�p�Ă�O��H�4 �9�ܕ�Wg�ib���[(�9#dоDt��.-x�k:vn�Y��R���W�^�sF��|�H�| /�*�o;ò �Am�p���]�.�mS�?�Ҍ:�8O�����:j���\��W2v
vP���������������҂ X�+�GHI5��G�'�|���׼M9��qc�WM��P�(U*b�"+���֢��M&jjJ��!
*�����!�H���?b��f�1/h�[��z>J~�NѰrƜ���c+���Vڵ��f�����;���>~Z-��d:�L�Qs��ޢ�^	Vu�/L��]a�G�rP����i߭��ڊ��X2vǨ��WTC+zOTl3B g�N0��0�q������s�ꀶ�S�E���Gj� Y���2Y8�cƋD���4�Aa�i��l]�G�9c�ܶg/�Vr+�%���*v}���l�w�7z�YP�_D�^��F>�Y�ȳ9�u�=�W�Ԫg3.�:F%[j��yQ�	�E�d�4�ّ�Y�r�ˠ��!���%�Tt�R��U_9�߁�:j���y���a�������؆&T��ءo������W����WGO^M�Ex��<*ж�b/��)gb���A����."O.� ��
n3ױ�E*�9Q�7����<��E�~%`�e�QW�ɫ��jt��B�T�RW+t2�}k�����Ǫ_8��r�v����*�����r�7%:!p�U�1|���В�����~�W�ġ\]l�Y��A���h7�|U��_>�~>�"m���[R}��G�fgޟ�(����5�4>�dA�Z3莐V���
��m���M�t���Y�L��iC0��i���̄6�Nr�!��+/J�bd�@d���N���"���zcy�����{)��x���E���H��k�<����:�v}}�y���g�rY�V�&+G�)���:8jz@V?���rĮ�*�R�7t�{l�,�^�|��ƙ��kV��r�:�����;�@���jp�9�V�YU4]ʎ C�3_��U��2�Sbu����>�'�b9 ^C������R�DP��YFu�:�	�T�<�X��b���	�sT�@G�r}�u�Ґ�����iʪ���W+ޏ�V�D����t��j��@�H��"l1LxG��׻Xq�L���d'�vv��rq���8���+g��-�3�7���́]j�vl;�~UyK>�T�3'�:D(h U�$ԯej�ԏs#��j�v�ڈ9��1�I=ٮ�g�ֿ�<�����qW�*IL�[�P�q/��|_�g�8��3�D%s~a��K���ݑ�K�������ʮ��T[��K�:J�#Sc�:���J����
k�qs�����n����5��������_�(|j	@��0��<Y�b��|��n»�=�RӋ�QL�7����
[P+DWߓ�SQ;��D�a��"�wĭ�����T����ݕUz2R�&T�V�_���t�6��� $L]����sZ������V=���A�'*%�Pp®'^�p���ף�{�l�-V.-{Y���S%�ňn� Y!��2EQ����iԆ���.��b�h�WW�;�#`˱���y���*���|
K���O�y,|M�S�\uڥ��dX��$�6Q�#�����g2�:K�R��{���Y���`�e闺gw��R���
�v0s��J��0p���O��OD:miZm��7V�hF�P0
�U����R�h��ǝ������z�$*��JU�H�k�7vAw�v���lr�󴩱��l�ڄ_�w6���'��{W0T���T�Cį{��(~ޑA�q��_��
Tp!_ѥ!^U�����c��K�OL��֭m<���2>z�2o2���UF�u��Gz�1��ᯕ��w���ߑ�f]���N�%�Q�eѓ)�Ŗ�������#˩]!�������s8���ۮ�t6@�\�Tcr��]��U|j�XQ&�
���!�b�o�H� "�s�4XC�M�j�r����w�̗�/T�����������b�y�����~���i+?Z�bY�_�C&���`�\���O}��r~��iRw�ҧTSg6(�W�V�?4İS��a���}��#E��z*oδ�m3U1u�8�Y�{���JqW^w�_�Ȝ4�;x�V�=h��i;��5�r�_�O������\��!�`۞����	�=A&��yc�e��<S��lV�gcD��P���^AC'�ZR2�dOt�f�R�;�����g�w�GiV廚-Vt&Q��5��Kwl��/G��_6����K����w0��OVq���BJSYAW4��Xe�$�F��Eo�@���NC^�(]\�^I�G��f]�I�=��J�X�(�;��T+"�Z�U��`��d����URT�zCW�/�Ҭ�'��P7����xF�*���z��6�3�?F����n���I������)2����<75��-���Z�"�s����|�z���`A5���v��1�H�։��4�͋*޿�U�`�)$+�Ia�������};GN�"ы9�k�<�9��+,��:E��3JLuf���������VT���*�*�v_f�8�1�W*���Z��p��]�QA~c�1g�ht��g��&SY9m���X��,q}�*�6���~5��~E2l%6���\�8�2 ��[��%$	�}�O����}�{���ֺv/���I� ��o@�[\uD�@יԕK'��:%�túҪd5�ao7���5=��D���F���]$�[.h�@�`��u`���< !� ]�h%�5������
3��J�W,B��r!�M����i�{��N�cl2՛�r�+���[�x�к�)9��)8�P����i&cH��]?�8n�V�SAת��H�hfWU�7������a%ɵ��×p����m(�++��k�Ƅ�e%J��M�_��/��$��<:
�F�h��u!4�=������Ўer�fe� �`7�0T�Wb�����}�KM�����YO��z�n_B�CV�{����Ԣ���`>�;��to�FV�Y i�!��wۅC����|zZt'�"�a�v�h�K���qU��ِ��ք��]�l��~�R��4�� u[oXEIG�X�P�L���fF*3+aP����6`Wp#�]̟����B��1���^�r �I$_���C'5�@qۉ����:�^��}b�+az��������dxȾ(E�7�[���VFgl1��O?�0�~\!�KPRa��^�o`��&�,N$/��J��2@�/�Z�i�+���f�+��@�
M����Ac��,۾|���:���=m����.O���s	�=�<��s��jE<�/.��:�e�H�1�k~��ߔ�Nb���/$�-�S��Gn�X��w��[�A�X��v�E�3HZ�jp֠��p�֊��d�E��&z�` �x��x�B2t�$L��;���Б�X�f��K��\�Gޚ/Sg�YX�C=�nЎ�j��I0g�MB�!��f[�3�Z���;���$�`*k'~�l���""l�g�8����%�^�?�!���<�p�-��AI�b�B���Q��)��e����'�Q�9���[r�׵��	o�i��P���%M�B�2�b�ƥ
y�hw��iԙ�v�f�:q��yv
j3���*9k��dN�d��/�d��?��R�a!��0�N�W
)x�3��trά?���W�v
���5��ɻ��ؒ���H���T�I�R��0��瑾xJ���"ŉ�#N����C������t��PN@Zs���w	�(�j��c�*ٱ��l��������Y��a�@�" �RP_�C}fĥ@Yu$���S��f�͗��v~�i�6�!9�J7��Q��_����Y?�f����g����ԋ�,O�/�shn��T�܈���z�_�l5Z�%m����w��O������*�M�?��_"�{g�w>FB1���L��\88���2�9t[Z��DiԝxpfP'���1k�|:�.
:-���2f�G����P�1�d�e�F�0����9,�&dz�����k�98j�? ���F�W�b��~}? ok~~���L��0�BH=��pC*�ڈ�E1*Bh�y.�������M�2�'��F�ZR�*�ɓQ���{����c_�~J]���C2������,coYX�֛��1y�D�������XP�!�s�0ᵣ����dhɑĵg�L�S`��{	��#[�5O^k�ԕF�4�䢝ڊ+�����XD��:C�m����/�}��o�J�N:=> G��~�u�ˋi��M��y��$|��b�q7���e����j���:di 4KX�BY�y��0�m
�/!c����}[� ���3d{���K�e;ߧ�m��P��2>�ME6t�W?� P�Lt&�LGf��.6^1f����F/��ul��Xvɠ��6y�lı�~���/19L��!�q��Ȍ"�Z��w�:��-P�(��ǡ��[��A�1>œ�*"���
5�kTHv�mYFG��k��{��H�o!~�;v�uk�)2ّy��Y���l�F������`���Ezv;知��5�^~�m��B(�5p�v���i>�@�v]����ԍ,�'+E�L�t�w�!�N
�h�A��w��a(ÿ"CQDnUղӀ���\����$���0��g?�I_��|�G�=LN��
L0�f>���!�gnZH�f�����U!�S��J7kL���tӀ���L1�m�!�,���sɐ����^U�4ΨRu!f����t�`��\�
%�V:	�C;�:@�K*p�'�d)�Aߍv�o��$�c�z�Z�6/J뫳w�tSE�kK�JA�0��=pKY'k�� >�G�5�ـ��A1��#��I�ѯ�\���N�̪����AT0du@HLt1Q�i��	_/V��2�g�(�j�lʯ�H��+k<�?[�N���R�b����_�}~bd�5e1u���)�$tC0Ȫ�]����iWг_F.������{�oK�z܊�m��(!O�[�-7̾�a}t,���>G5�/�{@�^I*�'����*5�6��Y\u�򤜇�����R�7�]Q)v*Tm��_�dN��[$aN��I���B�FE�z��|�ᶹc�)� #�v	q$;f��ğ"4������e�x�M��'�SQ]QA(ql�7Ψ��ܙ�S�A.F�Q/?��%t��`��h󹒺E�X�^	�?�����T�+tv?>㧦a*xxM�E'�f�O�<��DU��?�x�]p��GEӍͤ����bd0~����A��Q����BS�%TkQ�^$VF��M&�۔$I�U��R�Iq:Ȅ��j�&�P����3cV�����;}@�����i\l2�E�'K��J���u71 W#�G��D	���68��v�ܑ���w����T�Z�)�H��AM���D��H�XPݗ��pQ�yX�U;��v��U�p(��ݳ{H!�G�q�F7-9l�}�`d���^��?6�r�'w�y��|���s��{L&ޝ=y��]�ӍT�܉g? ��\�0��Q)�#�Y�Z�d)����5k��5����=�'��a!=0��Ɩ���aP�"��C4B����w��hJ�:���iĮ�[̜Tϒ��@�8o +�B��=� ���\M�H��v-�-xTx��ä��ǯ9K���JS���+A�*]Hbҧ���r�t���a	*�YYs�����'���xu�8��hl��wڠ��[ƆTq1Ӯԧ
ωZ"� l�:��Z�Zw칸�]τK)ELTi!Ӌi�]�$,&�ù�kO����4{/��Є�X�s����sfߥw�~u ��e� Q��QV����V_�n�>A� �y׃�w��I��a�k�=��ыf�c"A:�R�+^�d7�lS5���vG��WS٫�C��r�Q�6�'@���@1��B���ϗ�$k���:T���F*nu�brH";�/�������q�ڊh��_��#бN��1��Jŧ<Yw�qm��|��M����r���7��
m��*��}r�<�@��<��	V�+S�Ӱ��FH8�"!βm��D�3�z�ǫ0ׅ��oR\ʶ5>f}�'۴�ũR0�tϜe�'E���S���� �fſ�[��BOmhs�#Eh˓�{�(U�c�NRڋ��������H[����e�ZO���Oi�S�,�ƪ��~b���l�>)eC*a�$1~;�,�8��+�A�{n