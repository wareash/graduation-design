��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@���$U[H_#�/8�y��,��F��`G�m6f�f�aiI`������tC����dl���=eZ��^�٭����B�FYĸX�G�����݁�]}~�s�cC�_�V?o6���p!��#��9~̢z�x	����M�8�DӅ>q 6��n��  �	���Oi����P�ª�ج�9���Q3��eS�&�ʟ۹����:�V�ۂZ/'m}�Dv�Cf��)B
�n�ݘ�I`���e,����i�����r���+=���%{��V�ݴ����{��L�����3,{���<�@�3��N�0X )b�t��~����=����y��(�l\�m\���?��B�*"Rߎ�R�ʃ��t�6
dw=y`j�2�e��J������^��ò��-ƀ˘��yqXy��1Ȓ��h*�׈��.�T	森�y% \PU�*AH��i����Q��w�YH�#�k:����db�s叢]����8�Q�
���d]�5�h�Vr�(��C�c���¸޽`f���Y���#�:D?��.Ĥ_��5c����D�Q�{\l�M3�r�������
n��b�������6AZ3���r���%���Ly����7?i4p@�tƛW "�o`α����n0��dv�qnh9!��П4��[� k:{��ERS4�ۇ1"5�E:ԄxDL��AFqDu ��b��e���6ϛn�?;$�=_�t�s�RL8��""#�Z=vv|�g�t�嗻CYY���m�n���
����|�E}������aS0"d��*�q��h��a�9��Xy��1uY-6��Af�����F_���Ԩ��|�Ч���_�y��\ g��H(����|�&�D��F���Vv��&Y�kP;T�7چ>�tH�w[���W|��5u�S�p��[
�>���B ��{�t� и~h�j,^@0��Ƙ���(6�ɉw�ި�Q�D�je������g�����M��i F᩶#�q��Nm_��_�4p벓S��K��v;����
�~jg���vD�P���{�g�l"���Y�M�t���;O��K�!R��!��;az�E�BBB���%�_( ��m��b�W���@Ѭ6��R�3Ed�\P��.R�	k�lE�����Ԋ8�(�5��$�j{3�\�zS�ϪK�3(��}���_ �c�J�CJ����CY�z�mZ���S��B�rQ������O�͒��"V��!��8����H^Q�������s�^��H�N
іZ�3�����D��� ��&��t ���9��.���������C���A찺e��z���1?k[�/}|u$}*�҈��m��K��B0^��Y�����b3�T��Ճ��CW���w���@[�[���!r<9k�犑��_ٿ��Ȱ̃ə�&=Fa`�~�Ը�N������U:Jm�^Ow+C�Sq$��o��j ��ĩD
�/mw�ga� �78�;�P�h%������|��>��[.Dp����g���6!�E�׫x�I�{��1�3ū@��F��u��^�_��ݙ�Hws�0�����w�G�w8���N�7?{��xbD%�l�����Ua�"�9�HhH�P��4:�i�P�H&����u�� �
.|0����j�N��c�ꕦg��c*"%VjJ3y��&��l+�,/0�;g�~�m9 �d�&ED�TL�'Z�,�P�z̎`�4����M�� ��*kӴa��H"k�E������L�~I����C{8��Y�"�'��qy����iS������Dg�%@J,f�O�}��qS���U���:<�� l��.�u<D,uIS�����H�ه�$j+� ��^R�-�������d�v4���i����QԱ馷z���ϡ�� eGt��x�e�\�4�XF!^/�u��m���e�"�/�U�w�����atm-�,>a�"X�-NܧZ[Z�J���j����}�h;�'�G�sW�ʖ���6<�!6{;) /�V���M#��ӅF�M���ı)�[�����ˬ�'�^u{yv����t�Bm��l�t �*h�!�cM��N��6��[���B��]��.��
ELJ��v��l�_jV�~�¢��H��n�w��8�V�dy��Ѽ���,�pQ�i(��	�!�h��W�����g%,pq{����!v��ܖU�8/�/������%F;�+�e@�d��#j�6:�&v�<����3I^?�$�!�f�D����.��ab)C;4 �H����H-z��K�m�E0�dACǘpn~�ZW)�p��~0��MʰN�s������[fN��������MD�.}F�X��86���c;7�La2�����zv�w䡵������@��P�ۼ��򗠸�J��ԟ���Yl��3�ԄB��	�����5���
�o8(cL�	8؊�?�I�EuDU�f�*�1�؃OM�������ii
��\;�B����� ��Utyf쇞�|�����o1b��˸2�>��  E:�}b_�K�g:�.���%R:h���W����ƱcT��������u7�Y���h��P�ȥyVp�����=�?M��`�J)�<As�=��|���TЗL�om�ir�o6���rA�1�P�OdM]f�ݓ�F����Ui�W
CP�Z���&�
K���K��B���Y���s� �F�#5�n��n&4v39��t�:;��?J]��D���)�3�y+�PH�?�«�f Kpn
C9�tS۠{s�n5���2���$�� �s+݇�0��C�TNxI>���eB�!oF<_�=e��h�����{���Z�	�R�ѩ"��Gay+�s|{�kH�Ee��=D�(�ۂ�a�{�͔��O�|��#ٷ�]���s����B,����~��-L(�ѫ��׮��M��}�\ֽ}�A"���)����&%!�<�b�[���X~����������<� U�s��$=�-2��D��STJ��j]��WГ�����6�Mm��<"�@O�&��ޝ<��`�h�w�f>Z�@�=pS��W�� bvW��*�4���_F��N�7��}��F�O�R�����˨�ws�+"�ƛXế�҈���kq�N�_�5N�&�iܻF�+��QJ;��T�a�0sY�z�߅GC�\q��W�SLB㹦���)�4��&r���x"��+���Q���Z;n�n�"�)?.����s�}��m^䔬�[�Gυ�72n�Dؕs5Q���mق#4�.��N�z�l�S���1b0�k#�TB�%�!�Y&}6F���K�A���A�]��̪��r�in�+Ju�D翝oJ�ԀkPro���#���!=3�q�ցٺ�
����TǪ�T[�:�N}E[��k�?��bK�D�W:E{�z���Εd�J�^���K�T��N��7"���"S��A>�b߆EI�)׃?�`��~vy"�jr�-��j��W� VḊ�h.	f�L7o��������Sǿ��?\z�7Vۺ�#X�)�Xd/��v�/ �[k�Z*�2K.v��MY>����E��Ļ5��r�+O��U��e�	��nNUbQ��$��fj���ǜ�x����R̓�"�C�*�f��v@�׳�ɋ�xm&0���]}Ox&������Jђw� ��,�]d}�����˔���"@��S�������x�Eʜ�#�槨�f@���r�S�g=_9��@m��5h�9����5�}ޥ��M�&m�]!�"�(��s޾L��gg�B��%���?#��]�΁$r2=��R����M��6�<�����������՛S��l�eX|͖GK{$V�-����3�'�s�Y�Ҋm{��K�p�Β2?�u���G����*����{�4ӫ0Fx�t�1ͫ㍪/@���]͂�X5�j�����t��V���2���2$a[���N�8_?�T��;<e��1@���p����`qr�m���x�pw�ˡ&