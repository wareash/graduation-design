��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@���$U[H_#�/8�y��,��F��`G�m6f�f�aiI`������tC����dl���=eZ��^�٭����B�FYĸX�G�����݁�]}~�s�cC�_ �c��2)�}ma�dظ��v}�b"@@�c�
l�bx���,���M�4A<�r���w�$�S߇��`w���~p�lV8���
��%�4�0Q�Hj������8�Wnwx�5|%�B4|y��<���C�bA��T�N���Ζ�:U���J�::��;��B��O����k�q��Q'�O"�h$ZrgtI���IB�Q��s��P=�=�F��Q�4d�mM���v�#��D����)0 G<��^� �_�\�y(����¬.��	�y�* ���Ob$�}h��@y��y���ѫ��A�".R�]�hڳ��2��}Έ:�g�wQ� ��)��E�w��V9w{cJ�d��(�	0b�9k�X�� mKٺf�רZ�[4D��<0p?���T�4)G��L[7[�4�l+-
X�tv{Z����N�8O��B�埑{�	"�=%����Q�FF��bi@7��J�5V��n��fo��; ���Cn��m�s`%s�*�+u+��p�m�|:��d�%Oʴg�6�A� i��8��tK�K@k�W��'��X�@�0���K?n{ץ4Ej����=��l�=
q̤��+'<�-AOU^uO�����h��E�!A�M�]������w�l��C�h�a+�����?���{��}e��_����9�O�н1���8����J����j�H�R��T��f��ڛ�.}��դe��;rJz~ل!���̽v�Q(����O�i:
I>{��d��Q��r�D~;�������wB� �����AP��rB`�\$�Bg�E��Xzy#0-IA~2���A�K6Q,��z������JX��	�����%ӟ�ݙL�?��f"S���s��w0<�'���⏤+��p�;��]�<;�x�+;��~�J^��?�����Oɂ�r��E�cD�I*|=r�'�K��>[A�/����~����#I0`l/��?J��
M���ee8��]ʒ6$Q�uNK˧v�bp����Y�}a,���v�=�F�O��}����ݧFD���Y67lZ�:���t��
�M8�l|��w�M���Np�c�S�t5���"� 7���X"��qH=�eŸ���T	|Y�Y㧈nO��V��y�䁒E��ѝ�+�	r�=�Zs�=
�
V�c�)8X�2��B�K�x�%�^�M�+|l3����iW��_��_���b���8��f�;��h�*�QSJ���� ��ξ�;��
�dd�eK�|j͍R��L@�-�^��1N28$A�~(�vUydM��)�if��|�����3���i�4��_>I�
���0ܨj��
fǯh�S9lT�4�B.��[Q'U�KzKfʄ�P�ڝ�8����Ng�SۋIS�E��"x��H%ۺ!�x{1�UGN�U����?��8��>@&�S:?J�
��mY��������b��}W�Vjq6|m�tJ5N�(�p��U���ΠL�������SP@P�6�+�,\��L-'���+�&�<�d�ȍq��&������>�:�c��;~n��EtC����p'��R�7�t,Ժ���m6~=�O� Vh�C(�>�LF�`a�e�
' �Jl�R^��d"X7���J��(������\���@���2�ҥ>���4�b����Gܧ�Δ2��*��e��I�a��S���g�ɓ�O��1$�Uͣ��	�Wt44��|8>[6QO�� �;�LU���Z/� ��x���3ŃzfE �����}T�ݿ�S���׏�h�����*Ccc�܈�+uf~��;�����ù�㸫�hC�vB`%w�<T��vI��g]�QIV�/�TS�>�e��,S�/2�R�ayiΕ@�w<j�#;x�=����"q�p���qTPf_!O(r5G
5��j���Q�֒U
��G�}0����p��C�#c�!�A^��⇉�}�K����K��e
��Z�a�~�v�C�&�4�\GU��b�/�^R�N޷:�M մW �n�+��,ɴ�=)k�b����m��'/�4i�w��R'�{�脽��ӕy�$��:�z$����$z�(@�E��M̵�1m���4\���b��D��1���x�� �u��i~m{2B=�)�����ɿǏ����x�E^��qj<ρ;�H���_�$���]s�N��j7��Ȇ��)�G�k�����1��1�
��
�h�L�m�n��ÿL�ot�U�y���q	&�62.����c�!��2�$} `�&�+�(-��Te������W��T�z·��4���DM	����f�\�%��`�k�RF��
���k��n���=��� �9��nǩ���(ȴ�c-젃7 ��	��N���o�l�ȣ�}���D�jz%v�?���:%�_�B&+Mg.�XG�/�o�J�_i�y�����å^�� J���|20���ؼ�.�Y
�����3�=Ŏ�P(��M~�-����4��Tl�ӱ����x�=�����?�u-�!��6+�Vټ07Q׏��{x��O�j��*1���F�y�����=�>�z�DYӆz�E�v��ޠ��v�Y��17����D7������_mjՍu��U���������6l����C���z�O��!벯	Z�����_ʳu���h0��튮�j�����6cC)�P������0���ޡ�O-�xzm���̉�y˽�lS�ǝi�B��=C0��7�_����A��b�
6���
1�a�ԞjWՄܽ�T�PVY� BB�%�S�]$rk5�+�'~��˔�$����9��$C�F���ůV�渞ꐪ�F����֥:�~�B�8/#���V^������g�5,@q���K�N���3irI��NuO�5N�Y+W��ux���<�M�-N�$�J?��������;��q�Z��B������f2C1��%L]|<Dr��"��I��HS���q����Yaa=�?aw�oDb�sТ��gnqQ��u4W��FH֭\�T�i'dޙ)�%Q6�(J���\:�4��`Q��S[�_�e�##Ի�$gD���^/�@�39�	��paS�{$5@�*����z�(E�nx��l��`��2}iIUV;n��KrM���e!�+�׎��o�#Ո�)�����"���Hgy�z<�Uk���yK�$3����릫�(Ud�䮮$����t�[Ke{��Z HO��s���l>���%��ڞ0DZ��~G׿`~#��{��:i?���Ó)�W�_�`#�>��v��缬M[L�A�#Wդ��J�/[�ĥ�xBd���(bRl��-FH,���v-Zhِ,n��?�8M�ǒ��0\��Wx��������fM��Sh��a�=4�-7x�������Y���J0*~0�T��,�"�0�P����x�r^X&0)I6��Å���`�ѦK�`���BhI�!�U'j��md��+�lד��]�3ic&d�]��&P
��Wf��׊^tP0{d̳'BU��XJ:�|1�o���Q��\Z�jJ%z<ZRQ�S�:��	% 2m
�^,LXu�.<��J���EW�Jᙪ�.�/fǨ�A�g��Dn�rTIЭ�kQ@�\�S�g�[�a��XL����V�+_t��-��U�%X�Ϧe�Ibo��z�ǤvW>$��'a��-�6���>��Q��Tv��c�c '��YU;�=�x4T�S��Q�60�
�{�щ$�j�I.1�t�ً{y2�����@A��y��PF\�}tܬ��Qhq�3a��#�7��<ų�]�W��R�y�I,z:@<<��9gKb_:�]VN��Bd®SA��$��A��쥙�o�k9Z	�9G���wB4|��G���Ԟ��w\3�?v�d�o�^�T�͹ߟO����"Y�b.Q�~���3ߧ:�+�q)���J/+A���)ݽ@��y��#�Y���/,w�`�Ƒ���� >�<:�h���UwZ�_����@"/�����/.AE2|���SM�c4�A��%e���A�&Y��2'ws( i`B��#(�P