��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e����d���f{��@����S��>���4{��ת�AO�Q{�����"�\�h��Z��~�!����c~9�&�wd�B-����pLkl;}Km}�v���(>}�>���m�+<����4��0��E*��3��8s�:�,E�LA2�uXp��Ƨ0K���X)���z�Y�E��hbBBvv<Qߩ-(;3Hf�����"��,����7&�.(�x�\��󈣯�<?�����_�b�-���7S����.�勦qG2���!Z�l��s��+2��B^�B�x'�@��,x)Ug���P�_�r��:i3�in,���| 7�����:N��2��aB��@���՞Z.G�᎙G/��`A�e;�`X�^+wa'�����~�ԟ +�������,��
����cL=���oO�J���ͽA�5��`ݖ�����ܬ�k�]霹�FQ�^�(G!�!�-/2sg't��U������tk��=�-���#�3ud7�l��nI�I���~�J�z��f������i���C��e�I}�.�L#U|�	�"�0Dv��|�{YsJ���YMl�l�[�vb��R��w����idI�,:h�a��M�vl0E����ih�u���s���%ժT��2�Fى!�; �Cu{P���v�j�p�3�3&>{7��GK�C�^>4ӳh?�H!cL(G����%{U'1<�o;���A �]�,d[�V����ˡV��_�(���&�J�;4�m�GjL�΁�=��=��o	�����r��ψJ-̎�&��"��O�>��_�iH�j�a$��*
�K��9r/B��_nd9��!�䃂�a����2��FU9d:�4^����a��ǅ��E���Z[��A�Ʉ(�VS����ە���w�*�b��?ڊ+|��	���LKSxQ����|��Yw�9^xc.M}{��*9�riab��R'�~���ڄG��/�� � \B�^���S"�c�5bO��i�0�a[��_���{��'�R�bb<�V��b���GgRo�_��êv�	/�m���A�k��]��Mj:n_̭1���$Ɇ.�N1l�`��S��b����:�j���R���x�$~�
�M��ZMv�1��tPXPSǳ�A/%�����D{�EF�OѰ(A4��4�Ǎ����L���w�}��3P��� �u�K/K��h�o$�%H���e�����B�S�GCP������q%�;6��X���[ũwV��E�M�V�`�4rqYt7	��[�ߙ27&�H�F�J�w�D� d!!F��&	6&�8���i�V D��w���O���O��]fu[J~:�����3	��Ǉr�`c��cȽC�9��+��6[�]�9Hq���t�^�Sd�5 Ѱ���t)�k!k*�P��P��/��,w�z:	�4��v,Zk[���	�7�^�p�\�Yz�a⿭_�4໊<d0�	CT�����f���ܽ^�������Q�� ��Ŵ�u@�� '�~���hF���M�{��ȴ��`��.4hD�>��qU���e9���-�XQ�q�-�3p�*�V������v�tT(�6����U�KF�@�'Ci�^�����
hu� �O<������V�(������	����<��圊"����B�R=oU��˗���LI##�ē �.4�%vBh)��!i�
!�?�|��ξ.F��iB9�[:���t�H�Ÿ�'�54Q�bBT��/�G�)a�j�II��	����
@@6���ձAӳډu�C1.by8��/��b�M�^�W�=O��h�g�gO�&�GkDi�ݪ��W����R���"�DBk�)Y!�of����t���.��%���k�r��ZP�%8i��1ù�{�ZJ"'k���T��#8TE�7>�'�\�����Jo�ijh�t4*�ڸye���Z�����3N��)��%���<�#��T
K5�$n��`X�þ��zEޥ��N��ٞ��_>��g�T	�N�L��?���4(������OPӷKM�r�Y�G�A�i�+�pR	��~"�Sa�)�/�S��E;!���C�ށ��\ :�h�/f�\T��12ay-ۚ���gY��4I�C@�4l�:�k��-h��<X������M����0!Էi9U���/9���e�+r��8���u*��._��7�l���ZFD[��F$��3)��a}��
��l3�(V�Y����Hb���0B	�v-�Ɩ�N?Epٲ��Pap5I��B�F�	n�Y��}L+�v�=��JM��ֳ��80������|�]�"_��o�98��3c��Ղ����(c��d�T)�^3�U�w)�*8g�9�Dw��b��2��s̎P���rf>�m�%��Okd:�w�o<�'̆U�),r��8B���C�Vn�&��Νx��#�Y+��c�����dX�����M���!+0�g�
�}�{��F�a���e�?��v�9VήA���BH]�C���&5��.�������lt`n�{�|O5���@ł��'n3�&���ƃ7N�Ka�ki���<O+���_V$O����uf0~�1=P1?i�K'�C8(s���!C<T��z�.��ɬ����k�v��c���;F�����/�B��RX�&��W���Ett��K�:5��;[�e�&a]�`H��0�*>��Mkr�ς_��j�`�l�4�U������'����N�]KQ��^,�τ�Y��छ:���}���)��)�r\/����gr���n�GS�V�/}%�����v���?a^�4�izQTq#�MҟRZ�9^8�}���F��1s�0~0X���.�E�/�|e"F�U�4��c�XW��O�y�;�H��`�G��q.z�U>o8$��־��Y�p�d>�+(�����@|dT�f�;@��q�O��r�v��K2gQ>��\�ZT��t$�jZ�K݊$���,� )nZm�O3|Q7s�t(/s:0r3�$%��msj�%�_|�f�zԠv�^���殅�3�L&xJD�Q�տG��j��{���Z��OA�
�g)��c�2f����\iW#S�)���)�[�m���;�J�G���5�ŃS�x.�]˂���zc��������½)����#!%3P��_�Q&�������ġzW��s8��Y��c��i�꟬�O���ТfA�~�+��T)lz����U��;�S̈f�~�//��)�����%=���Aۈ�����Ss�F�||�`6�S���4����מXq���	�����/�Ψ���O�����Ȱ�@�!#]��3�Ψ/���_׬�C�Dhq�����O�Y�1�,��g8���1B�������@)8���7�jRdE��hť]5�pf�0�4��cɧM����i�b�?���wi�	�?���������3�7�p�k����R�6��[5ݰ$�:߭�`�$�L�d��(�摗��3�iҽ*�e�VDC�5f�n5O�՘�i0��HM�g9��iw�+��r�<R��=	�����h�5��wꁮr��3��q[~���rD4��\X��o���Z�~���hzKM5�p�\��p�Б����XA�T�4BN�u�e��Ѫ��C�vl�#.`<��K�1�U|�H�B���50jU�_5;J�.�<��]��rdf�V��`���/ j��Ai�^J��#C���{�ήL?t^�{��h1��U �ԗ�:�CЖ�I@��S:���q�6S����|��#��T��[�[(�]#�+IL��r3��p�mn6.���J )3m�>�ۿ���#
77�'�M@�#��g�J����m;��'�:tu��P�&uԢ�Xh�~��������j��檁�czt:�^
����o[�zwօL���h�'7��>�s��f��[��=�Nw�i���6h�L�2�����12�t� �yE�nr^����E���]~��œ�C��}���D�*
�R<|�+��G�V��[��۝q������'b[��;���P�u��}�B����X'��w�U��*�}(ҺG�+9�x?C�o�,tdo�G���w�e�{��U�>!�DgI�Akn��Vtk0�8����ؚ��CD�W�P ��ǭ�-�yr�}��F�G�5�$���m�qI��f�a��%dz�� ����tc~�:���� �0<3#z��S���U�OE6�f�"��qg�֝�����5� ��4+�.�+պ�N�;g�"�wXՠ�B(�������8�e;k�����=�R�Q�r�+��n��q�. 9�+v�I ���Ü�5�,��� $�����s�Ì�.,ހsh�������2�*��:�/�Q^P�7$�����6z�"�<:�E�3G#N��I�;�L+��c}����&)(q�{L�a:��/�)0Qn���|`u�p�|/f��ߒ��Vx�	N�Bӓ1�*oy�d%�%����<i�\^G�6|�ڜ����l2F6,�r�z嵢�� ��2*t��"^)�&ud{ �Uo��p���G��Tw`��>�D�P`�Kt���]\�A�w�����>��ǀvǉ�EE!�Ä�Ѝ�:��]�-oT��kه0y Ȝ��"�$f�2+@�1uN��]�$I��u��)�*F�ާ�,p��ÖG �9Vؕ�H��{X��=6)���nK� �Ox���"0�b���|J�8��(J�����`-�
�l�Mƣ��:T-�n��w��FȜpF�'�)ڮȣ��)K�,K.�M��`���;(,��wn��XN(ب]�l|����H�����#m鄢�N�_`=�d�#}1c�S�c�ِnܾ�I��E�*U����yv~D^��qWI3@��m4��ӧ�peL����e���ZN�F|�����κ6��<P� Kc�ݣ�״}���q��L���4u�H��濉�Ƅ�I:Y�3̖,�����}Y�L���k��~f��#��R���b���Dlv�x'Fg���ݍT���U�D�K$�9ppɁ/�=v�o"�,\����.j�Rv�e���b\����4l�b#d!��dR�8�j������eL���kK����#:�9V��
�&{�J�j�:�FI�裱j�@-�٧<9+�/s�Ԧb����_0d��+g�L�[V���2 �3	�����٩'��@���@z6](rpL��qN�!
RM��f��P�J��TN<e7�t�ņ�:��P���f��$������}�ڱ�$͖�AqaۮPP�����=�K��<Xإ�����КB�Z7���Uc�֣9�q�&h}�CM�W�+\o9�(���)T������p�j�B�V�ll������!�.6L(���B\���*��Z�c]����g�~X��T�ۮ]ٖ:#�8n˾�y��oڒ���6kZ�(Uk%��'��t�a)����V�@��9����_7r���<�f/}���|�*o����f��"؟���Oߕ�>ӗ�eT���n����\� ��Y�lM�$���&�K��|P�rL�&w	D+�'�����yx�ô[]�-�1�$��v�\�-څ��̠�`����0�p�zQg;��.m�7��Z��\畈س�A+{j�62�ܲ�7�N �`>���ʒ���lf����Nu-}���`k�o�+�����u�A�٩��	�����;BŹv�O�O@B@H�ޮ"��R�G�T�qF��۬�]���5��vJ�.W36Eb�����ʏ�L���9C �O���^������g���� O��j��<Ẏ�u��	���[��+��#T5��e:@D�j����<�w��z#�n�7�z	�2��|8�$Җq_�,|�C���*'ő4Y��h��-&"�B�K�N�s.hy�[Q� ���N@b�t��q~��-��L%.�.�G��!���9*�3�?Ps�����㬘�=�Y5n��Ի���5�����B"iv(��o�����2��y����y��}h��������_� 1�����|� ���g|�/6��j��x�֩�-Ú/W��w;SS�d����´���!��k�N�U����F��g7���8W��9�:����Gv>�kr�}M�9��A��FQm�ʲ�7��'��"����탬/�����J�y|\�e������Ǆ�F�U�!�"f�+n5ĠQ��'���v���8�)�.^��*E
 3ς��H#��fM\n%/^$�9 �i7����l��`{�����Q��U��o��Kw�����H�v��g�R��b\�e1��P����vS�bO��-
S�4�I@�Z��f�KmπjC��,�|���LPe��Ը�5����[f�Q����|S� �Ӹ���3���87A�����5����k/[:Ǚ�������{H�
-�`��O\}F�x�L�cԜ�w������Y���i:�{��j��j�'��ꐟNO62�c�4K�q�}Vh�5���p]8EL��� ��_��b;5$���wF�flwR�[�7m���Tb��aؾ�쨪��I+S����k9��&��؛W�2<��2�=��Bw�+���g��_���٠6��n�)������lMp�y
X����{�����+���� |}�b&�.�?,ݙ��j��	_�H�6�����J��,Rq2D�sd���>�A�O'��
B6�v��-:�������
[=���ҤW���3�:4�n��=�|��w�O9��wjRZ����(����HsD(�*��pQX��
鼽/7ɦf��C�W��b��٘S�F��i����	���~s{��0��Կ�S���LY��e������CKc!�Bw�hj$��I=F?F�6ٓ�D#���͇9\y�\�2&���4T��Y8����/l�WٴbF��9��F��������&v`E��\�#c�K.8���o�
��g�X���)7�<k�`�#YYښ݃���1���n���~����O�D��980���U�ȱ�_ʨ�&<�-|���k1X.�$V��-e�,���ݩ� 3Ye��p ������^N�V,='����!��67;���6�P�{��Qd�b�l��6f�	�s��g�`��R(��%p���++�r�œ��w<ĥ�nө{���V��`�w3��34Q�6bf��-��f�[���4�H���fRZS�-�۪o[�h�5�Ӥ�hQ��"�uc�6�U@��E�7�d��ûb@\%]ʻ�0k9�ȁzw�,$��l�zM�������ٵ�� ڌ�*���Z�@o�Q�J?��<�i�=�'��+���=~�����K�� *��ɸ3[���4J�"N-�١/�����yd�f�
V�:��2ˆ�x�_��`�"~F|�ZJ�x\�?E���G_�Dv ��~\���	�+K�� �<��Sē�祂rVp�k��w�|�8
��F43cj���ڕwu^�	���V��n��lot��rϡH)p�VvLN*G/\Ԁ�n�����Xv���	 �4�Wx���᭲��LX����.�f�(�n/���*P�S6��F�=m����ͫf��r;�שR�?��x�ADfN����c�����Fk+��a��%�#;��,�'&[����'�����J`�-0�,9��M�5����du�j�����������E�t7�$&r'���QTb<�o�G��L�"������}e��C��5A�Y��^z��Ph>�D�!���G���w�s�%k�B 5����UR�uy�g9B.f�F���a/OpR-�'��7����(�P�j�֮��rf]LZܶ�)��T�ӧ�	�Ȼ��Q��6Q?mqD�0¯�ٕ�EnxŠS���U{���x;8��Tsz��3-��$`�O���2�D�tF��#�D-��ŝ�� ��1���;������<Y�)�n+l�uZ
%z麁��D��AXu�Ie�e����k-kr+>���$V^)dߍ��5��jB�s�X��;�	�51ΰ�K��=j0=w����&]|���B����6%Y�%O�t�H[�?�+{b�Bۢ�y�!K���ExP�oBXd�Cz(���G���Q�����M�ɝ�4��P���A�̙�=��&�p�d��zb9�/�����Ù�e��YW�z� �Y��b\_OW �p���;���xR����x�e̚���:<��]o�	�J}n��`+ ?
���h�ٍf���\�o���L	c��$��U��/�-�9�t�G�{��'IF�F]�v��e[�I17<L)G����m��ǚ��eT�{��	j �q!;;ێҳ�m������֓7���Uʥヘ��)�.��n>����M6ލ�wL�L�	�ùK�b&[��f�hF�
��/��. w�ܻ����I^y����S�I�ߎY�VK27Y���*̴uU|7p�3v��7�6���ICt.q��_����
�Tc�!���o��	��<�zaZ�*�������c͌/��t9��x��Tyj���%���:"�=���B�>�\���hX�7����@���v{��΄�Yxj��+�{��/'9Rz{�ލO#�u7�2�Syj�:�L�}��Q�A��VW�����s����]掱����� -�O>�˯�D�v���nC�8�9��qKuT�%�%�A��2q���s���|+��'SoX)����&���4FaN	v�*h�qn[�6�=�ѐ���ڭ����I��6M������X��FJs\WW΄y���<�-���A�u�_}[:�֐ (�/�a$A"��=�3��?55//���2˔v	pF�z�����_�m���_��]!�O@�#j�$���Ua��#]REמ��?�p�2;\4�U% ^��1�lJ��>o51g��H�OZE_d�(3j�ۥ\1G~(s�d���_�X<� ]S����$Ĵ���҉���r�`�yzdudu_1�ja�$�p���ↁ�d!��6
N���wIM(ux�tJ���Q�~+�`�\f4[	|$�.q��F�ŕ�޴�C�W��X�h 4q,a�v�"�>�9����X�نk�~y�D��N�g��}�a�Z�������Q�DKƉ��qk�pՒ�@*i�u���D�����B�m�;�<g�:㟴�pj�0YA5+��L־�S��b3��c��nE��q}�ą���[�gb+����E�e��8ɮ�j��w���_���B"��g�T�s���b�)�G�_��"�����:f�Y������e��@4ߪ,�$~��`9B�.N�����09a�B����Z#���.�K�}���R���(e��q]���ô%3���?H/.�(�{�JU�Cu�w�_6�T0pb�)�9����N
�w�u �⵪+z�Z�-�a��u��';�r�oD�!É~�j8�WX�ha7�љE�E�����Kby� -^�r�U2�E3�B��W���f�S1�1$iB�u�w�U0�:�����yn#��\<��a��/]�a��٧֔ܛ�[FP���*d���T�q��"��l2�x5�禉���)��n,f���;Ǝ���ض[+�eju!T{Pu�p��F2��葂T
����u����a��	CBTGA�jݢ�k�6M������6SGN_�P���삿݌�s����EDf��i!,L@ i��8���-Bm�I0rI�Θ2��XN���[n^���!.��q�dlJ6p3���CC��n���L3b����}8�)�`�zP�Gs�Ľ`F�q�蕖�-s("�q�TSy���(6����d=�Uף[�&�V-=d��ނ��\+ �d/y_�L���# �]�gЊEf�������/�p$���h��<L�3���<h_ѕ�張v�Eu����'X��C�&XV�:�p�h0�|c��5�W@9 z��"���֫"�q�TK��i�RER�dy�   q�J��{1��Y},�'��0}�_���f�CY'�Dk��~�"J��to�F-1��n��ɸ�Z���wu���Lh�V(�dg/e���6�m����:wҚ����<�Иo�֚������(:B����li�����bYdݑ��]�R�!xe�>��_��$��ό#wgm�� �}�t�j�b��tM�>���������,{�������ƠY�W� 25������3�}_�$�hd.D���ca�cD<C�NY�d��X�[�ߔX�烄	f��$�+b�
�&�ExM{�Ͱ���Ψ:��GP��s�,�M���<��h&}�t#6-x�F�Cf�vȞ�<��E�ۋ�G��7�,����"�-�y�1�=U��;я<�;x�E�w]�8��9���ͭ4ր}R'L).N@�7z1>���40�_���tZ\�\v�����ގ��<��3αX�3�8�=�?Ĝ�0�+���b��1J��W5����+��KH��H����$���&ء� �n,�q�K+*H�Z#�Ku
�w?�`��.�t�d+C�F�K�Xv��5R�[Mݠ{��C�'�|����!�,X��Q=�Bʕ����& �u�9���ێH^��ṵ��WF��+tV���g�d���vp�
]��%�׈��-ˉ��$Bp�����#�i>^��&���$����+��������R�]<����bw�OVk��+�#��4���:�4�Q�<�*v���8�+�eh'+t'v��j�CJ6���,������J��ќ�ar���0�pֲ�E@:ps���)��q� ���m�T���M\ �6dvQy8�^^,��!�銆ɽ�w�y؁�.+�6f� s��: !S��bcޭ�[�d a ��T�����o��U���6CkZ�0O���B>�-�@<[E-��N������W��,�k�.҇1���9a�l�n�~C#Q� H����M���[?qT���
�S+8\R�iϑ՞�R�=�[�E���d���0�[r�k-�����t�Wg�Y�d�q�*�=a.��G���1���KR%s�5�����S�%3���5�T_|����OE�n#�CAh��9U��BO���˄�����n@��wPᘧNmS��n��p��F6RT.�j�EY��/=�G)��z>Ȇ�t������ݲ�$�47�I�$�=T���6@�M�qVnZQ`�/�Fﱱ0xf��F/�u�a�	2OBd���BCii�i���<!�����P7-H�My�\<�Z�M�����?p��Չ'���Vɜ���P)W5����k�]]#d�;9���1~���WJ6�C��u6���[?GǱ�3'����H����-���*�^e�)Z>J�<+�����=���N����ImYO�hmgZ8s~���7⃠�FEuB�7�cP��^�-�bqݺ�Bʣ^�\��D�4���^\Npo��9Sǻ��CbZ:9)P�U�y!j!oȫ�����fr���e�7E?f񑬎�D��g�Iޣ�*G�ں��1��<j�%���tG��x��8c��j����²���;+-ﻢk����W��U�������!J��,�?���<�1�天������K��U�Ų�����֛2�<��.�(�肊�!�W�K]1sk���n�*Nѽ�ĹA8�؁2�ǜ�����Sz]�i��fw�Xv̘D�A�JQ3�΢1s�W|��Si��`x��|w����qUQ���É%#���8�'�XU-èi� v�ێ�,dƗ�e��S>��J
�I��
I�ڢ��t�!@4��O�=L�xK�x6y��g��q�V�5�g��R;��=\U�)���EJ�q�����%���f���d��}��$���|���l�������4V�3x��vV�{<xU
 ���(��Xj����v�h���VP��V���*�����s�ί��峦;ҳ2{��@��gj����+kLI�HZ�w$��h8>$�����H|����ʖM1ie�7f��z�a��[�sL�/��$��L��2P��m�� �l��+Pq?j����־]� n�,�o5P��/xԒ���#&i�$?Ӹ���'O�&FԂ��Jo�ѫ
Ss�Y#7��:�U��7��}O��y�f�{U}�)�|�2�|▖3�yu�A�j<��g<˖�%i>�|�����@���1SV�#���}��?ݾ�+��>��ۜ۹�bD�T9�F	�� ���d�����<�	_�_�����@���У��G:�;�7�/y�句�R��w+�Pf����	�k�@�.S'��t����J���J
�{NX���ӱ��g��w�M���v6ͅ"TX�)��Ƞ�� ��䒩���d�2�x~���5��MU5�u�p������o��oނo�^�B�eq[�`�j�N1�v�D��.3�X�{�U����:�)6%�>o)����<���=��=t�:���m���E�긛g�,�5w�CO���	�nW-�P�h=�f6���*�[	<����	�"��w��KB�ꭧݮ/���'��3��V���J�<~Ja�l�G;��z�\�߷=��\K�S��"($�Di�q�~��0L�'p3R<0
�B�^��񓿑ቐ4�&2��@w�5|\œ֬��_)���Q�Yއډ�N���^C�%�0�K�RYsOB)PT�7�U4q7�P�8�=m"��:���Mr6>j��𴿻�'�#
�s��Km\�Ҳ�i�����nC� �l��g�o�	.��A�KLFmt��(����S��k�@��"-�K'������(M�p7B�}��}G�gw�ҥ}�WZ�����3A
�x�-�SP��4���{����!=��yg�E̛���z��J��ж7}�Ӵ��k��@E��	���I���
�ø}(~v��7�KKTQ�;���,Z�C�wm�q�U��t����S�¡=H��R^�6[�Z�����V�qݚM��Gm���Qτ�Hq�!�.Y�h��Tx���{�Lb�;E=WI�p�=����G�k�!����"��B�x΍]��>�������B	+���ԬI�zz̃����Z.�!!.��}�u��VAP������#��\���1��}�w�̆K7��H�,(dPJ����n�`�ǥ��ldp	䳪S�Ierv~0]���j��C����&Ȕ.c��� ���+��{���������T��ǝ�in���@�~�����\��0��h�н'�]d�*�a�������Ӧm�?2��&P0 ʚ�C�� ����y<ӳ7�C�3�U�৖�M|�\s{�j�Oj�vgop�`x�#��q��ٔ܋M�ɤ�.��l�*���ڼ!K�s"B(޺��6A��냎���մ��G�ؚ�u��chP�y�����-.gf���R�!>���(/����J�&�B��@EKg�����3j�!��i�y=ߏ�<)�=��)3�%�"���8{KAudRd��=}�� ���)�$Be03)��)8�y�r���g�`rǩ׺	���۟iʿ�H3�ҹ76���E����P��i��6�N�Y� �p��n��ZU�%8- ����W����*�x]liq*[��'��֦��^��&�����@ϻ �3cMR����,��yU&\�^�%y���$�~�а?���/�4Z�g�R�F�����6�u���G�@��}���1�C����v�m; N0����>�I�GI^U�|���F.�{n�~��4.����m�1��a&.�ј��p"/_�L� �F25���pp�4�b`�K0fٚ"3��U2�8���q�YJ�b  ������c
�}���+m�]�~/f���\��i�������<Ź�g��|s��ԛ�+��[�t�=�}�jf�>'�5 �H\��j�Q&�b�,)���P��Rr�_ĵ�v�*$��2[�����A�.�+�Y_3�Z�Ev����E١t����7��/s�C�j�b<>kh�ds7{�H����T��6��/���O��iVb�>uf�wp�0ޝ�p��|�eA��.=�K�������?���xwG��7�}�6@���Q���δ�1��hs��Vw➬0�:^u=/��h����F����q���p�35�e�kWH����Q֪.r��0e6��z'@��@��	|��nL�7�FX�7��f������觺0|��{-&y�
!����Qh���+����ͻ�2Kd�<C�������qsg5���VHH���?��N�P���� �WXLȦ���W�W�+�{-��Z¼��W.�m�!N�!��	��Ƞ��r���_�Oj)�P�Ķށ	#>G!U�#��:6M��5�OYW���RCN���nX
	�v'�'�%?�Ý��UC_�O4�׈{mфTd�W7�,���+�Z��a��M`��#��|�ݿ{�n+>�<⽘+M{���U9�,�2g����{0�/(}�|��L�O�*�C��1���eԣ[m�x)m1ub�Ԇ�ND�R,�\1w1��{�f�p��#v"�i�1/�nʮ�� �_83QR8.�S��y�zJE�;O��� >�b(�z��~�W�S�}��5�ۿ� 
|�Z]��ڃ>�e�>��K�_+C�Ϫ�.�lp��
Cgj��_��pv<�qg����[e��`�T�nyx���]�7��Z|.0]ծ�I)�}����{�D��m}�����cr>��v|#�捖�'�`8��B�0�'��ԿF0)�����B�w�Ocp��JM���cM��<%����pB����*�U�� ��$C��֨�I�i�]�u�	�ҭO-a��S��'��G��B		�N��V&x3�2y�e@O.��ꄵ�<�>�Q����a,�4�ZS��I؀��,�zY�-��nCp^�a�B&�o4��[���&�\q�{�@���̚�Y��ǲ�\I��n&���nU�`�a��IؽB�2�\ޑ�ԩhTyl=�C��������_�>�L'N�j�a�'١P�:ZR$n >f�	��6���Q3���$��XIGe�S�@��u���Y��P�I�����N�a���HZ��fKz�!���E?�D�*�Gٲ�u��0T=�A���|%�jF����m���Ko�\���[��v��,8���^iS��J��f����C�?#�"&�1	M�QZY�#/�j��Xp u����ݨ�W���I�{m6'�R������~;�'��Ӊ��l5Ip���!�LE���u�+{��F�.1�[Z&�¤b�@w�v	���q&�����0��Z�*p�A��i�W���O����� qz�����
Ʀ������grli}q���d6�������$�.b�O)Hu+�ռ��Uw���7���m& gU��]SY������;{��DISݓx�j�\ҙ��fF-���4raY������[1�׶�V�z��o�:IH�fp-ڭ\��-�i1�{ω��$M
�lQ�2��O,����/)�#�|��=�Qh���]g�<W�|5���c�-��;F�ժ'�6Z\�@�b߆'�}����6�_5lmBˆ�x�Q|���V���c�S��k%��t�R��<ԙ�3J��tQ��#^"��z��0���	��ٍh%6�'O�hJ|�'Xh�E�MWT@"�������h`A���˿�-�?p�w��m�V(;W��9��g�E�w��&�T������mKQ� �PD��_�^|���s#[�5�.���;8F'i��M� �^���Ao�©��,�uOe�ƞ9����mk��+G�k'�T��=g��w�q8�_/	1C��x�7|\+��	+���q��*:�G�>i+ӐHEv������1"���Α���G��j%لԟ���ׄpuB���u��O]��E�R��x=n��(�y'X=1XaJ��� 9�h����+��,��zH
-��'j`�ik�M�c��.).
��"|%C��bg�a6@�y��ػ�ُ��lC��qR�ģ�z��K���M�?�{�t����#+�t��T �V�b�2n2Hx���C��C�}��Uf���V9���ì�� �j���(a�X;�͠X8�Sv������g}#Q���<I3�h�e~��XX���7����r>��C��@��J������e��l\ڶ��۱v+a��R0�a����6n�	��5!Αͩ�l��������/w���]�YH�Abz�G�_��Ee4�4�<�|���2����D�����g���/�r�ɧ�16�|�0���3cA
��aQL�4�B�}Թ�>A��a�OB���h���1�ȯ�̷fk��*>ܦ����up����I�Пf:��z�����>�1�o�? �:���Ǭ���ü�i���X��d��Ǳ�ŏAs�*��i���*p�{m�1����˔a*2����O�e�_���������� ��ڨ�����R���?>h�}�i`� ��"erg�2���HHf���f�� U��%�~^��Nٺ�7W���,gԲ�w��I��{�<����?O����n-]��d���*�L�:�	��|"R��MdY�r�qt�����׀�0]�36��(���]�G&�/11�v؝����4��C��}��lҸ��K����u�/�����T!��� �}~�.��`ћ��52Vf�ա���%+��P����]�^���ֺ&Y�r�gMq��ȹ�՜�o�ޡW6�}u7�-dq6�TC%B�Z��ۙ����v����u�X�	@��)��" ���h�jm�VL�Fxz�
�M�$P+����%��;�n�߁8Y���p�R]�٠�m�{:� yE��Z%��w������l�{aU�!��LMI'�8?m� i5n�ST�v��9��	.YD���ҡ�c>@Oh���rD,~hƙ��ߪ�V0���
%��o�1��ko��y��� 3����@gn��W"��Y:8�7Z�❐��UEH̢�����ś�0�@�������Wo_}Bb�oͳ*�/�����lQG=��Cv.o�)�޹
s�m�f�{�����X} �m��EF�ƔN�L�TL��u������/���"����]ư���,�CA's^�����c��Ŧ���0!F� �SJJ<�9�pV�0��;����0�*{�6)��h9�,��&__�<T|нŴ�S`=7�0:<���We�Y�Lɣ����0���|T_z�w�yF��C�3$"4�U+��k�%��ǋ�a�s�|р���|�ˠጿ�GͯX�-ɕ�e��'�ދ�ًC��JK����}T��v�H�O?_I�� V�N��~�����Ys�`D���W��=����Et���[-���l(D�J��� ��N�]%��ʳ�ޓ���&il-�C�@1jƚ'���\;]�.�3�)��x�!;��̪��XK����}1��Y����=3��|�8�7�Mx!���Ef�w�:u;	<��pD����*���y��5�Bg^no���G��%�z��^g��;�(������>��O������J�z"
T�]�!5U��5Ϛg���9=9ҥP4�T����}l<2CK�q-��1�~}'P�p����m����C�Z������m��}��&!W��ä�M��r����]p�!��xZ&~�]�~Z�,?���6KaGQ��/AH��z���f�6fBu��C~����J�M��Ga��˱n�xn)H�֬D�t-F�@��p�X���v	�1u������tx/�p��J���F<�M�����j���E��&u8���/Fg�E�)���˚�;S�a'�ڴ��x�Tc,8�m�Qdƛu�;|K�C>�zIoF3�ʫ�Ơ�-&_'�*4H5�-vc�28��ϲ��i���Iz��XH��C����F>zps�_�,h���jx�;K%G)մ�%3���Ϳ��sߘ3��l��v�5D SH�>{���*k��H��WːJ���0R�t���,6A�蘀��N�զ���%���[#Z��G��!���S�)�����O�0G�aTBb ��7Ѥ`3�bq(�b�����t�M�
jAO�7�S� t�ڷ5���8�I	�Vܔc�rl�UZE���)n��V�|-��I�ge>�ϡ��W�* 8{kUsQk�Qz�g�Az͔�sh}�\��݋�=x�9]�`'!�v�����Q@�j����~]>�d����g p��(��s!+?cP�ln���箅�u��wܸ�M�)�����?B�_s���m���RS�;�L�ꥀq�_��k[�%�0nJDd���
L�t���d�GW�b��;*H�j=�ͭ{���e��ç�4ܓ\�[��p����?�W�������f0�Y�� ���Rx;g}���Y��5L���c�O ���
�If��iq���P�n�ۨ�wX��5�o��6�j���i�W��3��7h��Sh(F�.|nad/�7�K7�^���B�Si]�3>������ۢ\+m�I1����G��D�Uf��/�Y6��~��O*�bM�m����yEӵ�Z?<"m��Vt�����8<���қ
��c��'���p�8�Y#�,��7q��찮
�w��x��ǼUl��y�Q���O3�m׀ܶ���������JB�B�ǂ��ܟ]��藷�S��D��A[҂�2W�_�-C��W��}�D����/��v-b�wqC癔o���g:���]�#��I�mf��}�sS|�%p/N� }��=���6����>�<%�&0ї:3��B-'B�?����
��Pb���"V��\�@�K��<Z
Y^wέ(��X���e��ǻV�[�)�
�5�l;��VЏB�Y)��b�� PQ��93{�	�7}r�*��-��Ԩ:Ě
�A0$SN� ���Q�G�4��2�� sY%�Ɨօɒ�Vo>/k<0)����̏�L�f��b��Ns�U������#�U�o��A6[���ʊ��G��S�f��*�%��۱[�ؽg/��>��Jx�p��@®Aр�?������/��̷G��I�y�7�Ǣ3��V��b�˗�SaolĆ�lw0��������#BS��|弎Fɭ��S�x��-�W��[a��TR���ږ�:� �u�݈A@��r��U���ž�[I�E*�l2���]�� 4�#��;��k%d�/CO���6��������7>�7N�� �a_0Qɖ$���[Y��-��t��j��Q��;�W ܯ⩅�]������~���Xcf���5k����u�*?޿���}2�M�PS����Ek��S���.3�{�b-P�����)�Б��> ]'v܆*�����:
��4�}Z��N�P�a
��ȡ;C:�{e���׀��R7\������)Ֆp;L�=��o�aT��㷵d*��]��}?-��%0��
V����T��j�=LTf�̫`90u�T�B�L:�Y� �6�gV���?)P6�f��E)f,���]��\�%cG����eN��K�5������ú;��b����ӱ�D�?��p��L�vT�L	��Σ^,�	�?[N�>�tW+������$ +\@��h��J�ZA��1З�G�>��l�5T��Il���6łzٲY��ʹ�=ԡ�+��^�0�Ʈy@�/�~F�.���x^�;�SK��Q5{o���S����H&�]l������U���N;�w�C��&�0��g��O�Y��¦{�:4���"�C��,��!���0�=�0�; w����j�';?�-��{W���ڋ��ޖS�ѕ����
��hj*��̝��@�ް�+��Az� f��ĉ�i�x���댌l?e�!��c�!V@i�R�G�rz�!Q{��}� bt9���"x��¬4-V��W�[G��k�$��yj�|OIɌ�ȣ�,5�'�#��
vA�$n5y���t�jyt�N;�7�2?<�DxD]�.����^f���iS�{<k!�~-��z�[qi#C��Z�֨�>+RT��M����W�%��~�I�A��Jd>~����6!!Q�5_���Jf͘��!T��ƣ5�-�L�q�\"R���"÷�X�,vW/� c�5�*���D��C@:������%{?�
i'�hX������wR�@k��� �ؐ˔�S�z����@�ⰱm�N���RǱ��������ȹ�h똈e	���v�M1:tc����$�����g��֩M�2$��1q��s�a%�f`+#0���F/���U3UC��bV��#,b��.3�<I�a�w���Z`Y�x�?K!�3����#�닞�=�$t�|G�\}����}1���9��U���֒l.�&̿�z0�n�]ٚN-<!�_v#�g40��x��,>�Ʈz���)��f��/���-;>d%������8�����V4��ݿ�K��Y��W�Z,U��A������$?�p}C7�
<l�Й�`K{��+1�}z�PQe!�%�e Zc &�S7j$n� �>�����J.O)��A��6\ݐ�e [V.z��5��P�gƟ�#�����f&��7ο$;�j�L1��� �`# �L����J�������|�d�-$cT�I�i��o�N�������%-�.EK�����睛A���8v�C�7t��՜=H�8� h��O�|ކ��$���q|7��Q�����*[�L��d��io�\ ����Z�d#����N�,�$���k�lH�gU�eci��i�������P����M^]��>�f�k�����Ju��Z��G��l�hk#�-\1hpr������r�����#��9�O�]�ը��e�����HSg�y��Mk���v՗�no�<b��{�U����~���" gV2����(i�r�'q���٧���OE�Vj��{��s�&l��|^#���@P���ǺQ��Ȅ�M�fx�ig��$c'�BeyW~��p�Ζ���"�/bG���vJ��B��f�zM�
n��Dtr�@!�9X�kb����3������?9ʈ�e�2��V i�]�7��3���8CoV��P=[ϧ�v�����=q�����	(妴`M���"���n�mCcwO5����.�mb3&%����S�������>����g@C�`�8}�ܡ�C��G�擴�o
�%�GE��uD S�O�q�sg���HOub�j�>1��{u_�Ȳ��W�9��y�?�.Uiue��J�wI�6��(Q��ž�����B����㍾/�V�S����5��� �3&����UeZwR\�/J�R_��Iv��Cu4�`#Q}�3zc�I�HSo~�����ZOM%�������׃���~7f3y�hD奍��};J"A@yH�grL�������o9&�u
����� ��ź�뜁���=���8x*L�������r���O{Yr4���0�So���mp�Y'�]ա���usʇO	�_a��暶5�D��*�|/�إ
������8ٌ��(F����2���2�W3*>;������z�Q�g*��W���!����"�mM<�@���O��Z"�Ao��]g��a���ne�#lji��������e�>�Ʒ�1�al,y�K=��*�(1�����㓰�&*{�
^��.���u��u��â-���Kғ"?��:����@6A�/
"�����	��T�z���T�iZm^�PL��G�*2Lk����ODf�Sq�)9+����H�^-��Ъ86�ݛ�7���g�"q����ш_/A1A &����C����2�BDJ��K/�ڬ���w�I�Bb�ʛ�R�zXÜ&���.�oI�}b���	]+!��j�T��s��Bv��"� �prVE��Qۤ������4��P[mr�_0.1_HT�d��JE��������ޞ�%��U�cD������]}�)9�Cٝ@����Ӊ��>�6��:�
��9�U�1|�:c�X����S�'�ե�N��PuiS ��[7��1����<kih���+	Ai���� ���0.3+j2���TQ$�׽!�5��gf������/�T?��s���;:7�P���*���zm�ع��C���/�z�4��|No�Q#��i�3CEv�.��]��}�?��ռ�&�d	�-��!G���^�xҎS.������V�&Y�Б��pc�G�ۙ�SU�Fh��>(\�Q�Wx��~g�+Dh~�pK۪��̼���	gS���vt�I��
+���{���V�E�Ǌ���.�0�����i�s,D���h��	��tD���Q���'��a���k�,4p�F�寈���;�r�i3��I+\A 0Tú��n��Hc�X���p��k��J>���� ��TY��������Z��/K�ẌI��G��m�^4�B���d̯���A�%6�Qu~��G����Vk��O�eυ���5��5�$?2�l�1w��[�A*�j�E��(q�m&n��4��3�����U��/A�b���K�nCљ�7=���r�q��p.X���m�:ļ�qB�L�
ܨ˃��W'31��/A��d[3�P��@�|s��R���7~��f4�9�J���C�ȼ�d���:����RKl�����|��.ޕ �6}�2�]�&��m�ݫ�^��<������g�^c_�R�e��KP�f�D��߰yי�.�-KR꾁���}㑥gbP�1��K��	g��Kvy�W��|�9I���\5+g![(�R���W���|�Ѷ�܉�
I�7��$��KXn�(<�Swy�a���[#a����=��?F$��$����ꧥ�c�4��j$�?�O _/��n��[��1��/M��m����S�P=	H�.:�>Մ����xJ�E�Is��������TV��o�.ѩ&[ ��L�.��XZ���a��.��X�#T̈́&g�qM�-��L3Eo��r�5��h*"��V��*s�a���HqS�-{�Y�`��_�/i0]��CMg�Ö�ܦѽ�x�O!&���L�Fb���CT��z,�_���uW�0�Gc�j{���Ӥ��gG�!χ�]k�C�����9��&�4_� *�̬\3��X�\�%��C� �u�ZI�}�������<�]���w	��}�v���i}�F h�E���Q��$lGCx�c�"�͠�܏��'���<�D���3�lN���D�pI^lr%  ����ύ��Xօ�I�]Yo��z���x^�."�B ,f��)
HUigy����i>��uh�,^U;�p����E�NWN�I�jm�K�}�D�<j`��#�8��f(���
�e�WA�\-y�h�qyP}��O��w�ٳ�t�l�p��iwNX>]����peq��|\_�h
�s���Dqp�Sȩ�d��C�>������s���1q���WZw�,a��d��O-���r���Q���Ф6��\=b%_�J�z���6�Nr����/i��ə��W��΅6Nn�-��6��y�~x�6}�����+��H1����O��}���"cN>kb|�d��ֳ_ė4%c�s7L����E���q�.�4V�,�{��!�E���^����1�&�0C�'����"���oc��dM���WPb�c C#��aYA� q��<Aݰ`6�uS�2	������a��3�2h�y��R7�m&����Řr��}B�P<�p��v����v� J��r�8�Xeӑ�O< C�:d�""Nb\��V��ߊt��~������z�V��A2Eb �Le<ѐ��i���fy�Yy�I� �Bf��wuTӥ!"ݟ�� �^%T��sh�s���!��G���jk7��Zy���^��i
��ND_Kt��h=y\�E�n�����:[����IQ��$?6���T�0��B�5櫼e���T�me����JF����I�q+�#�*IN��ƂMo��]V8#���ަ� �^(��~E]*
�]H��q���ƾ�)T�bNk�����wg���F%��`�����㷤h>K�L�Y��ս�o3�1�wz���z�rWmZCT���Ә��\Q2
5���h�3[�1�6`E�b��G�A}B��oV����4�(�
a>.ؔ�0 !�H�ޑ�OVx��z����A��|B .%;��=�2�Z�l/���:0����Zp���C�����0�	�Zs�L�P2g"dQ�^��#��s�e�1��\���r�w�=�XD�>u�-���D���5}���z��w�O�b��X?�O=�]�nڙ>L���s[��+k0���p�t��z�fFJ����
�L�<Y��'�z�(w�Y��B�G��O�x�2�y#��?���=�-2�'���3o� O݈S�&�ZF�y��~n@n�Q���Īg�\r݌�`����Y�9�sB klzq�j��}�'�3�A3�M�d�%����њs^��ȫ�O�}ze���Y�<���5.M���
9��j�%��P��܊�K^��u�@<FI�� M�^u!� g ������TZi`���h�C��F8y祐�'�{Y�V�!�τ̘ɟ�ΐ���Z�c���?��k�'(�3-��,�E�E�����Ч�W�;V�iR���S�]���[��n�e ��e?c��6ś�6�'0:YѶ�k����Ж�|�b�'�����m#��>z3O���w	��Ɇx&=C��E����k��"�EH����`m�=h���C�[�n��I��pD5��qb�A�����FB�R��������POq����hqU�M^���
�P�6%p ׍�dv,(�xe��C3�a���CFyيR�P�*NUDi�?�d�`��\;�K�$��Xi�d�Ҕ%�w�/�w-��	Ez.sp���q��A@ %���k��-��uu����)�M�^�	9Q�nw_�IZf�Ӗb��S|����h�������bIB���ҟ=�q����i#����M,=�L�t��;�������{Kn ��S��ޡ1�'������D�P��ՋG�P��ӂ�DȞ )Ro^X�H�c���*O��vE�Ȏ���Y�&ڙ�ܪeJ#TK���	��u	/��v2J�o��N��>����K��4/ҝR��}��פ-�1N��D�vfd��p8^�8�J��~=Kh�A�6u���E�ݹ�*N7���Zz�b5V3F{���J��p�'j��oD�_������}��V�o�������:����j��C������k�^�g}a�WMg�2�Xp��"])���kE�A{!���^^d�߷1=4��ce�}(F��������"�f,G]���'U�-��]!��2��[�@3鴓�sr��^��������,(+�������� %�@�S��.L�U�y��0�!�Uʂ�n�+r�������ܲ�i9�ϙT$�A���u[q��DC��"{Fw���^Nħ���6<��U��T�P�-�@8��/�\r���s25 ^P�=��i�}8�#�P��хQkB��9��C}Rp���ls(kI���/F��o �R^�URr���D*���M�6I%�90��#�B��d���ꁙ�2�~��d��+�o���(�Z@SV
��g���.I��_�"���� @�e��@$���k��<�����Q��^�N}�B���cg-���	�O���	V�h��ӿ��dʥ�e�*_�����i"�`d�|U��쳙������t���K��^!���l����j�@�n�s@�6^��7����L�ׂ��e��KkNX��M��mM`{0;�.��Z��!�+���Î�^R4Umk��C6L/�K�g��>7����9ր�������cz�lX�>�$�\'WqŤFs�q�=���m��| ]-83p�v&8F�,r"�g�e�#��;m'�ݳPoJ�Xg�+WΜVlW�	$`�s>r���b�^_�3g�D�I��v��A7/cE���k;�1�(|8^�.�.����LG�?�nպ��G̒�}���[!g��zA
A����d%��n~g��{�[��Z��^,0�y��^��Kr	ݖV[`X���S������f��>�B�9}'�]h?��
��c��0��!����bt�/l��7�XTP/vb���ˮ�I��H^ĵ�^}��uQy*����Y{��Ђ$Ώ�sb���?@���o�Wl��T�9�qV�\#�D�mY�-��;���J��?�{vK֬co l�%+*j��Cb}MQ`/�F���now�5�Ԇ@rU�Q6�/�0!�Q,�]����J;,{Oj�u�Y~�v1�D��\����I����ʘ'9=���nԫ���æ��:r�O�F�QL
斴��-�C��s���5<H�B�	��-?hQ*n��#�f�Բ�鑂�&4�;���,2���SUD��N���0���7�d�ܨzd��3EU]˓��R'Tny���pzRq/[3��>tEB����;Pd�G�e��%
_,�L�6�D�|%��.����Ѻ�C���y<8y	�"#�3�x�g��':�0H��@��/�Kju�a�2���>P:E���T�7 ��ߞ9�7-���' 4��.Y(T�O$-�`�wЯ���ݿ)�[���v��x����ƺݜ8��BC�]8�%��	�!�"o��?z���R���I
�*,Tm��
�-��Q��v�*��5��d���c.��z��,�1�e�-4T�hY���D|�w��F���E�T2�`P�͟]��/��r��Ɔp�U�3�^�(�[n$b8)o�?u~ܰ�v�s(�ND$S�X!PԽ��Ja����º��s�P=m�l�ڻ�z�%P�� ��\�6b�����ѭ�4��Vy���o���E��`R/��2�x�^"�(����S4�rP�Ă�e<�d�	�/�2@u9�tL`��~��ʤ��u�|�9�h)�"d��tj�4��Q�?�D��>�fs$1��ow��Uq���;[���͔]���l���B�OZ��!�1�U`AF��]������u/��y�k��\�����n�1�w�{#d$LDuі����RZK�!^�ꤺ�ڛ��&a���nuq���V
#�	u��ROۈd-m�i�k�5ϋ5L�k�}��w0��s^��\
����a�Z:��dQK!��\���W	�fN]��ly/+���v�<r����!ڏq�R�� �bG(�ǁ���Y���nd�OD�΄U����H���ķTr�<���Bm^Cè��b:%����~�R�2�(Q�{*��rzx�n��5��[�+�=�)8�� 8�N�2�����X�@�թ�����^�A��H���в�.��A9YZ��i�w�A�p����k,3��U���Wd��fV��9P\^�	ƐbUeq���z�J�?�YT-K�"�����)���^��������(�E��mw .�!���œ��o����
�	9�j7IyՏU3�Ϛ����$?"r�'a�r�sg�A���ٵX$�+V�^�kR�#ͬ��|�o(�'�Z�u/;lU
�B�>�C��f�]j����t��_�h��Z&��l/��=����2j����+�v���ީ�?NO.�[yH��4�Ee3Ug�'�a#�PH����,�\`������{���?�!fo����'�Ũ��`�/���^�*�-�\��d뉋�J�o�r+�旯�8vH�_>��V��ES�ʹ\_;���j�C�K��V���l[�	���GN�_ǱN.�Y~wݾ�/q�%�U������8���Jgci�QT�
^��|l��Jd%�dJ/k&����)�8tR&�d��]a1�7�T5bJ\�6!��p�@Gg�iB3я��BrmF��޶8�te`ro��L1;��s��>#{S�8�%�G��Քn�:��hL�����)�q���{�;`�����/fV��G�Th"��'H������[JCY��y�d��Q?0%�Q�d���ں���e?�M(�c��$Kg~�@Jy98��;��"��7�� ��ռ⮜�a+��R@>���+�SC�+�N�3�)�?v���ڔ
Ĉ���1V�!o:h��Z�UU�ړ�A}.���7}�
S�|N)�X�m�\�������E�{����dz�!�̮�ݰ1�㶞��p!�cJ8���a'uο��V��Qg����# �]�MзQ��*�rُ-�F���ﭛ�]E{P�UF��֠�)�?�#�|�EGua��g��-��Q�ρ�y�V�ݒ�u���H�9td�-�5xĂX�^��x�<�?WU���ő�@U\�����B��7���(��
�����+:� œy��tj��bu�bi˭�1&\��D2J�Be[nE�?d���ځ�YU�YB�=���"�O����$.aü|�t��Ǥ�R�� 8��"3���0�1������t�%;�&Ķ�^h$�ԝ��]@�
��x|�"����u�
��I4�|��`��p��8�����~�����qu�jǶ�sܚO*:����<-q���}ʅ.�6S�5��b��|�Z�2(b�Ɵ>�K��O�*[�p`̃/���d��S���B�Hc,I7�2O�CNx�MA-\���+$�+�܈�*�>�e牝�Pq'L��x��U3�1��\���5�]�A��c��%E	ۭQ�����c��nQ{�Z0�}�����6���*�q	tF\��1k8�w��	.��zf�0ʹ�|V�B�g9�.�e�-���[�؛[���ou�
xjd�x���Ii0�����Py�������\6=��|��q��m���l�9ު�� ����9ɍ�d���w曝��LA*�=L�����^�3.w�� 位��pP����̪��؁{��V���8ne+ʭЀqwӂ�l��l���	@�ό:����7���c{��7���Ҍ��em�[[����U��.��.A�֢%��R�P�h�:]���KQB�#����<8ʆ����Ψp+�11RiUL�~Ξ4�}J���};NT �z4/�pr��u�"�CK#�����������q�C�_��Hg���'�t�>%n��I�{�z�,.R���TPlB���YVq�z���J�� ��Kġ����6C~}�Rd�
��>����2���O$a��Dh��x ��6�g�
'"Mm�3.(k�\?�ea����E��X�P��O^�;����i;�ׅ߅��?=K�� ��G���%a�B�w���\}���JBpK&4�{O��|17���A�a���$�\��'�B�4�t.!4�ݱ��T).�n/T�Yv��kh�yt����R���j��R�Y�=Ǿ�K_�����"H�^�<^y���mo����űm�c��\�x��I���"r=A�.�޿��rrV*i;�P_� -�v��hE��ٻ���Q/�ဈ�)#��� R�:#I�yv:�o��BJ��M� �`�u
rr��ͽ��-�R�d���[���J��$�x�1�C}���s5+�8WHr:%��U[�m���
��M��.+z��D{�����Y7�y����"�8L���kb���ߡ��Ȏ]��K��Ft���Z���1 �V�y_ "��*3��<���Ŵ�w`0���F��rT��[к@3�c����R�(f�uud~��*��! ��^����~�����Jb�T�������c�Ss�Za�
����|"::.����Gj�"& ��v`��~	q�Q0�:��M"݈=w(CVd�'��c)`涗���:�I�҆n�A
���j䜙o��T�J�^[xŌ3+6ډL�Ex����%�M��I7�`�|ۿ9�ǧ���; ��ؽ/���v���􏎇7�������"bTQ&�j���s�=$�!������)[�����|͇.cw�tn�`QU�����/:�T�Kl'��X�_�bٹ�u��T<�L{��c�#_�uE�k���o[��JX���ߐK��QC �zl��J�ߊ$)e�1I�W��͔�4R,!�s��=Q�c�ײ�*_ߕ��^R�/��2�JsW��@<�a�/Ut!zS���OO�����ehH���}���$�����7�_�~�`�xJ~���N_b-&�4��V?�Ԫ�D�>��F���R�d���M1D�M���?�M BR ޾�&B�y�'�cW�Y<iY��O�Z���T�?���h���ϑ\�҇�e_<����fV�i�vl��3��@��Q��-'  7�Q�ۋi�0-����3�f����55Z��P�B�b
��[&�|=��Na�ۮA��.{JHŋ��[H�*G�9�啳�8�A��2���cK����ޅ��n�χ��5�E�q��??�罷@�b��j^�`W(��7-�
o_�4{�O4
�Ӹ�H�9x�7���ĥ�T���Ʒc]�V�DC�� R���Vy�\���B�)K�(��N�+I����giix��Eݲȉ�W���?��Gz޼��DC�v�mq�Qv�>K�d�C�j�k�g�u��c�����]5��\��S� KlR�;�Ԧ���:�aٳ�0v������S}����)���J�/6�m� ���.Nɚ�Lw1�;&}���; ���fk�a$T/(7L5��kS#૯u��>��$�[��A��ө�\�v��T�R��[X[� G<r�u���b �ؠ��8>z:�d�%}ͽ���4/ʺ�U�]-
�WF6g�	+ð�R����_�����e�y�u��Y$�X��$�1Z�����2�+���$�R�9���W_���kNc7����&O��/�B+9�,��ص�.��V���¢|~H*8���9�Yb�6yGV�|�+n�x݈/f<�	s�;��Wu�UA�`Y���-�0�rG���oG�^�#���O���?:�!깁T#���"o]�4S�;��L0z��s�����[Oh�ѧ�D��;X?<k�υ�	���ˠ��3�
^�La�-ȧ'_���-�1kGVj$<"V)e�l�����}� hcB%�g�}��=bL����x)Ga�r��Ǒ2�e��h�c;���_��h���o[e��u	/E��g?��_:	���?�IO�}�����Y�&fe��'@~�i�Y�LbK��J�k��V�X���-OZ��ø� �O�<O��v �7��7sV�)�T�9���]G�z�S�U8i�Cvq����fF�g�KfQ1O��I	d�k� PqC=���u�������S0�H/�T�Hg��3�H�wQ��]�[���Lh'�ms��Q)��0�Cc��+�|R5w�.:F���fXT��/5���@}ql�7���߰��|¹�iОa� 1 �LO���}B���lS$��������V��zD�(�E���J� �(�(�Y�-A//�ZX/��k���P_Z�FҌ`�:�d��4�M���EE[4�v����~�1��EBԈ��r��D�"+<WGr�����d\�8�"��J��a�~$�B�dg=?��7w���Ꮘ�r��1:�&6��G�X�U��j��u�#���.���m#m6o�BD=��w\1$�,`�,�HJ�ԅ�{o�zS�iBk����[y������Xn����v���W!�鈣���M���\%�v�qq����>�d� �3Ѐ��~콅�������~�,��釅ڊ߼���_ȷ��̗���Î���ž�|:�8��sg=s����n�7�k�)bq�N; 3�a@w�2,ҷ��2B�@ι��M-G�-�s̋3���= B�=���}��&}R[s�m�:sQ����x�L����ȏ�\ڞ���1@g�Zu�D��oZ��T��I<��ڹ��X�r���2�K�Wz��B�}�7�u���DW��4RW!��!�)�rp���/1l+��ilq�1���q�:��?�Ez��Ɗ�l��$ u�^����[
��\���āz*�mM8��֕s:�htnE��.�����!��NM���J�����:�%1�Ait��P��0o�I����p*�:�A�n;3��>w��|�v�(�A��ԮƯt�Gq (�|C�ؙ�Ļ�?�h�F���q�*��h� �6�~���ey[<7��g��,+�q3����)�L�U���Zٶ��Sx��v&�Ǹ�Y2��x.�<^�U��&�q>��e�eG5�[ �+R�u��b��5k}o���f'�d�	���m)o���l\Im�{��X�߁0��
?��ON���=����-w��D������N�M,L��Uu���V}�Fd:^�k�t��MQ',8A�~�1zk ʨA(S��|�w�Q���ez�דe.�+S����^��^�Z��F� ��G����`��_M�%-�F`qH-�M%���>�(ȭ�?"3n�7v��Viw�w_�r����}h���j��O,�%}�o�c0)͒)($\��0f嬤����� o �X�B��8��
�:aq��<�a���4��E�p2*j��؛�D������*���f4����P} :e}t�v��g|ϓ ?5/O�4��	����q�(�I90�բI�%��}/Hm��1��-cA�N�
<K�9d8X4.�c$�
������c���*̱��z��u��d�z�R�0ؼ	�%�����v��6�S���+��#�S	��L�T��a1T�FR<v��8o\�?�ά��p���F��-Sї�ޓí���T�� ���<�P�ui1k�[#h((�n����yضb�[������� *~!���޵���al�U�J_�/�w2m@6��?��]��, 8��V�D1� �y6����w���ζnɨD!H�p��j#(옰FӝigkJ�������J�D�x����`��_��.�eK>o^Ʊߛg��f[����dT��4�����R�K}����4��#�D��m�L�������2��&Su�A�Km�� M/�5=R�&o���:M�4F�A���x�j�5p�-�^�O��'D;rs��f�e��ƿ�B~��ȒqG7"!��5D��b�C��ɏ[����)U�i��_p�992�G����Mg%�fêԂ�z6NNTY��� ���A�E�@1w�,b{�]h�f\-xw����g������L�4��8�I�_���rq�?��f��iE��P��S�=|wv��p1��jW+�]خJ9d�Ҽ��0>��yO��.ť�{"mv�?ʜjH�����5�j��AQ��b9�p�Z�[Yu�U��5� ��yY�"r��Wa7r{�߭	�&��6�L>|�P��u,K��8��3��;���9��EU#�(&�FƷR(aɕٙ�p�\.�G���D�/纖{�`b�Qޮ�d��;�Ť�U�h��,�p�K6���"�O�Xxh��-�_�m�J��!����a�~*�,����i���v�5������fyȷ�ً��|�\+�I���%F ��h��>��=��2�;Is�#���eI���HU��IGܕM$mߕ���\�(d�vX:	�Cܦ��'�P�#3���A�N�\:
��ݞ�_��׀��1tf���������Oҝʡ$P��,/��+����5蓕��ᏫnZ6��r4��e)��/�9��� �2�G�d[ɿ�=��c�P�q��+zR��RHA�\�h�wHW7�0;�a�G��9FX4�.mj������d!$)�d��0���=Ql�Z5��	���������d��W��=�CF�O�jКP�S��/��˫|�[�`Y�vK�wC����CJ���������K%D���
H�k�� �OXC_�����e�7��P�TCn)��b�;�:��f m2�ͺy��;����O}����y7����D�0���/�����PV���+o�U��3W��f�ʿ~V��?P��?�:@�'(�<�M?�2z�{����賃E	��t+�a�6��s�L]���{���p�G�~<j|�p��Vca_s7��B�'�w�Z��.K&�5�W�IR��g�W;�:{~��l3h�<,d��73�]ዻ�������Z/F6��㨣Fg����7�~Z!m3ނ�6m���:~*�w����M�e	��!4Bû�o��Ф{¥�������^Q��U��*33Y���t�E�P1��9%��>r!Ǹ�CoQ�������F�f��t�Ą��2�����R�1�P�.ZdjԎȲ��Ș�v|/u�w���Xr�r�0��pAN�FE��u������T��3��n,��L�Y����O�LJ��OzݑC����W���_y����_�����Z��x�W��4���r���ߗ��0	 ���z��ڤ^�	��E�y�܉\e=�>�w(����s�D2��Q��9��x�X�l��H�Y�꒤��4������x
�H��o�a��d�'z�����ZM	��D|�s+���xz�o���d�`�o�[_�f}���q�تy��ȡ��R��z>�c�}�]�>�̵�qn�RM�ܰ�[D"�m�S��m������{��>��&� �-���ږrZN��KR��#�.����E���-d2z�|�C�M08��������FY!�"�YÜ\�u�U�
4����(�58�����`u:;+ 8�Ř�R*�@�[��V��%��ع�K��DΛ�UCL7`Cfn��]��T��Ite�s;���m	G	7O�9\C�S;&�V~�N�Y�����ic�A�����b8�Y��r�\nz ���6�����t��$����auei��i_�yRU����Y�`{7/�0�!AuFi�Z�@о<cL.-�,��}�.iL�lH6N�S�j�ݲ	�}~L�?�jm��h\��9�pӆ��(d;�d�	czd.�j���|��iPn�aBρE:�cV���y?�z}܁��B�ˆ��!o�B�׳�����[=�mT%���*¸��$7 ����'i�U
�J.�/�4��t+�B�@�1�&��d�HvsG����-P$C�&0�f�FM+@H�<T�|��]�����ϱT�U���G�0�������P�����	�润�|L1�����
s+�6�_-g9��U����S�K{�7UB�L�M�&5M�*`��+�^NzR�iř���̝�A^�iع-��ϙ�K�����Y���S������p6�w�f�k5ز'�ʮ&�{{|�"b�C[6�����aQ0�r�u"3ĝ�J2��Z���.\�΢�ѿ�D�*#u���ձvɢ4%U����C-��\=�8!;z����I�Tv^�ȩʯ��<�iA�%���3��eh��6�âu�ؓX|$:��	/�V���&o*F��m�M�`a@�A6Q	�|p�����u��#���bc+�I���:HVɏZ�^}(]�}hWS�	��ٍF�ђ���#�n1���'�5���M�*��"9�p�ԝ8$�c�;��,A��s��i re�8�������dtRC��R��h���ӄ���(�p�ΚR`����fu<�����?��8!u�]�d�QG���\�rO�j�{J�d![�xݺjח�㝅d��3�%7�/�x,*
B�������g)��QH��_���gI��M7ǯ_W�����Hi��.�� ��T�6�;��h�d�E��A��3Qx��;�P$&�����07�
�x}ww�n�%i��oe�:�t��j^@~�|z:Gn]��9�cKat�= �]���r$���7k�p�O�k���ٟ�zD�61x���uI�6�T�����Jm���>Z%;���xb2��� ����J��i���1�p�wpU�N�� �v������8L��,�H��wݾ%�kV��T�TX�sȾ��z�䟎�x#C*��Q����R�5A�{ec(G�e�����g?��8��v_ߡ�ò����� ���"�_�n㆘5�P^�"eQ�K��!�un���3�W�3�����w0Y���i���@�8�G�W�8�2��V�9Ppjv�7�2u_Lׯ�� U�cr1^(>�%9�az�Z$�\����O��;J7�0L�sq\�,Ӝmfӣ,�m[N���iW��X��]A+������	 H�2�?C��,�6Ù�|��OEUY!���ޜ_	tO�g��J]�7�#.n锔�`s�##�����9d� 9ɶ�{��mޔ��2	WQ� H˥'���[ۢWgL����S�g����H�k�so����|��ۺ�ۙ ��Z[+R,_S���5�0�#���uא�������WM0;�EO����_���#�<�\�ι�5�1�rL�n�c�^Ihu�k����w����������o�����yW-
�cUKZY��u=�t9�*?�BRw�<G-�������n�
�͒���?:�Wrz����p���A�fJg��0��v@�Qn�9��,])AX�ˑ5���,b��KϡA��� HH�!���!4G�IQT[H;�ƀ* �PX�!��ՖVQ��<3�?�S����ҋYW������EM��Um����n�[�1ۖ�7�|�t�=�JO�8|�J�����z�A&RJ�;�~kd�f���o��!��v^=��+�N2�古�t��z����o�j^SzCyvG�ͮ��Cs@X�p#mh��^�3<����E�a`����PG
���y�LP"�0w�n�h�@oR�8�n݄�����+����8��`cB�P�Ũ��������F賢��=��v�WO���T���i&F���}DG���E��f�R�V��x�2�|A�c�S�ʇ%�HJs�NU�yW�:I~��i}�b��D~��
��A9�]�'��ERJ��Wς$����3�|M���8�$���؊#��m���)�r�#�����q�if���1��!w*b.u��mo�V��D����G1p��}D�������� 1�u�'����=��Go��s$#z��-G�:N8��aY�*ζ�;��1͇[���\I���E��A��!��Q?�@S���Z��X�����@X�LZe$�EaM�u]-�g�d=@o\����ˠ}��[�-�jV]� c�$����s,�oY:�5����ϽC�g�:l;"�u�ɠ!jӹ�W������l��׃�0TI�d��=w�tܲ���H�Z��fX��K�J���H��ne��&��"	��d4��e�8:���7j<(�K�l�`48[ˁ������z��wi��g�r<�2S�F�ya(�Mfd4��|��ޤ�oV�1��E�����䴦3�5g*�^A�6(�WP���n�T��8�j�L0a����5��jY�d'ҙ��옼�}��`?O�A��Eb���y����D�z����:<*�x4���y��Bc,�^~����LZ��I5�7g�ED�P<� �J���#�ɉ��R��2��$��7��/C������܌mXQ�9��+?�����3�ڍ��9�D�6ը;ھ���sھ'ȸ��#��m�M?���$4K;�m�I9%y��Z�:�^�����#Z��]�]_� b��U�7���{�"���.��u5A<�E��P�M�E��Y�:�]D/r���:h�#ʛ�'���z8]K
�Qa�~&U�вL�x�yP�������ߍ�,{���}I�v�#L\;�R�3ӱq3��3����/WD��W�~T��tM�ϧ����x�b;p��(s#(����d
p�<����_��_�Y��0��j��P����eM��\AS�콏0Cb=��Ak�D��P�.�0z��Ė-�;Ln~C�H��	gR���
hx�J�͚����p�H��3��D߹F3^&;>���*�朜'����v���kT.�V����v��N ����7q�0��8 �{�����x�s@GB�� #�M޳4H�M���r-\��+��%�R@$i�.���;O�m�W�BH1r����X,�)Oؐ�V%�V\et�.�>���`/Fg�$W_��{m0�ʝ�jG�������Hf���q�M��l����U"<_a�	����`"�BĮ��xn�E��J�(f뜚���?�w�	��KȨ�@�\3�����A5-M`��8Nu lf�|�����S��Ku}?*(:!�$��aO7�Jyo�.p���.2��]��	�9��mj1�3	 �tj^':�)��񺞃Ώ~m+�����o|� �������k��İ������vL�T�K���%��|����� 1�B��ӄO��rhW~��Ҷi*����m3&䱬6اU\1.��Vd3�S�%�Їހ�0�u�L�`�j�p^��@�z��#x�r:�G�]I��#���H�s�:1fx	Z"�I��SSHG��k�3-/�v�0�Mn(vٽ�"l==�����N����6 �&j����A�f�GHn�x]�� ��a�-'4�R4�ڴ�a��G6h�d���^�!\�tK���b���$AEA
�0(�~���*F����A�A���]N���i�G�6fSbq,�� '�Kӽ���=guG*�Иq��N��p�C$�Ns�l�9}'?@���rj&:�D��d�P�&.��|0#rY��o����C���+��[�p���g���9����
��r#��C�
b��f��U�J,�ɀa�ρ����]N�4-�V����/?�d0�w1��� ����**뛆lI^�Q���X����Kn���eL(+Ft�o��M	Al\i�����o����V`ng�?eW��Vܘ�/��[�<v��E+H�������1u R��@$��$�W~G��)�y�S���3��jxOY}���lcM�a��L�͓����|�d�u�pb�cf��MYgHbk�_��}Nj�;�{��c�Y*��l��UX�{���h	%�����(*��fLP��B���p�t8�^��C:�N0��Y�?Pc6��(��00��M��g�ݯ���2�Q�{�?�)�=��e�,���^����Qǌ�� ;^�X}�{�β-���]���v6���[�7��c��Ҹ7�A)��C,��8/8��: ��:{V�|.��Q�W�0mH��qo��.��_#�V���Fދiy��܇�uNWЕ/H�LF��H$�C|�X�_��^�߱���Ŕ��S �#䕙��O"�ޢ��|m�!!,�w��HK~c��\V<�g�n鹌U�;Fo�:�T*��T/1�'?e�o���:s�y��BN菝}v}7��׀���j��� Ի2H���i�<�	�D��A{o7�p2�hܜ�� U���}OWy�C��C�2�3u�b�p(��W��4ϧ@���5���;�4)c���pA!��9�`V�����C����5DFN핌u^���95��#��t��6�Q��<n�w�����?$��j���It��8#�jO�y����v'ֳ{|�/P(t�%�j��̅T��� �Oog�^��Ȫ�sD�a���"�"���׀�\�.#k�b��@�AB2�p���8����祭�T��d��ͻT�w�M��-�a=k�az�u��>]&��.�<��3�eѦ�����G�K� �^��-e.�9��ǠN]���&�"5eI)�߃4�0���f OvS���.�ڹ<�-u(ށ�N�BQ���6�RJ�Z"�e=�S���O��R�B�"����Z�*�{�X7&���=K'l�S���=~�a�p�I���T��U�B��/�mNԴB�K �x����V�T����x�>�ZiQ��t��",@�Q�ϑ5�;��E,\�:Yе� �Q'���c�������ud���%{y�J�~��4���,| !�qғ$��������0��,v�����.n�p6�0[i!v�NS�������������-CK����k��Q���|eF�锃@q�ɲ`����K����\��J�jȉ>
;�1�r���N7vc�e���1����!��Ս����=�o��x_p�#/��U�$<�
���Ĝgn08.�����ل�P�H������EĎ�+Ѕ\����$�	�`�C��MAƆM�}T_$��qR�w(Q3A����J���Dq��,�D��˯fQ��&}�ҼΜ����-���RW�>�.��r9��f�fG"�~�Sׂb_j2c�8�{V��`D����mZ?p��q��/:��L$%�-"%��è|OX������׀�@����#��s���u�mg��)�$_��+|��h�-���2�hii��*@�� �ȸ{��mzJ�qm̓OK;�?�0h�)��2�VD�(�r�嵵��#��G�������I�����x����=?r�F5��"ʉP��+�����x�{���њ��(H�rzL��O)q��F
�9r�o�s��,��͊-B7r��>��4ǿ��\ܶ�9�AN��}��fj`_w@$dC����zL�қ}_�G9����왶��Z0�.�q:�ĺB��y��،���U�6ꊜy�8in��Im�e��uT*rJY�;{Ie�������	�D��ڂ׶���]k}�i>M�`K�m��u�]��1g�Mr��$ź�0/�`s�([r��#L�.�f���kJ�:#�3��-}�#�|p��m{e#(�VҰTUg-�uV��(�oǢt��+R�t:�?��=BP��F�[�v2}�i�� L��v�J-����1���W����g]'�sqX	~C^��\�����]'�\3-;�h˸�����ԩ�Ӊg?4D���N�o����
�`1��(��3{�������Π7D~`�:
{ �(�0�u�'{)ر��#����+NeY.)h��C�8�I4~��k��t�L���n�Ә���ʪ��M�o�k���	��k��_�u�'��ѻs��(i�d_m�X

jf�|	�A{��kK{X�(����x�VK�_PT	���~;TO~I��Wk-9�?�߲��8�ؒ�;��%��+t=4CG�PO��{a�ME}c��4�,ܻ��ϥ�.���~�`��{�� �9(��#��<Q� B��:�`cRt�{̑�M.�
M��,Ss���*34�#,���a�[�	b��a���m����@�sV����F��,�Rk�M��v��A�"�3'曦$�h���Uj��;	�ק�@KJg��|&,0&�����a'٫�ܷ���6����^Md�{J�\cN�텹�g��fC��Q����ʋ_3����A��\b�K���5�ٗ3e�u��_��h7�!��D��4f)M3��Y�	\�+���MN��$�},�5-�X�k<�	�®=j��y����v�CQψ���������:��u��F=%�ޢ��v����� ��� g�GVp��k�h��Ӏ��k6$��n�P�?5�L��*�Ejk'�u=ԙӳ�:�4玶����Z�&2����<�Ψ��������	є�<N���(k�nU��W2Y�4�q����s��If%~S�KG��y+��Y�q𶙯j��i�W� �E�4������i����2��@1��oW i�ʴ%�x ���L�F}(?%r���~��c�B��Z\%""�.e�j����C=�E��?�.W�Lv͚�7hP���L��� �-��"ݱ9 �Ml�cүf?�~��/CU&kc7P�d|��y���m�ہ1�����ώ�ٟ]G{�ST �y������i��8Co7���O	�՟SA[-���^��3C��	�c�v��D0d����y��I�b���NJ�^�P<a��4����]���rR�-���ȉPB��i�����l]�e���g����H0�p�CSS����q0��o�/s$�;*$�l�=�&	���t����.~!"�� ��Ā�������f��8�6�bb��S��D������(J�E�S�YltZ­Mȭ�
T�k� �z=o��,;������%}��?�f�U�߫Q�ǖuaTyV�n���0���:C>�fz��b�~Lq���np���H6�����)�O�q�
���nf�9���Fz���ߖ�����w2��DU/	xvB:���(�N����<��Ë��{,��Iz���񊗥Y��ƴV0o��
yG�8'�;��4L���<~�Kc{��Ц�?D���e�^�$��������*���X���3�����?V���0@]� �M���	7�Ϸ�G�{���ک���(�&�FЯGB�I ��� h��А���p-5;2��]�)��D���5�&D��X�Mw�ʼ4ay��ƴ��A%�0ϩk@��	:��|XH��X�H�9;E��K����h��&��B�K�Ch������shl�X�ӹq�G��V!�R��V�?ܰ���VcI�Ŋ�J��Z*R$������@��k�����E��#Q��z����MM_�&Ji9^��G�9H�O����^��I�
��߰l/d�E��I �b�9^rg�~��1T�;9)7��_>̉%&*�Ih��J[�~o�yog<ud�L�s��D����tC}Br:�V4#��ժ)�4���r���#�
N��� w��d#;��t������&
��ǝ����0�����Ce�e�pZ��*���|����1T�ʐ���Ͼ%^�%�F^����t}��^��.+����هI ����ʢ�n��,x�f����Ho(Q�H���'r`�����k|��΢S����}XG��fَsT��~�&r�	눻��S�
�o�d�C�ż��3��Ov�4G$���5ſ���Y��\�,��_0Ek�vu�����o�	;�b��]�S��GHxѱ炞^��}�����<ˮ*�H��E�C��е�;��F��" �mx^y8^5�%�M5$��k ��@�f'HC�����ٹ�~���Z;(x�U��v��X��r�ձ,P.��eF��V�I�L���D�Ź��F��%H� �\���\/�zW��p�ɌR%Y�C �q�lqՔB��,�oB�֭'��w=fi�}v	FY����$�@4:��>��
�g���Y�T M ���[�*śӮ�uWr���������ѾB:�x�O��"�>{R�p�K���& �[�%	�0��uO�����pSq���d�ҙϸr��a9�s۸t	<K3WrxTV��-B$�iq"��O� d$�h꾬�M��_�����~�	��ΨH��`{%�7�nle���s�`\�	�������ͨ���������Z)辐�ɟYU(C��;'��G�҈���s���*�o_>n-�E�M�e��0^y��'�g�F����1y�����nM�P5`�@�C������v��@J���!�{�ᾩՊ#݁[�Y<=1'��m�}F�KkWј��E4.7/?|!�ti���%ѧ���L�b���#-�R#h]2t4.@��D���F��	
��nua@�ҵ��ͶI��X�B�b�Y���O�f+�X���-%�����!{��Gpq��s:-ʱ�H������:�n��c�D�I����-q{����:@~q�����Ω��82��O+3f�1�N���"��R����N�E��/`�T�اvXo�f^��U��Lв�.u61�\����	��U�����/1����B��Q#x�x6�����3�1ʩ����RF���h#ڦ��~��D �F���C���k+êc]�fW���j�%rUI㬧���OU.`?��|bgcL$��B�V�>v��8E#H3:ۢPz��w-"M�&�Վ�${z�TMB��A;1ê��Fy��0&'�}���y3(y��f]��t��u��xr"b	�R�͇5ߵl�-��@ޠ�iG���I|���t
[�)�ӕ\U��ѐ���,�|{�a��'��͵4��|.�V�;�8�^Bm���ۂ#k���}ٔ_��7h���{�T��2G2��9�F�P�?�:�ݯcy��)�녁��d���^�5f�)�k�������K��_#B˂K���������`%��3�������$q�+p2t��8���2������iw����I^�C�:���Wْ�s�Ϡ�r ��.�eN��bw�jĐ`�1\��@�+��m�
"8~1����?{�
,��Y.Ԁ$��?^�$?.�����p��æn�G�kܫ�G�'.,�!%E'�E׵l����	�Kmt6���6�(5�c��R*�b��ŭ
T�������e���e%�ԟ����i���޵x�X6C
������MsF�����r�_FKbGED��'�Z��W
���U8�k�Ti��-�,@7�n�i0,д�#+�a����@I�hmBtv�S-��f3�*@О�mp�>͌��;�8����{ݙ�jN�7l0X)c�����K���tG*/�bF�D����6�e8��z�1h/�
�L���ɓv��u�D����C-y�ԞK�OIe���Mc7!k��V��/d�v&�;���؇�P�*����s��<�:���6����o&�j�a_�-�����#�ch��������,�����a���v_������vB�:�tT���b��z����q��&F;����H=F�눡���Kb�3J7�[cmd��ڴdy��fg����}��Bߦ*�ġ����ڛ�?\���v�(�Փ����}<U�v��m쉂II	��{�sɹ��6��4���T�i��a�I�z��#��6n�,��
�S5O�!�S
�g�|����r~�y�@��-.�o��� ݙ
3�)�����2��Z��H�'$>{Æ��7X?��w�KA��y��+��	,��Yb��v��"˽O�	�0Q�N^�X	X�����0�x�ͭ{���KfZI�:��_5���@��z�$fK������^*	,pG����ZP�:gro!������s�� �.t�g��Wƪ����2g��Q1�u����8��aD���ŏ� �xߕ-���0F�#Ɩ�5�w��+��]��K�{O��+Q,�>�RS)�ꊔK $G��/�-�'w�׊�����:�[��Ù9��Z���S��k3�F&�2���?k��;	��y�囹����F�AttI�T�h ���.�1�Ƒ��[ �}1vc�c�O<q����s0���G�q�C���jSaB��γ14�s*Y�D��D�`���绠@K�����<}�O`�2�֢��_9%�Q���t�L��V"Au7y�l�JGj�)/~4'�U���pw4�f�@kKuu�v�<�62���u�Msc�ڮL���|�"��R�-mZ��@����u���x�՜���������u'?�5��/lt§l�6r
0 ����i���`|�	�z�!�!�����t5��ܰvЂW+7��J��AdM'�����^6��6��Tu���hrׂ����O���B���}�@�p)+��q����i ;&'Q�(�:1�����r�~�x�K�CLw�EGmrj��ٴ�ˁ�t�)g�>t.������M�om�W©?�[xeC��2�[ն�׺����hX��<���� g^�a:�N3��]W"�$`]!�L.���g��ad_�pM~Fm�t�=��xgd?��b��^��9�v-�m�1�U�I�Vp�^�0Τ:W!B�R�HR-޻��������>��� ��/�J���(�Vi��L��S���/	��Y	XChk�E���^%GV6)�Q�ߘDMę�FB�b�Uρ�Ҥ8T�����t�E�畹�^Q�wt��_\�_ 8^�@�Ʋ��Ո׷H�`����a `��G�b���>f��Sh��o�ϑ�7s���!k,ʴ5Y��{�����yq�� �-�+d�6�:aK?J�z�Y�rW��Хfd��?H��U�<ϜR�B����0�b����A�c�Gi�Fd+(ț3ʚch�0B�C�N���l��"
m��v`H4n��j���4��f3�
�P#}��I��Zq��ؤv9k��Sg9SH��><|tFxM��^��՜>��}��}1�x���+F���O����(��"qM���/��p�ѦI�`q���3�g�|��s���&wH�����%�������>�Q<�ʿ�A���������7`RFhGn&�Z��<~b_�q#���V�����Iak������nM�UV��|=jQ-��M=gҸOhb�՜sA|;����V�ig`G���!v�uV���_Sr�	��K��C��[�^��{{-\M# ��c�o	Y�����rM�5Z��F�s^���$���eȿo��n`w�*� bLG�#� �О�j���:��nqrբ�]qь��&*I�B�sZ"��*YhPD��M���T=��p�AK����?�[�?��`F.Ӯ}G/Bi|r���n���4����`��_;��ˑu��e�d%��)�(�;��ڕ��U��u�*?w������d��z%��Ծ�K[�_�x�ٕ���A�C����fw⒔�A����R�(g^���S�ɲ�����C>d S��Q��G�,�e&�N�z8v�\���g��T�;��Ó���<��5��J�"�d��A/�d	F\I��� 95U�oAJ7��Ҙw�x���m��d�"�]32��W)a.&�ǁP@�&N�fL8b�QS��͏^H@���w^�e�� �:G$ZN�?���M�Z��7��<v�Zf&�� �348ii���I�������$�4n~�On��^�5aMBט���N�\$��/n��0C�%.˞� Ѣ.�USq��ӊ�ǘ.�3ŅEt~�k���R?A	l�$&�z�"��\\t��bY�&n�ꌠ���M�4g�R�P��:c��E�w�p��\Z�/��(����A���r �f��j)<��i4c�F����K~j:	Q�[��:��[X��L*��i�_!8�ܧoi{�gC��ԉn��S��S�	�L��X�4�Y�V� ��'T�H��y���?�ل�	�Ǳ�����P8�#�5�VqF�D'��D �ii��.S�$��V��-�@�WЁ����'�
)�C��^��T�P���}k�5S�O3ֈ3%u��q|��ìʦ��v,@K� ��> K��L�'���#z�v�~�n����L��NZ:��\Z,�o�J8�� X�އ���J���L�IkN}��]�$�u���0u��y�bGk�J�

�f��^5���%�ݪ�L��M��{lJe�˦D2Cx�d�3q��19�"k.�q0�&�-1c��u�W D���g�n)�o輝�i���$)�_�n�˝~S��WL�^DѦ���]sd�7�H�O�}F�(҆F\�bRe��]�Y�$vTo�K�q0�VS�f�iïyt������(鼪ؗ�u���!��uw��nh���/�We��2ʘ���%��p�	�h{��{8q��W"�2���t��m�( ��q�VZXq��Z"�uw}:���S�eݦ.�J��e-۔o5vg'�����^x��lj�����N�ޕ�Xl?q*U��"]F�^����L�҉ �s�=)�	� 6��i��d
m
z�F�t�F�Tk��dFc^��s���H��
���q���y���L��C���e�ߧ�n�#�>��d����5�0�Зb���|�@*�{P��~�[�ӂTW&&�L/���%�l��O��x����26ũ]�3���NV+7�e����EQ�il���=�@"���
4f�z��?u���ɹ�+Q�����̴Kr�@���dp[�¥�6�[�BQ���*��� T/�l=]��-�4?�J�;�?y�1RK�:.YA��,Ɯim���������/�&�f������������U����1�*�Tw4��fQ3�ђ�m��A�� �RR�=�N�E�/nD����b"����3&��j���D3R�b����* �E���p�^�
��l���9��?0$���K���7���c.�M�kv+/�,��&������C���<�w�/�a��� ��(qB���	>�'f������/ߊ#�9o1�2�P�03�/�Bq�CZ�j�x]1C�.'Oy	�X�uK�,Ǹ�w��#��J�óPaO�(��i⳹U.A�֒I}ZFC 9��<�jҝ��-T���'��OHW'�p�"����u�Fl��"Xh�\�c���0Hp��Fz�Q��2ϧ*�
��R�G8��q�(��__��q�I�T1�A�Opy�*�q��6���zI�m���C�sq�>x��Y?Y����F�9f��U�:�r�dx�4���fO�"��+��_��2�b�c�^OĴ�+��G���f�R6��\���WT��)���y���/9r���ݳ�e��!Rl�� ��@�N�<��e�C�;Eڂ�)�0�=�J1m�W�n^����g	2hQFQ�����޷��'9���]��)ۖ�]J���i��	�1J ��tڨ�r�������c,C�g+�y?�d�+M�9e����j��z�Gd08j����Ył��O]m�V�{ԇ�����*�w{�}o�H�_���_w�W������ ������b{��?����_�������+D�`h�=^{ z�ПP�M�%[��>�:�{^������>7�C2��P�v�xt�|��8e��3�����"���o =�P�X=��	��	"6�g:M��熝�Vjw~���sR@��|T�ai���4C�4Z�.S!���@1��N�K�j���3_��vb�V !�3���S-����w�i�a�?vT�e6x�a{�;f!�F���`���d֑��tb?����� {��P	v�򫈢�$*ļ�>$�"S��AU;c�^��6�������9�|9.�[����,ޑ�B�T�q�!3�|f�ӄC5It�w(�I-7Q3ن�:��CB���R�n2l���UG�G�jxc?�zh"�����r�k�\,�a�&;�� ��|�%d��ʝ��bY��j0���a����$����O��M��<9d�U�D=���X�B.��v�RKr����vxk�^����a>9����0%��Cm�^�!���O�������*�װ�U�lY��Z*��v`d����<������E(ر�t�s��xf�<�G�9���p13X>s	o�36��4���tAz��>k�F:��O����Ӓ�"�a��r�_rc�Y?>c�$A�]�f�z\���e��;�2���2Aޯ1q�OD�;=pXD��eU��~s���h�y��=��R���m��3���EL�v��g��,�'qP�~Sլ�1��E݌��Pv�M�=�w���8�}��TI^ލг��u�l��#���xJ��xG�{������:tR�j�T�~���Щo�T���ݯcQz��u��tU�Pa@~'�cǇ�I-�P|P��s�1�˭�*�$�%��	�aۉ5q��ס� �ֿ�s�?��^��P9]�!a�5=��S���azi���)�/XS����ˣ��X$xH�`r���-���|�ka���Ŗ�����5�/j���ѤqUc�;�4�\����*?�!R�6�yh�fsZN��2H��W�-E�T��L����5k�;���t�G��� �������b��KX��[�x�~���첋�Y��6H�M�ngv=�������	�W���>u�+�^!�A.Jqrh�&��-2�shKO�}k0G�k?���۾Ϟ���� 	���Y�'Ue��?b7c�gc?�5'�KyK���{�@
D�ýc��W�|_$�|�c�Q���e�Ȏ�#SA0�4q%�_ �~���l��]�k|U���Ǽ�\�E+ћl
��I��8��C�!�R�ډC�d��*[�)"�7��2�T�3��#:��^e'8O�Yh�
��b
WvR���H�w���e�cs�����e'��q����!����4-���6)��(�v�P5��&�e�Q�}M�L JW?�g��d�~ԙw+-��IqhA�E�,	��>`��>rnџ�1�*��U��\O��d���l�\ri �ԏ�:=�i1ߕ.Іg>):?^7�َ\£u�󙧚��P�1Ź���E=�=���D��F@f|���!d޶�!�ރm�E��²de���(�nH����b�;���r�d��il�yb�^��d�?z�0�?�4�ϾV]�E:I�՛�U������+��!{xn�+o�>��i_-� u<؜�%4&��V������J�V�O�����q{z�zx	�vA� ����M��V�J���a�u��,�֌Z�`M�w�:)����t����Z����a,ۖ/S�tG_P�9.1&j�^�uQV)EJ�iC���#̢�����Iq��+��Y��9_-��B�@=p&�F�ޗ���_@N�Y�Z�JZr�g~#n�PN�<�J%T��y/�c/IK"�ځ M�o�%��G�E��>(����Ȕ��_v�J*?l�Ad�Sa���mH�'Rg3�P~fx�}�\�3?�zو'�8������V;5�ۻ���/�J J��"S��O�j[̉D����@� ʓek�Ş,���&V�b��2���}GQU��X��O+Y�jAkh$��$�B��AI`���#�*"�rE{U�.�����ᅂϢBZ�}���
Ӎ$�V�S*�G+/rYucbr��p��EU���ѥN��j�]�y����c(J&)�퀋�����vj$v��C$��A �Y'�n~=����G�m;�@x��zެ���1H�K �5���*���T��lc�I��~|G�Ƒ�p�6�5	����s�A�\G	H��}�̿�Wڙhre�%�R�eKX��ȉ��`�������䪢�]����
�~��{���p��3�f6��Q���S�!]_�ị̑8��U�,��_�NxЃU���#����KF�1ھ=I�]��+�>��`�0=���?��= j��}#�C�T�A�+�K|@�J:bĦ�_��iWrs�k�ay�e=d�cG�	���WC�3��OӴ%�E��V����܁ǆ�}:���3�𒹞s���e�r����Z��!c�����sq��1�����)�Z����(T�>U��R�q6�Î�0z��ẕ̇ d��,����b��Fџ�Q�|�~��a0.�[K@���J' sz6r��ɫ�4E3�Ly�R<g%��OJ'��ʻ W�*������u����U�X㡫T�#m�p��$j�D���ᦤl[4�i��e��cI�w��C-R|bsoY��"�I{6��ľ�Y-�w�,j��) ����|{T�@���"�?�6Gf@>$�&��vޡ�\e��gh� �q�u�>�G׍�@ƋCpy����v���	�ݫD]� ��䑅򋎃B�+���:���`Wٲ��\�YC�`I��GSiT`@H�	'��c���T�D�ԲQ��)���o��'p2��ݘ��5;,�s���qn.�T��m��@z�ԡ���-$��Z��~�K"�J�0�����@��g
�8��fd��[�TC��� � m��W��tO7����>}�U ��m���w����s�	ɫiKޙ�덦���8�-��Q�g*$���e0��͉U��,0�v��сNN��K+������d�s��D�&m�33
�q�8IL86 �_.�R���&�ƚd$���)l��2���7[ݎ��&򞹞~�j���+��{D���&����E�F�n[(}Or�3�Gy Q0~�[�1�aP}'��S�'�^�Y�et`1[��B@Q=��ϕ�%Mmf�z҅3�0V+��=����CTy������U�Eů��������r���`�>ƢW�"�W-ـ�H�����aP#����D�L���@�����7�1%9��]嫙Ҡf�P��Cn�/hj���������F���I��\�<�ر�*�8����t��ە��S��Jն��`�x$I��X�|X��K@g i"���G�H?�y'ĉ?����Zm��oP����Ae���S�NG���V{�aa!jO��������m7��"�L���q3�sl��p���/�uq:h��Zyb��7i�B�������'P��DPM������1.�/4`Y��&b�����s)�ԧp"G��Rn���J��'�	�Ka���%�hqPT%�i_���������Ib���tʍ������h�
�s�V�Zc�մ��&�WrM�1�+���'��-s|��u�y���|�^��p�c"%%��@ ��g�~u��V�������� �P�:��ӫ��= 8)B��쵅�OCΓ"R�)�*H6�1� ���N���uK�5�W�م�(�-�Ma@��t��}����$5U��9��~����7:��`��1�!�6(a	v#B(SA,������]�B��s#[n:��)}}3~^���~ju��q�]Z�^M^s��rL2y���=w8.�����2p����tm��Ɔ��m�ؗ���T&�6(���Ehg����<�3��i���Y ��q��i���9cԔ���"�ǧpƒ3�NV���m�_]$���Q���B�5����d��4�ﻒDA' �&�>����g��]"d���6����셚�����W�O�7a��Z	�p$/��Iwv�%dcx`]*ͮ~ce�P�U0܊\'�u�X���rK�<�S�,xx(��b��B��[B��<}pB�u������(��X�.4�� ޭ�����T	��Ô��ۂ�"��V|7�i������I������5 6g�A��
 yu��Y�]P��[���f�D����>Y���+�]..�~�\��#i�R(fƂm<K���oL$[L��_��J�U�������t>���V��;�0=��=������k��y��B�Q�{�� ���9VhEw�I(|3�eO�x�`���ƧHBi4�i��P�.�P��C�n�@ϴ�����1uB'P&�\�6�^�I�3��S���3U*�A)y	�#��9>�d�G�u=����b�-@d-��*
������X�~	��h�ee�h�))>8w���nɠ9��� JpU�$
:F8�3���u��E:'K��?Mn?��?�x�z�j�����`]MHm�>�*�*��r�7[�x>Jd�2�;V��B;��#|2��m���j��/�ۜ�4�[�z%x��h�3F�`��h�� ��՜�IA��3Ŭ��(y�B���מ�Z�f�K�jX�3�f���(�G޲�/c܀��U�B��#����=��ݽ��@�N?0���a��N!d6�J�%�7S��Xgu�W�_���4,U�7F��ws�E<���HB*EGC�vµ[S_�颣*GA��l��q�#�B�ٚ�3q��z�L�f�fHy�Pӻ*q-��V�[���O/�P�=�F��$�*�ԕ02��eK�+;z��l��en��lE���(�[�.�>�cP�/s�b�Z��+phǎ:��~�_�J���Yg�_<?S*_d���ګ�dh�������=v�d��V_@y�r+;Y����؉M/T�xtT���R�/B�L��C�=r����=A:���CYɷ9�>�K�{��r����s��T/������ݶ���L�Y�L�3Z����-�/R��!,�ؾr�x'Z��H��[�h�r�Zd�e~�%����m���ރ����q*4�a߅��q.�ѯ��.�G�c�Di���1'�r�S�2���uN�K���K�-�ժq�L/Z:K�b��WCg:�j3�%���ݕ+	�R.�Ѝ6j��](�x���qZ&Y���A�;�`��Q;�
�Q����A}�;)�^{�	���t�&����}�>u�b�v��6i�2���������d����)�5����M<�䆪�;o��$k���֘�e ���0
���xu�{�u��o�t-_뛢��ݥtq���y��,�� ?�C��u�������+O
_R���@�v���XY�8�H�İ�M�F���JKDS;�P��z7y��&�=�H �����3\�Hsd�Q�+�x�����In��[B�yA]�͹Gr��{�o�,��Xҙ7{�g�ȉy[{��Ƶ�E)�c���R�� T֝����|F"��)l�����>�]�Y�x���;,�snf<=��W�P�Y&��Z�20Hma1YT/xd�z�<a�u�-��8ǌk#D��uH]���s�t�>����V�y����0�1ţ��Q!�ܺ4���ϲ���]���&:��[��_��3��� �kf�g�0����d���w[٪�u���������FX5.�64����Wv?��[Q�wj�:_�M�D���#b#��"q���s��	x#�%S�����1C'S�Zy�glD�;�՟����+	���Ɇ�=���^qZ��B4�Y�%�<vة������ة��L���{��=n�n=Lu���61��<Dl��(���A��:FQ��EK��%�"#�0^"��em�9
:P{�>-���uy��\�D �.���v�v����＄��JL�SC�R�IG"J�mc)���9B,�4x�r��nԃ�����E��2�#��a�.��g��.�(6]]�(�U������Gw *:lA�CK:�*\#�Df�&�R�Ĩ����0�6�U]F�#&����F+�э�	���}���.� 7�.�k	��I�6�"�����6�~�S�S,��#��~�vؘ�V&y0yNj�|�8)�h����� n
i~���P'�����y����(FH�P�щ��z�A����@�����g�S�����f��1T1L&�a��)���E��	�l�۹5���X��i��Y��47�k��A�R��?2?%�����g��S����a�Ȧ1��Qɟ%�}7�n��/¸�{���`���R3��~��)�k?r�~��ߐ�)�]y����k�����ڨ&=��]���'��j�چ��H�d���\�XCl��c+��Y,�rZ\�,)��/��x%���4�3��,��kS 3�&��-��[u���=R�1��R���4�����M�0ҳ��\��U�;�g��xD�*ޯ:��8��)GN��8Px�H[��Is�3�TO5�����q����׏�X�����_K;_�#�-~$O�y= �����E��-��*D��RH&{q
��[k<T��lT�J���l�΀��Zȱh5
��~۔8jf�tjV�l��1�Y		�Yza+���s���zJ)�/���,[ 	vG�?2ȓ�m)�l��Q7�c*�JFV.��&p���l�`gy�m4!1���J�������Q��'0����3z���G=_���O�	G���������c:�z�O%Up�^�ZHH��3<�$
�����@�6*f���������9�d�sT�����LY
#���$éD
![�d�' ��`���9|�!�>��mܳ��~�X�܀z7X����D�v�O���!e6� D�5`�:��wѶAЬɰ.���^�nÛ?s�*�ׇE���Dx�L7��6�%&�� V~�=�p.����u}����4[@�%���ti�l@qWc�t��8z��{,��.��S�lܹ�`��"��I=�,l��(0v� [^y��vXK�o�K����«1N7g��r�e�9E�0�2�������U��÷�w��N�و��5�+'�F�6GN�[��@�4��FUlPaF��.)O�C��3�L�&K6�8#���,S-kheBK�CX���s��`�WK�T�~���O���>��Q�/P]���Њ[&��˽ʓ
x�Q������bW��Yf"�1G����켭"�����נb_��@/��`�+dy�j��X�zMk@�5;�̇f�ӳ.��4T�Z�C��l�[���襙�%�����׎ql�~t�����Ä�4����o~O/5��ǃT�o���j`t��<�[t@P�_sܻ�����FyТ�ZGxu��uS��u�/�L(����w���*��W/	jR�ĭ��9f����p���G]+
�r'��uNW\�@R�0`>{_B��57���K�T�3��2lk�l��8�~5���v��o.�ДJ�N4��D�v��읣�C �:c%z���%|6�hFxg$W�f�ݟ&*����T��}2��
�K�>|uB�T���\#��>�'k��������%o���u|7h���~H�߱|ܴGi�J��	����^��C���C �̷�|��I9�2aoh�Y����P2�^&^@��n`����z��d<�1��.��ʑ
ޒl\5�H�pY�Ì8q�嗪j?ls/i�]:����ȅ��4��Y�e+ �%_�	y,�@h\߳ćm��Γ=�x���T~�7�5_O���fv�����Ү�#�H�ijR
�"wU��\7�:����}WK܍WT=��	~c͖hY�4�E
��,|���� �QYw���[;g-U���د�C��g�8B~3i]�f~�w��#*2���|ΛCǒkHm�K�nU&��׌����r�S��%�
?3�\P&�C�X�a���l�im����~-��d*�Os2?�P���Ҧ��[����v�<�U��,z�0�:�8�sW�GB�����n��c�M�ܬH�־�~�fJ�u�7��4�������Q0�{�m8N�Z;N&[GM�tjPF5��@��B/�T���Pc_�X��v�iz2��mS��tR��>�a{z�����g��� B�XĴ�X�e���-���d��ݵol���y}�b�B�� �^T�׺_��i]�+�6�HM[D��7?'�Zm*�tVc*������e9h�U��)�&��Sv��orԇ.a&k��]<�$w�y���ȹ��=Z�x�������ހs�4�7����ӇYPy��"}�M?����l,�\J�*����Anf�PqD;����~���%j�$ɱu��Y�BU`oJ�8����Sך�A�Y�pF�gΆ&+��W}7!>��S���=|XI���1a�&��(�!�cG�f�p���l��k���*��n�m%<����d��G�8�zB�	KZ��K_q�'��*I�]
��fr��(
ғb��G��d�V�rI4�Q�����\̠��uΗ�&dOvK��%)J��IO��j�C�a�X*���9�r�jߔ��6�6qiPG��;b�5���ް�$������(�@u�l�/�U;��֩��C�~���&�d۟�#'���uG:�k�N�҂�́�	X}�%f�׷��~�'bIB��|�H�,�f(��R�	���`�x�y�
T(5��=�*�y3�þI%i%Y���_��׷%�U�
�3���lȕ�j]��݈mF��*�?�F�{�¨m�!%���hD�6�����d��3����=u�[Ė�,y���q�W�
cG��!1�&�����=D��������8@�h�^��Z\#TU�Ne�?]��N�	��@i��U�@��+zy�d�S�����i@�eE0���Y�!�pi)i�8�����<��,�8�����6�ê�ɀ��[W�����pn�@��&0.�sk�h����ﮢN�u]�����NG���f՝@�!��8_y��"	t�Ri�._��9�
6��� X*Øu�A�����ʵ��e9��	N�[HKWF���$������K�U&q����֠��~�Ӎ7�zc��G�]? ��	�I�����M-1�/����@��������9S�, :�֊[���⧄�z�2��j����7<�~�\�r&F�
Ύ���XBY���{u��{	:�I�դ��G�UX^�Y����`�I�n3��b*F�('�N.$�AJ����`�~Y��A�]��i���цܓc"
_o3N5W@�����L���*h��#�v{���u"�yJà��5qdM;�So��JPԔr�P��Y�[�&�B� 4CxR��<��|F��*��oZ�T+Cu�Tj��a��Ur���D\ۦ��>�i��m�����]�4?���*�/�SI�͎F��6k�9�#/��u��� �ρ�3H��LԆ��Rj�����n��T:�n��C1'���G�Ue�h�*��n�@��ϡ ��?1/�6l�2$�rG����Ȏ�8I����kj�a)S��Uv$��#y�d_��N�(�� ����=�9��"1Y��N�i{$��zÆU'U ��k��8�0�6��Db��)��MW.:�^!�,��]{��KS��lX���-eO��?M4C^��ۮ_�w}o����U�މ������=W���Y7�`F�)��wRQ!4:p���,�?�ȋ��`�В&�:���!�y�藉?%>�u�+o�[]i�S�ȝ�d�cB9N4��	���7�����nw��L</��c�\�+�Pp1�=��M`��yIx�ɾ��$i����K���^V\68wl8WQM
R��I˧��*j��s��#:��!Qq�M(�������F�v�WnV�Rg@Ʒt&������N�f��o���2-]�^*t+!�n��h�h�&�e�0�#գE�9�MX���K�*�{�p8X� ;uE��.5�2���@4&"��W��l%��zw�Ô�2>���5�q?qj���a��^�:�c�-����K*�3,�Ȟ�d���E�ذ~-�(��]� I
�Cib;�i?5U*KBO@��� �ǽ\� �E
�
�H��t���w���喢�倜yo��P<��͖0Z�Q�.��������P���^��](����B�T!T���i��Z�>��W���F���ٴ�z�����no��Q���0���;��g�����?^�Y1��E�u�Ƭ<OR��,��8FŸ]�����"�`#�W�6s�<���Ð��
���(��l0�8�!f�rV���9
I�	�����<��G�h�����v3&��5����=�Em��!T�@�����V���Eﾁ���6��d��/q�Gg2p�t*�6	s�G����F(�a9��M�K�tK(wi���)<��z��$Y��� bfd����rm���d��|�D���d)7�Z���E@�ë)n��.�1�뜲���Z���ݹO�s���䚹pf"��
�˸���֞hɯ�U�fՋ���|���4aM-���*�	�����F����w"%F�馓��Z��v�%^��D!~�Y���m��x-ȣ��Zf-Tj��=Ȓ_Дwu�"���h�h�u����2]-Cm�_3-F����SF�Y�ܖ��ɿ��n�L�QY��|������<�����|cT��y�w� ��9����m�]I�Yz�>"/����(��!}�ߍ3H�t&��e�%ޝ���`D����~���N�ǯ�sabg�	�x@qA3�Ⱥ��� Ź����S��l��A�[׽�{zs���RqF�7��EH�%IX�$d>Sf4XD� w�o�����;M�Oo w��OWN?��%7�wY
��]ش�����<��l1���7��2�_^�ESŝO������j�51�0
�n0;G����ߛm���UpP"K�u�l��51~�LZմ}��T���^���Z�
��Q�7�"m����DWi�i�L��ð�Go� �6t�.�>�d�UN}�u,B��ZK8�)#Ů<��0@�˧�����O
���Z�C�T�e~�X4vt��W=0fĉ���nJ����EDNEy����*��1�fJ���%:������
����`���rA�6��r�h˵��:��[^C�c Wjgɶ
 A~F�����<BZ�m0T���@Dw�0N|,�����<��[0o�!TG~��רn?���$$�����0�)���z=Y�ls��y �JEg-�@\���a�K�ګ�D2cA��7>�"����r79���!�VL�v���1Q�P͎&�OX#�$:�#�i�9?�:��`;�ȝ�.���ZL�V�_��T$�3۸�8���]% �Β�T��z������=\�����OJN]��򽂊�`i��]X��҅
ߔ&�����9$f-�
	!�62����	Ǭ��ۤwФd�43~�V���(PW��ا�:n�n�J�9�Sr�YǕM"nC7 �M!*�ˢ��� 7{[�8���o�Ӟi�Џ�RC�gP�zȤ-��I�CtRMr��M�(�����7���R����0��U���Q5C� ���W|G�����]�G�̂f&���I�g#�^������k��kѐ݇�D�3�(������ۂ!��M&!���(� �|^R�Np��h=JМ�F8xJ��n6�F�{+,�A� 5&���~�4>J��6��d�����
>��Ě,�����6��#�9��1�8��_^w�����sV3��*�����@%�S��� &"6.�,���r9ߜ���-���$���1�����1/�G��X�edU�M�u��X�k	҅��%<���E=���7R��JEz�:�#���h?��F�O�(���%d ȍ�e�`[_a��W=ƽ��j��/�{��cQ���Iv��<4�5i
��&��3��Nҳ)D�E�a5��{mՌ���N�pB$n�4A��3B�0H�7��{���X����\����5��#N��T����׊�"��%����UB(�3��h�
�|��[���.{�*�a&��$���.��҅gBy���dR�*q���%VU��EJn�����U_���d��u�8���R`�'P6�kJ�=�A�RR`�B\DR�䂯[�+ywB�`�Y��铳�a���t�&�C<�aZ�,!��Q���?���@{&�n9��˳��@��vec�(&�=�ޯ���l	����Jh1��A	��$����?�=s��cEgৣ�g��%̰�72�~���q�bvG��<[���� =ҬR9�sY�	~���^���͖��<AQ'r����|�:�_�K���M�J�N�>V)@��\:e�v�ǁ��o�>�h�H:�z��:�hƜ���o�B�CVh��[���n:4�#�eϘ=G��Ո1���H��|�C�3�7�~�����Z���g�;�Ҙ��-0�}�AO��	$�9�xu|���j�~��^�-.��ADI�W�ZL�/7��;���������JT�<���`�\���>�nw�g�G@�z��{��D�!9׌���E�O��%��^92פ�W+!<���f��nB��y#f=+ ׹��_�;�����x6��9rG��#�W����	���B?����Y�篁�S:��wc�ZzU�o
s˒�K�$ۿn��[O�+&u����)�%�>&y�Ɋ@�Gv�핕'�n�=V��b���Cn��-��G2�f
��G��}w���TJ�]�����{]�?�������2a��G4���C��36��sp��8{���#����[���`J[З����t6#Dr���>����;�_���i����躩Dk~#�"���G���"�q������`/m���~[�{�pF�O'�#���/����q�Xw�c�^�\��Y�� 
�o���i�r��U`:]�g0������*�](!y��=A���Q�'3��Jڭ��?��
E1Y��������Q�%s2��솬��v�;t�,�̫ӽh}-�'�'�"���C#���/]�+�^�N��6�U��FmEJi%�x��'�A�'��4R҃�_ch$�G�4�pI�j1ˢɷ���b�\�-�N��xA�5k=��68�Ry�������`\�+L�$�0�dOH!�$��ؙ^ ���1��� �_�)oS�E�h�l��d@��4��yc����7׷&8`ޒ�$E)��g� Yb�_C��w �4`��=��'������&�}}�D�����-�'���l#*����@٫!��
Z��H��k�R{mt��#��"E���Z>?���rg� ��*7��\�pȰ͑�
�� ^�	۸��&^�X�Ztt��D���%�<憎��	D��L�ݶ~�/�B:�_��3	l	��L,J�:'m����IaXI�g]������d�"1R�ՍXK�L2Av+Z� Z��m�~��Fg5Iw��E���{��|�|����Fz��C�ܻ g�]"��>;��]4���YDҔ)�0�\~�T<&�t�َ��E�g��,�]���6�����b��G2	�vk�H�t(m��ܱ!�8�Y�e����~G����4�e҈{^�B8�A~h ��1�NX�\J�q���-08���&m^�!@a�>,nm�<ݤ>�Wj���$�qK���_9���2C����<+�\A�B,��n��5���:4?%�Fo�Q�Z ��eCO�O��F�
v����HY�/��5�Q�S�<��o��s����ΞZ�7F�]\-p�	d���Y��z�v�_{ ֝����g�&?5�>�^r���\����F/ݨD��p��XgQ���ܔi�wn��C�!���������\�/���N�F������|)Y+3�� %k=O8���qq|*��� �.��%�q�y�[k�r�'Ǒ�Р�d��jѥE>�+w�	�V�RRۆ��Nрw��|� �:�vcg�PgZv���3�.�G�0b��$ȭ���� �,eHW&-Y������u�����h�����Fw� ���6�_��W���`�Hh#%���ħpx�0W]�Q+:��hT��w�x���DH2��_[^����!Uq˜�sG{B�5����&1L��qV����U=��'��Р��G��T(��"�J\YZ�9/ZLj�>_�;D��y��W
�^�1w�OO��M�|���{��l���`ci������_�����Ń-���ڨ6*foM�~tD���n��r�O� �PΪ�ڹXx�%;��H�@�x����&D3Լ��0�M��l�n�f���	�u��W�_��cW4���9IO����N��E���I^X�~c �<ǥ��;�U��{uT,cф�f_��f��*�c��;b�¨g <R)��6vg��������⑔q��A|�P$3aN��P�����<�Uڑ�7�jVr�n����tF~_S&Ϛ����V(>_;�~J٫ׂ_1���<�{
��gF��L�x�`���w��OS�
a�nT��XXu�R>����-��+�-DQ��� �������P3��}��Ȃ F���6��������O��c5��JY7�/�T�����|n3�ڇ���V��:r|�8<�ö�6�+�Y_D��8��;S�0�8l���X��� ���	������|/Ht��.�����l�\bI���?/�Q�^�Y�X+�8���2��ݙV�h�, %��
�	�i�m��i�`L��k7S��4�����u���&���38��<����GE^�0��#G��Nx�i ���*������L)oxSG4�N4����S
��N�C����C9@۷ʇ�M����x+�І�CF־���!8;�|"[M	��2����*�u��+� �bQ�:�S+�h��|*��K3I�R<9���w�@�֊+� C��uBw�����x;�lx_���'�	f�~dVQ��bR�+m��;S4�,=�m���5�~J>e�gÔ����~蓭*V6�.��X	ek8C��@D��l�)6�}vQr�M�XT�j�7��|
1H,*b���h}�Cd���
3l9t��>�Xu��=�7��2�3����BVv�Za�.|e�/��W���x��q��P[I�k�nI�7U u�M�M:2�*ZI�l!얧�[�P�2��4GͳJrm�_�Ye�A�8M|Jb�#2�s�+*���t�m��:�vx�*]#Kd�+���u��u��2�2�b��:Is$�*���<��
⒬���s~g��L�P�;�+�G��oQV�(�� �f}�����`,��E����R:�2rJ�H&D�@�_�'������2�$�F��Ÿ3�(!�7 )z�d����t�] "S�θ0CS�y���}=b�O���\� I������uצ؊qY����0��&�;^[����_9�U��F�A��NƸ]�d�a��'h;���p��U���7�׳QQ��x��J(~�ЕڲG�SZ&��Gg�[CҾ�_��G�+~/nx�]���cpTO�|�ﮮ� L8�����+<i�4C�(>�fo�O)�,"hZ	��]X�*�垩&�p�~IٻU���!%�i>GA�u��y7����uq��Ni]�Qz��}ه<����I��'=sjS���]��Hb�����VG�	�����S���S�P��p<N�6�D�3�y֎t"�࢒�P���R/i��}L&O��q�K���0Z]zL�z��e��9x	���l���J�g�/x����JΣ�����3��W���p�@D~��T���so�hyS�����Y��rY�!)��Zb�X�<O ��,^�1l���o���e/Ҕf�K�Y@�k�z�a��-���Xģ��R���**C���Bh7tJ�II�<a��s<����`TNk˂[ ���E)�<v��_����j���K�����%��9����<-W��6�b˼�R��_3ڝ1&��q<������lN� �$RH�x���)�zI�U�a�nصo)��OA����)�5p�Nnv��Xخ��4X�:+�{h۲Om_Sb`���<��g��̀������<��?����a���eՊi�$�˫����K�d�'���;_;��w�M�*�T*C�n���/FP^!1��v����`�R�+�~͆5����Q��vDiJ�<e�=���.�>�FT�������|
��m�3f����`�%۬��[x�E6#���D��TC����Ďºy{�բ0�X�N�}�	��(�C~9s/�/��vYJ��&�iF�9�D68Z|��e�����E#zC/^ֹ�vV�h�+Gy��-1�BZ��yN�;s�;�*�$eX��.�Z�����>r���!p�N��-�n�x�&���F�/vl�pߜB1듓_����w�%��U��~��u����k�~V�W;�d1߽k�Ml��XC٩�=ODw�;� ��UX��`$�h��� ����Q�8���@����p�4�BD�䓽HC^��t0j��������4V�z͛��(1mio4�����ZO�#ne��]�i<C jO+������pzns)Вa�o��2��b��7cW�8����*��"7�]KK��1��DǙ����uPL�(�.�� ��
M�#�~j;�������|Ф2��H����ռ:����Y�˸�-nŘA�ٕ�]؎�^C�<$q�ś����C��T7�R}�Z.µx=N^/U��^�B���|SWs����W�^E9���G�������RT>w���S"�Z����&�v���?�@
ɑ�*�,m�:��֜��:������DEt�9t�ʉߌC���>�_r~�v�o��?7��>��}�����"0�0�Č��m/�K_�����rO����^�P��i�J�^Y��P�'�1�qD��I��T�J���,�3ޅ��*L$��,����6�A��)�#���y��޿UFg��w�����c� s�6	i-�2�#*�M�f �+�����&�E	����$��hW`�j�m9&� M>_��y�*�_�c^(����(8�2rG����bWXҹݔ�����:tx�M��hQ�|CU��]A�*f���z_c�I���wr�Ey�ը�Yt�W���1nY�iEKͯ528�Sb~��G�@׉�u6KF����^��~�ew�
� ��1�c�ϯ���r(* ��n��MG�;aT�5�� 	yk�l׈1� ���Mʧ=l^{<]w��RL
� hW)QMq1`f�D+��^L��5��z(��L��5�	�aᾀS�\3<�h/tft5#�c7q��Aɀq��iJu�ݢ�r��1��t����P# w%�^~ʺ�"w�ϣ灝��k��^���U��F��8d�Q�7t0FJ����k��O����cg/y;�*����Fc��;�}l��>Y�#� ��<�z�1�����L�)�r d�Fn���oHC�ܢ�hr!/@�ݿp7�5��1!�h.��ë���̨�A��Y��TR{*�����)@�p��>��˞�tV��~��D��yif�T����Go"��_{�=L{���� ��~r$Lu�~���1t�vf��R�X�Y�ؙ��,���-�����;H�:,�mgc/�m�d"]�>a��d�F�*���^��k��*�f��V+
�jt��7��뀥E*�Qo�v���Ы�8�|���l�����t3!���[i�Q-;��[��XB��Y]�Itt&U�#�P�6����gFEk�d-I����J��~��Q2��ϊBҚ*�1̿���n"��eX��L��v�׳�Ȥ}��dQ8q��� �&��K���,����0�ʵ��t¦ ��t�7��^��q�j���3��]��a����?����8��hK�sWzG���2�Q����aqjz�|���W�{Q�먂>7��!� ja�|'��u��j����4Mq5�?���1�Q=�׭��d�{{=�sŇ|�%�C�	������������������,� �1i�TAL���¤U��(��,Ejr��4���sc�0"�X�&�-St��[:>o�"�H��ii�	����m7F����'UG�� ��l-!�uӍ�w�����I��;x�0����.T�by?cHA�/���N�ZZ�6���ND�h�S���ʇg��c}�_^����f� ���o�>�Ii"�+��#JMt����R�	ZĘ�����g�:�7>>��G,-���s-~O?_�^%��
=�a�Ѕ'�9|���1_�N�Br��!�_��=*��ޕ2�%��8���這%�N��'t����渆lyR��R�DB��w܆ �@��NG��QY&y�=(ԅ鉌��s�\�� �����HB��E��V�,���#�(�Zĝ4�	V��b?�k��_{�|g���2�R���^���x\EU
�-)����AdXG�۾�c����'d��r�����t������>�Ƹ`J;Tőяy/�6k���Jb�_`��7㦪,�r6#��M�lY%5۪m��qWؘa�G��xWq�I��J� �J�'�f�O]'�/B�ɗ1��G�1��)}���#&c��wh�$�����ON1��-�m�H�$�Ґ�Odђc�˿�LP���൹�D)��.%���2��]9�����Y�2��cQ�Ʉ{���:z�����:k���g)�r��
�F���&�Xj]p�'��N
�dw��)/�λ��-�Ǟd��ER�E1���f�FX�y��g,~�B��s?�,�]�D�E�����k�m�&;��Ff2��;�}vk��x?Y�wrfWF(h�U��j9�vjl�Q��G��`_�b&_�2�?��PM2}4Wd����8%�r2'���W� ��c0=W䔀�e�:��ĂKQb�{�9g�:�ٱ[�.L���"��Ս$+9~��ʛ��R��f7r��s�D���{���y��9q�^^��"}#}�<m6�̰��,�#/A짹3�V�� �"_���u�>�L�4�l��R�!^m�^�W��!�����?tE���Ңcq|ER�Uf�ڿ�'��3�7E�WZ�l���cyE�����J�P��X�:E�{��p~W��G�햑/#d��K\ �{ݡ�m^*�8R�vPk�^�p���]�玑�>Rp�F��+&�FT�;ZFk�ȴ��o6���t���l���� ��\��1+HԺ����rx���1���	3���LO([ӮY������e���UX�AP=��������Z�"2!��[��N�T�E�h6E���p5��uV/�����#Ĺ��RhX���4����r0K�7�I'q��$BS��c9k%�b�R��.68^�뼪֚PL�8���N�� �p$ސ�Y��D���$��=	4$�K~Z�0
�8��b���%���B�҃Y�w�[$��q�]���x^�����d�ŕ�T��[�8�O�Z	�>�m'M�u�$)�
�v�ybb���[v��q�`���UM��d���2imw��A}��!{������bPT	�	?f��q.���W;����5�ޔ/R��҆��_�!Λ�p�|�<�R��mpj�u��[^*s�c��߼1hF���K�hD�q���#(�s�=�������j2�����<��F���}��D㝡J��ͧ��O� �q�7e�OɎz�ۮ�F�a�ۅP�h��^q]�[�%3����/����K��}�M����D�,=��!�!p�Y�h�z�G�0��a���ɜ�UБ�Ӂ�ֿ%㥵�u�\��<�n���\�ь1�[�d�5y2�k{s���s�"�pE�D�6
��mP7��-�U)<��N/��3:E,D���1�rN{D�Y�fK�WJ�~�k�vR�9SJ�|�>*b&K�X�ֽ����$��o6�d8��ыr�������FZص�G����`�}�����3$Eg�E�G�2�Y\ɸPă4*p��h��?$�t���H��Gp+M=�⣖_���-�Z�c��?��?N�= ��	�^xa�:�S`��M̯�qɃ�Pԋ<f�7�k�x�&d��ZC�8y1"n��셌�
�^k��}��y��8>�$`�s��*�N5��q��L8�|<�\�zf`?�S��aEVix&�	@����ٝ�Z<\������К��;{%�I��aK�hW���2��ϥA��?P���MCw�D�N��fq���]�>�&#�M���CU��� �L�G8i��9�p_ʫ���%x�`�i	�a�L����*�������ꞱR�Ë��Fס�!��o������=Q����
X�t�?PN�(�՜Bv3��G��B�d۩,Y�%��_
z<�q��?r#Ep쉎y��x{?L��3����]������bT�wa˪�c�s���+92��-=�C��E�n�
q���m�QڵP���[�Y��^<�?���[!��	$ MCl��,uo&����q��zN<�gt+��;#al����slcw�#K��/�RUZ���Ȝ����o�"{ ,n\�,�wߊ�n��Z'P�
:�H��]��2�@P�s�$�X� �G}�\7i���(��<En~�R~�3�l��X\�L�����Lȳ�+s}W)"�Wڶ��R:w����J�֥1�:i�Ow���Tۂ����K�1cۍDS	����nHr�����K�@<0Oq��xL�B�h.�H\Z��0��"� (.���Æ*�i��4�Ą1~��W�X�K8Î
	HՈJ��=��S�{Q��Ո�jCӇ�Pt��+��M{S��`�?nWO��n�h7�Kߜ���={��GV�pƪH3���mmFŪ̯���-���h|����+���d�:f��iݰ"K��K���C夘í-	�ґPV��)��h7��w����8Ƨ�!���O�<<����B��=�Ƨ�G��d]޿J>�zc ʺ��5�J��zK����F�P94����u�\���: c�"mu�S�]�?z3�3
�f:�gv�?�y��� 1X����!h�!�F�^%#
��F{A������P�U�"��k�nu�Ga���|ɸR��.+r��(A��;�w���,�����ә&�����J���w�1��:���?fr�7��l�2}��{e�;^�x qw�b^��αBe��ZY�s�X��.�18@A~������KV�؇�P�a�eV�������J�LJ����Wa+�Q�5��$�c�+͟?�k0qz���	嶌\쳴i������|�AL�m����6�z�a^O�E�}�X�6��bvL��[��VF���ʀÓG:�?����-�	�;u�W���1Qn��m2�
�נp���S<�hH�Rd2�z��tfq6d&^E��[})}La��,���_��=�49�*�tD�9p�>'G��I���hJ"�����3�a��S]`�mrN7(�{�5;HMs��#���A�qɥ}��͇��!Ym���]%��B�B����X[qwx������.��O�Av
D(Ac`L�m"Mu0�JX���N���g�5{�M,�-�=#:^%����VJ�c{�x˵��V7��V��&�)��4��V�!����pR��kN�oD,k�����7S�P�Z�J��q���|~���l�>}3Z��uv�+��ca�]�m)gj9H�խ� �M�zkT�\�g�ݭ	�x/������A]�#/:s�7�������N�?w�k�yMV5�\�f?1Ź�:}��P�.��(��{�8E}qvt��[I����ˊ�Bq'�	�;���jm]�W/}W�MjG�� 9(�$��>����Q�T4O��fS���ʺlٮc�둧��G�Yʶޤ�QR�gd�<o �C.+���s�n��j�:ddAQf�����_2k�*	;�B �Ԧ�F����d�p2��*{���3	�4��*לsٓ��h1-�9#���f���ɧ�;�6�	n6�^9�{�	Ο5e:a�V�:�D�s����|-�d�����?w���n�m�e*W�d:����
�պ�rh�E,V�;0b���B���َ�Y��
tċK�x�v�������%!������-�cg�'���2Z�C8�h�xܼo˥�b�;>�"ka�0�-��l�N�V.��"
�%�\D�!�6*{��`ޓ�["n 9�-t΍f�#�y^��-Seʇ��~�?�B�9�e`'�'����<��zˣ��!l��_�+�p���VW�1��l����"Z���şd�LG�e@�,ɒˆ�,�[<?�J��'����I�F�-��	��ũ�:����&�2
���3kZ)"&�-���n�E�6%�o�3\���o#$���P�@2C�EU\����zYTA� �9�.�&J�__pN�}��x��M
Wv�f{cݛc5�p�6��� _���q��?��D������'C�8u*��M۲n)������n�/�K�wg<v���|}�*}d�5�:z�yx���i:���*+����3+ݶ�wUj����}p)�����x�7	���C��M�-�o��F�������_1�п�<0.0uvsD���6M#>K#* �P�����U������w]���z깨�`�r���i[D�d1���h�&��E�.��F�5b����Tgݱ��!�=d��O��E2���^�sܞ��N�캍��1�kXy+�)_��z�%�z$���i�� mB�K�ED� ��w����;���[�]h��d���=�{d�WvM\~�7լ�{�I�ýu�ы��SO3{�i�e�����:����$�!�#�� ]�O��zy���Z&�wӽ��덍P���)�d�� �]��R��il�K�̒�rx�7��XC ��j����o���_k:0=2ЊP=��U�t��"f��ro_�Y�+I'v�乲%�WOv`\w�#�Ccv��h�;��'�*$?�el���!�]C����ܫB60K��~L�onT-t���cy���;к����/ئN)�we��6H�^�=��s&�vS~�qD�ڛ_|����W��Q�f�7�^y�}w`��4�E�#��"�i���(�ǒr �Ǘ��ܬ4L�Ė�������:I��m�*ԓf&�CL�]]rE�e|`�(��E��Cݿh�I�W&����Q���0�>��2K�������/-�cb����0P�������?�G|i��3�B��BܜM��<jws���o��.�xg��v��V���o�b��ϬG�9+�j�&B��i�7Uě,|DT+f��~��3z&k���*.<5�>7|�9.d��P��4 ��^��mB���u۩T�����E�t�D�񴝕�F:Q�N�}ZN��o{4����e����ߔ!��*��Y����	Ÿ}n��9bfT#m4�!P��Xb^�Ӧ�ּ�E\�C-��л���5qj�����Y�f����'9�!^���n0��U��+��	��KQ'��pq���S΁����;o�
u�5H�˗�J53��d޶�)��vi��@ �ְ`�nH�J{N���ނ�2���s�������?�zό�z,�o,�7�E3�'�r�����"\0����\xp���Z|����ҏݺ?���/T�3#9��sy�7�zK/3�O���D��/���D�<�&S�����pm�S:��a�+��������9d����f��ĩ^�揥���y!�M��
�=�~VR���OՍ���)�#"�
�3k ����)��h���U����:����Q�$��_�� ���:x��$A�p��=yO�W�o7~G?G>Ԣ�L�bOH�3�5� ��[5�F>JR�em?��q�3�"�T��_潛e4�H C�-�-�+�?��Fp8?�h�Z�� n� o�Xm�};�(*�H��9b����{? [�7pX� =z욛w��5��?%��!��'l�L+�_ߔ�\P��ٲ��r^:��H��L��I����sP�C�uEk�H>��:���̘f��w����.8�WJ&�n���ǚ�Q�-Nu�@;W�Yu;�7���f���v4���pА�]P�ÉO��	��(�A��U�Mii(\���e卋p3� �D����:�~ [W��T	�tIP~��{F3�EA.v��Q��l,x��脌'߻�fQ�L�ȉ0=L�<%���e���qu�b���ǆidh	�7|(���R�T�1ƶ��T��[/�]�a�1���o��k������ͦ^�f���n��O���LI,�w��C�a��d�a��F({�\+\��pұ�c�v���U�=/�B�dHbB�o.��O=�&b��;�_c���5��|LB��*�*��Z'ړ��e�-��	LDq��#�-Т=��8�E����w�p�/���+W���˅U�����<B�R.W�^��H��m���J��g_$@���L��E7]p��z� V`���'��b������<�v��|H'R��N���3���6�I�#�!��C�u�Zޛ	Lr���ݒ���A%4�����:%��k�U�.Jᩱ#�-$'PT|��]�ǜ4�%q��ıf?n�2(t���I	�=�ԕˁI?+�I�2�q4"1��sw�g�w���qȥ_�V�SS/1���`�%�0*��V�2���7e穿��W^��*�r�
��X����B��V9 K>�<qp�d,pI��zf�z3�l�%���(�c���F�{��3s��X+���g(� UX4���JEDH�&�%wu5���\�(X����j� )H�GU�p"�v�xH�Hⷕ����Q�v"Cӻ�ߓ7ʯCn\שߴ�0��.�g}�LS�>�]l��n/���M=���H����3�*T��b�4�ݍ�n��
�J���`�ÝE"ڬ<�9�0F6�\���`{���A/�>�s)�6���n�*��؛�U�\�h�?���U��m�0�ѻ���Z�y,�XL*i�=����ƶ-�8�aj����T�LA�:R��rX{d[֝;�Q�]��	�1�UJK8Ë����o�`[�v�I�W������_�f�|��- �Ҍ�C�WVOq{��x_�&�L�Yf:��*�<�(��l��U�:�F��EM�6���:������ ��I-0�����"��[u�I�5��ѻ���k�9EOɚ�`H�X����>ڈ�H-б�D�ІC����;�@�$W(�38D>��)�(�!�ݾ�6�JL��d��3XQ�˽��(;tb�L�-V��x������g�Zdym�����.q�E���H�������|��I&Z�f�)KF�G}��+�j:����t5\��`DpMLe7��n\���	��x<�7|+i_o�(�ľޯD0����q�'F�Y?�?��&��1���a�)��$����A�]ʏ�Xn�7��N�,��`~F�L-�d�R�g/�p�$7;ApA��*��"W�3芵����{��pO��E>^�IEC�KV�I��Ɋ���>H���>�T�}�� 0~��w�&ñl��U���0)*6���ݯ]`���o�3fqZD�����_/<4J[�<�D�k��ވccȃo��dߥ��\yț}���`����<�k��l"���E|�C��:�s̼;Zt�ȥPf;z��Y�Q���\$��/��V��ʸX�Z9O����w�Xw�f�V���s8>�U�e���*�*����Zځ�� ��?�DV�>��U�0��X��ƩG���Ly�`t��G��
v�������!u�`�����kS�������
�a��m�,��X:��%�-6�-@�6�>�RH}�M�]{����ܺ����d=�ӄ���u.7�u�t�oQ�*˥�!�<���f�hA�rN��A���?���-.5��q8?%l)�S\o��r�$�,�j$�U�� --eR�ٜ>G��?�QMNB��%'���#L�RV��Xe�"o����#�w��]A���4��2��z����E�&�!���N��������� ��6�B�����}��8XGR�h})3�H�k��cy�N����[��j��*L�GG�Pg��J�������c('���۪����z�Eq]��A*n�c��䝌2
;�m����#�'���aH��v^[� �Dvg�'w{s���nW�u��^mw��s�:�r����TEU�����Z���8L=9�k� )mw�b'��>-{����9���ά���PP��2���r)w�Q��.��/!��0��co�w�7�>	b��˳B҉1}��v����͆J�)]m�����Y;�M��'�� �3j�1/^s/x���Z�B�ۀ�0^�L�.]N9<��|��݁t���X��6t�Z��y�b��Hg�Ӣ����l��V�
V�vz�+!}��\�h������2��"'B�8�5�q�Q	�'�nk��#3�>����M�'b�D���~��gr��b���f�PQ���א5jWZY$���u��mTa�C�aAj�mJb��������C���V{�����K���r9zϣ�1�wը�~�gy�����
|��-��h��6c�5�M��[���j����Tj5�>���az&�њhù�>���?��[�.G	>c�\�����)�뷚����`]	�mbH���p9�V��W��1��	�ڪ̈�ɪ	,�_�_�#�sôk���c�l����n>�nR��?�	b��v����a���M�QſRI�������]���0(��_��q�Es���L����`B���Z�C�R68�>D:�7᨜��
��7�`o�*���5\�����<2�g�o�+ Ŀұ`.�[.*���q��������ʆ���iϻ��l@6+D���O���Y�����N�qa�/V��ŏK����+��lU�߱/�98X���(�rP]��9bxx�q}�҆��,����0f^�;�Ѽ��몠�y���B+h�8dmJ�q�����o;�ۑ���͕����Ʃ�'()�D�����/7�/-�}�o�Įy-��sL���eJC0͸TK����R�cY�(�s���yS���Yt *�(x_4��MA�C����wyDc-���px3�������$C�Ax�3����AX���[+:�!�����-�����pv��X�ӊ	��G�hׇJ�
�� 
��"O_���T�t��<k$]����JV�/���8ppA��	��2��5�?x�K������3�(Q����ܪJ
��=�ڰ.�q�0�ߺ�a�X�J� �U6����>l1��ρ<V��(;�%C�1;>>d;zR���0��; ��5X/	�<+��}w��>;����aDgKv	)`k��_8!T�lH�����}�}bul6h
�Y�H7.���%��*��Q���6x��{h��v��U�Z����\f��n���N�񲒰_t��bK+�T��㍋�!��ؗV���!�IU�����vS�L��NH�X�B<��⢚�y����5�8wy�ك2Y���<Gu1e�4�nD��^�
1���nP�
��Q�)n�z�L�-�եi�(�*R��A�j�c�4!-�7G[���~J�ޯ}Xn��D}lZ}_i�@��ɟ�kK���#ja�|F���*׎����F[�(�Y�Y�a�2e Ӭ�$��>�~�ᑑ!�����k/P�M��16$L������ϖ�f��Q��laZ�6"(�W���^����꟤ʛ�t���)�(A��08`8��0&��p�����1�:ͽ�s�8Ձhܪ�y�I�z���wp��ՀU����W�H��Z��tف�-Ѥ\]dR��]l�ڮ��9
�։�+C1Am��E�!p��nNTl��Ņ�d���ꟙ/ww̔�]����9�!�x��%x��İ��&�� �q��[�^C���1�����D�S�0��Y��[��wT,��y��&Hh/m*M����d���6�%z["��k���#r��E���sD4\��9�����>�h��i�	Z�<�#����Ĉ��P�=՞V����`_�YJ�&��	$nD�����	�)=˛��oآ��hr8�HXR���-& h�(�JT�e�ss�w��
��\��`	3l���Z��H�%Lū�c�ߞ��`տ�t���fb-���l���j��u�59�;��j��s�<���ld�g,�kNQ������e7�nZ�e���#�!���.�Q�r�,�_o����ǭL�7�ƭ ;]�=�rMn`�Z7R����np~eɒ����»�z��#����q��3@�.\�6���� w����dy�6-��ŅUE�W�
�׼���8S�XR�Z5H�A��v��Oy;�r&���E��?��7g_�1I��������U��&�R�]��3���|��2:�����$3*�ּ�5Uyێ�Mľ��sL�{bm�ㆣF=��ؾB�ќg�U��\�g׿��V/ݦE=z�<��HW'H8X�a/��	]LP��ro�S߱
����;H��w]�j�H����h���T���Ao?�E�V����Y��[�	���a���e��ȆuO��=�l�ds���iq�X��Jy��;�-����ہ{�ZZ+{*Ǧ�k4���lCFΙ��-<�`Ӊw3!��[c&&�?VGj�?p��Nq�k���v"�ž��8e�2$���Wl��0��*Պ�}�ᡚ1Y�+�p���b6��¾4���r/���1z��pVZAಒ�g���f�C\�)��O��tAWxe�6�
�go���[�G;-i+s���~�`	D�W���,���In~�B�g�1Kx"�[rM��"3����F"9�g�:�5�H��Vy��A��;�n�ˤE����]���뵽�Fn��)�d*S�I�e,@#������,)�}qM���`ѩ�/��j7��	�
��2{�,�0\=���0�&b�=5҂�D7��	��dt�x�;=�t*=`�C~ �x{z��
�b"ٯ��Djq���`���������u"M�`J���b7���Y3��$9HM��|��f#����3 /�_��~��u4EjI��ģuٹܡ��? ����)�O����dL��L��t��%�YR?[�p�Q8�3�O�(��B����O�}�����g���g&�*}dkY���b�'�n�d� we�OZuP�!�Y���%4�qm�H��r1��i^�GB?�n�b�z^2�nHُ���*�M���޼f�7����b��O����f�K	 �-@�NL���s���95��'�o:�f��yg������@�-A�W��z�|�'�n?޵������5��#��}����@�}2`�<�6��jO��=L,;��1ByI��̮p��� _�}S���p@�MM�^�|8fu7��b�#c��T����	��Xb�*������}���y�:��Aᇱ�P��Pl��5������-`���J:�!b���^�B�����(�ϵ�}Z�Y��n"�l��#��, Guȟ�,* �/�+9�5c\NVx��a��ө��n��L�#����w���g�����O����
IeG��W��mah�U�, ��4.@��s1�6���7LoF�6�������6)���,ߐ���LT >u����t3�jǷ ʁ�C�X�5�����U�/�ǶW��ħe~�"9���*��3���M�j����=GI����5�:�7�!L�o�ǴN�wuF- ~�g��~������p��OD5O�I�/Ǘ���J��M���\Xf]���܈�(�eݫ���$��En�I���7>��@�3�p�R&�0N��r��]���ܻjK�]h �� �⬄<@����<��)��X��Zɸ|J�t����to�Vl!�����/}�e�&!�|f�L���ׁ��Rp�F��s�.�M��T:�!{L�N���"�c�7&�Ks��45h�N8jB��~+�ߝ���k�}(�-�F�q�Rs��a��3��>�~�����o����[g�crgu�"����1@m&AZu�qM WӔ�%�f�^�Ks�(a�'+:Ȝx���Gk�xq6�����x{\_y���s�1��E���I��nUK��uF������.ODJ��G�XN��(�L�1�u+�M���TnU�Y-��vp�VKD78sQ�缺���)!�
�Y�
3�ڐR�*ǧ���������)��'�U��*㐌|W:N�ޟMdna�U�F���U���K�f�Z=�7����6�~�2�.x*�	�%��բx���hp��/��R���PfO�7���w)����|�QVĊ����=�o��݂��Y0J���`o�7��X�����^���聸$��]~�WB�����bԡ�_�$)���Ӽ�5�����
�O��G������BL�;{u�Q~�m,�Lt�?��F�+Fꈆ�6J"����W+�H\Zɓ��0P����_̕^iYfԯ���!���af&��D�H�&fl*:=d5�&�"�(è�w���Ξ�-����@��Y��AG���n����S¥$�N�b�[�F��I�=�x�D#Ξ�4��Y��&���Хy��4�Օ�l:n��N2�r¿��8�ݎ�g�!Q��.]AY8+ˡ�����8Y|�'k�N`dr��Z��|Z�����<s�"%��ݒ_V5�˜���_���������������Ϳ�2�vi��>R�%d�|ǟ؍eΌO���SMCΰz� |07O�UE��Ɀ�%����Y���%p��|x]���\�lfʯ�Db(�z��RL�3#�ݓ�n!V�`�j����qxU@�ai��<=tn�}����s�y�һ�FO�JTcx���}�Nw�]e�(�m`�EE��Ű<�/�� ��,w��˲��t��i��^�{̘�F��3v���L αC�Fo9R�gc�,Fާi��L��)잵n�-n=M�f�� �&��<�]T�e'U���ӈD�<��+���\XyR������S!��yrY�J!��{�#� 8��1��#b�!^�&4�T2Rn)A~Pl9�׊]v�4�B2�|�ʡ$��S�n�%��oj�l�L#�*��{�X(��(��Z%����a�i��\��o:�ǫX���������6t>*~Ȯ��[J}m�
V�f��̝<w�m��0��#�$:���_8Uw�'���ҰTk$Bu��݀?���� ŭہC����k^�j�D�Q�WM��F��L����M�Ż.�S����_F�]9-^sm��Y_��4��^��J���Tyt�'':�wە;��~-�`��i���j7�������bמR gh� {W*h'�#̈́+1z��Q�u�`���&	&F�d������0��g�t*�����0�b�!�#�v����f�M� 7b��gh�A���`֩�ɥ&=	R�̶��� �����ܿ�c��g��������7�X�r�jcO�n׈C���c��B�p�a���(��Jg�Y*k-����UQ�ɫ�=�Y�m�+���+�b�]H�#��bY>��*g�����5��P�������m��?�Q;	)�Wk?��0��ƺl�kK��H1Y��)�M�$W�1�< )O/�f�w�D�>xB>b���SV�1�n�
h*߳�f �n��E�w}#���R��(�����^eN�aĂ�թ6!UESE�'�z��iyJWv��h×��T�懇���Wd���/���2���0a��&�k*������tcL��-��eT*� u42�������n}��b#g�(��6�����ѕ�U�2\��q�x��,W-|D��M��D8��Q�W�1���]��)���.��o6���h�!�9���R�S̞X���=��X��Ł����77� �?*(P�!qA ������V����z���a
�PO��?�O�م�k�@����]�5y&=)H�|pp(��=(�c`��I���=�j;8��WU��{S0��Ǻ��[M�ň`�~�9��'Q%E$��3��Lu�7,���&�K=�%�M_&C̄iY�n���g���[?�,�|]���*[�҃]ș�#g-�����`Tx�[�s�kD3����`����9���I84���!4F�jqVy?���U���@��.��3j����7��ϋ�meԈ��t�V	�(s�e�
��az�DIF�P͛�&(�ݺ���Ѧ;e)�����	i�Mr�(��5�雝�� g�2�Nw�d�� �!���)�^�yU�94/c?�2���U?���\�D�yse�2��F�( S��:m�"_���h9P��R�>�A�����'�]Ѯ+�`<9���ACv�~wx�e�'��8���$m��Ή��R�C�ЍP�ZNn��6N�^l�9����@`@�OQ}����X� ��D�=i
]� ,�v��V�/"�h���@)5P-ը>-2�Z�Ͼ�:�Cs�;Y�$���#'�y��/91��L�f5Nթiy����ǆ��#���,#e��"$�n"59HDs:����Ʝ#�o˖�`��������5R�&D8�T�#R8���V!� �;|C�P��݁>�3&����k� ��o��QP�7��0����m>�����[)����1,��
������J��*ͽ	�S[����7�-�ɑ�Z�`��*�#V1��B���w��	�(i�3�I¿���*�q�"���I��0����(R #c~`P�4$��7�MFB,�G�X��f�T�k�������E/�G�&�����T����nP��A���|v�L�duE(�O��u��|ٌ:,Ȱ��g;�m��zټ@�Ķ�F��a�Mk	��??K��ǆ����kcw��ɕ_��]�Ԛ]����Qݹ�θ~L�r�.M+����2F�5�O����K�F�РdQ�N$<���-��ނ�<����-;��XЩ�5H��s!PO��(���
���^b�p� �"�\8�r�h�诈�k�W,���,����?�7�9*Z�4��p�	�d�'�&�˷Xחɳ�(,�~]�}=Yѱ;<�֠�H���d�j�򞂫������^Z6"vX#C?�r�}7`*��v�󠏤�ϼ��!1�S�	'�D�_0��-�$�my��a6������&U&#��Ӿ�þJɏT6ڛ&��i챰�v&�Ŏ�;F�@ӽS�1��������̳�eL�C���{R9|���O`A�gf�cRIf�	��E��U����KD���p�&ZkT�p<<���hJ�U1XX��W��l�r0AF�$�׎�U�k�;�A(�5�i٫�R.�6X�>�������_��^�z�B'��t��?1"\)^�?�,��L�❻/X����ވ�n��F�"8�d\X��d뗿��p��=�ZP$�z��!q�Q�t`@y(�bp)	�&tt�-�+ⵄ/�o�+�6�v��v�ۑ<h��/_nGm�d��lέ
��GfOD�c�+�)�t�ֆ-j���:GR�qS��W����5]�O���0���Ҋ��-g�G��H4�R�&��i3mS�2V"�A2��	��ਚ�m7��lϱ¼g������O��b�������?Jg`z�~9E�L�4B��C7���ö4�����y�z��x'�cW	7�]�[s^�(����xV�	������# ���o@JѨ+�͂{6R��r����ɟ��*��Q�.�'�F1_#wc=#,��f^��&,�������ߘ}�?x��'��6"��GW?�&g��,�g5	L�T��~�!燛5��=��"�
u�h�P]~��d1	�<�Z�q�('Ic@&qDD'��}�U�,	������I�N;*��WE:�J?Xfk�*�g������K~ �f��G��K���L6`-�������0�܁+��Sܢrӝ���(��O���:Һ*t���U��O��Cp�J�G�F�6]ZbZ��WC��@���ΐ���8/�Z@��ޖ������_��+�\��� ��(|�fIʛ��h� ׆���fn��㑃���^�ô���F_�����-��-��x��m ��Q����+�@2縃�
�=�U��=��N-��w"j�.B�3���h�m��O6��١�E�l�B�16O�r%%b�f1���+��`�����d
�Q�$n5����"aD�¬��ÜJ%�WN���gWT���K�������Nz��|�)-�Cn��:��@ĵR��>�[#��n��W{����2��j�0���1�ൾ0Y+LUݨ��^U떊�f8dT8z�w��� �^�[�EO��"�Z�3�V�Y��@������)�5��"������v����,vtjR'07� !�e ���3S��
-�#�>'t#I%E�h��u�o��E�0�^-��1Dm�vq�D$����9g�@�ʔ!q�P4i��[lL3`�x�QJ�Z���.�)�֨ԅ����Ѵ���c��Ã�{�'|�
��p3��n�����`0�aF8BQ��n����:���T�\E���HH{���v����u+������C� ��<<��G��n7��7�3m������� ��p�=���-�@�Uq�y�`btQ�
y���ˇ�}E,����FK��{��)˿@�N,�������"E�g�v�*��n����:P��ƭw1ZL�p=�e6�4�����73~�A��ޗ\��VZ�j'8���'!&�9'�Gm�_��T9�i5��R��a��c�J$Z�oQGE�q�//�y��Gk���bJ^\�X���H��F	O�J�	Ѭ�:��B��8V�(�D�Tv��?Dg�'�t�����l�]`&�m�?�zܸ�z��UD	��aCxڏ5�x�󀙸�v؏M
(m�4OKxc��;X�����ChˎJ:�]��T���L�۷F�~�ض���6z%az��"��@ZXc8�J�=l��2���~�,�c���{�ͬ�ޜ^�1w�.w��1W��>��<�S�
y!�9���f[:"��B6��{�|h-"�α��#$�8��t��ciY�*�=��m����ź5�ح"Z�)B�BR��,�b\V���a�*��S�תԾ�u��+T�̟�q� ���4X�ps�#-��=��W��8M��dnI|�)ܤ-|�/}A��L���0�É��
2v�;�"'Aw��o���	>/��|_Rw\����};����4�V7�$�)�/��,@����o��Ӯ�(��yv7��X>�*y��/�m�>����,)_��������%��22�⏈�c��4�%(�3�w;�W�l��B�����Mv�m���4�=�D�D_�2˹~n��:ګƷ*�ᰢrB�ܤ��材���c�[tQs)&�a4�R��X=�2~�����v'�\��r@.�},h����|<����J
�X��q+�jD�V�n�yu�{��s�Gp�h���V�fЃ��f���E^�?��S��=�������ԒV�g�>�P\�t�d��^:oZ�/a�Z2P˕s�A����V��(��&� ���S��
���&b��x(�$�2�w���t����M�* ϱ�ٕ>�j��Dy��MG_���k�Խj�q�c�N��U��ƚ^�����W��7�G��%hQ�X淡�"\ys�bN�H�|}zb��>�EE�T%i	S��04�O��>7Z�"�.�ޱs��-Qã���(�U���ʯ�<��=��E�[j��`fe�C3<��;�欞82�O�ճ�ޱ�3��`M9�Q��Ǉ?�T����UB`'�sf�Hr����EK]��\�VC�m���2����MS��Q]$ǥz0���H
�ܭ�=5B�2����N�+wy4��{S'\)�!����7f�F�ꕐ1� �T���ŲNHXA�.1m��<m �L�N��zI�-i�TC#�$1?Bs��=$"��󍸓%/D
�b̌����uN&��t`��wi*���o�6�R߀ ��[�.�)�����M�cA��rm�����ڏ���N8�Q\nw���I��˜�b�u�_�y��+3O�����^�ު����:~�\�������F��:��.mԤ��Ef�����
q��>Hn��L�oP���u�LTZ-�_aw2p�����[�����;��{���	8T�\��(��X���C���WbM�D�"�X�9�[K� � a�#tf���-e*���D��o	��_CI�
{��k56�~��'ī����f�Q�C#G�7jU�6���M_>@�������`��9*�����Ԩ:o����̜���,�[}N���8К����a�<S�E�&���Q���>�&���?����j��2`a�d�C2����(�7����ǃH�YkAY;�W)����4�%�.wm�4�j�Z�,%A2W��$��Z_Y�㐎� ���gnf�w�̡]��dh�ʯ��zP5Y�H�0�5sGl��m�LMg̑+q�(�B������V���AdRxl�y�ۆ&x����ٹ���Hk2�h���	�%XT~�M���mp9f�L�"&!O�wϓ$� ��I�c��k�9EX;DIHmZp�g��R��яS1nC����.��Oz�F���)�t�񶅉M�h�$`�ˎ~|����58��5A�"�օ~̥z��gV�xރ��CV�K��N�����X"	F��0�~�cmr�)���s�s��V)}�ι;�H�Ҕ����W�z��T�����\(�"R ����j��G)��]u�!�{�r�����$E�Q��Ztq��MF�*�[��-�;���n#�g��-L�ԣ�q!x��5g���*h!�{a4�dce��q��lqk�A�O���X%�R)�n`f;�-Rх^���ڴ!����]7f�$=�#�p4Y'n
c����O���r~�J��ʧ��f�g�����k�� �<4��4�"�
�Z�����H/�r0{�	(�y���A��� �,%&��q����H��lpn�Z�D��e����A�R��,9L߄y �QP��0f�+<����6_���o�<�2���b1$n3�F J`�ft$e�I��S�|2A@�g�:+�n�;m���/9�T�)�L'��!�(��S`2_b&*�| .
UAY�h#t�Rg��m�?��W�y���6����M���_��4BXf2��
�z�c��-�X����;���W�[�3��5���aC���6_��������a	�i�r|I'�}�aNWѕlIw��&�B	(kh�����9��MM���'�S���د�-I�����ﱭ�7T̈t�����*�S88���6|Ȇ6=�H�ɾL_�h+O�ٹp�O^[�T�5��D�
��>ַB� ~3�3���T, aZ�b�#�(1����j����,8���j�rH?д.���:�YqS�f���;n���)m���'A�y�$f�u�?��8�m�k�!������G��ꆃ��� �����7J��R��\�J��5U���%X�^�y`H��w�/!��r��J'��ֽ�iSh bi:
�^�	�a�q��m'�-� g�,v[<"WA�sJ��ri0ohl�o�P;j�.l�sI�KG�&bs�!m����e��V��~��7\�H�e� �ց����>�RЫ>�������E�>�f8s����!��5F�	JF�ʮ�o�"��ߛ�A�����.ת��Us�c��LE��q쐸���������?Z7�� ������7$?�kP���-���``��t3�G\�A�8����}�<;| �������5� h���%���Sr�;�\7I���Oͻ�l��'��~��3J�%j�C�����U�e�`�#{�u��-�0fY�4�y�����橼����|R�����H�b��9+��{n�g߁���{"��~��j��1o�s%��WA�V�zLwМ/�<�K�@����d����V�t:��^㥧�\�Xʶ�������|���`���� =���4���sws�>���q�$�n����P���q��w�,g1̋���,�����rP��׸@[��r��p6�V4�fI"�:Y9u��(U4z�+�StR�9�N��a�6C�G�x��~�&&��G����,f`<�;�n�$ CC����m��e�[���ڀ"������Q		�b�PR~Oޝ/���3�1�pԃN����^A{�*��0�*�c@X�N�Ω���מh]�AE�j�W��a������2:�M�Q��y�uY˿�{S�v� G+��p�9���g�5�@�����4�5 #��^�/>�9!r9l\U8����e�_���VI%���>雐�$?��nˋW�YXa!�T,��l�<%,˵�(y27�?4�,����4u|o���%�l�SҶ�5�N����`|��U;����.rN=�	�	?2�PyH;/p�v�Of>�����������5��"+~�:^����=J�}`KZ��z}e��<!Ng����E�k7�fͫ��xa�u��:C&��L�%be��#��E�H�^EdxJD��CNAN�����C-��Y�I�:��O�i�Yӧ��������ߠ�l+��uU�Ϯ^�*&�!�"�`3l���Q�����c�`,&����*�٠�c�9�~ze���Ed_��ψ����d�JR~F59)�EY�y�����%9�PX1��Z�3�:�$(���Ww��c�$��l��S<���PF���)]�H	�� �i-��n2�4��9�ǣ��� �X�-�f�p���yo���	������PQT`�-^��i���/�����f32�=�U� ;fT�+t���ҥ�8��sX��2,3�` o�u��@P^���
�w���ٵ`B��_ˋ��s������S-BR0Ԭ�]��d�cG|�8��S�1�x�5:��s3�F�:m��w̸1��Gf�F��`vV�m~G��r
`�Li��A_/M����g],��y�yP�_f���
�k�� ���qMHN��u����ĉI�M��Z�++��Cʸ����]����rc�)I����6�;I�=��4�!>ڣ�t��"�������dmWpr,��'ͭ�Z7���IV�I��d��-�b��;��!��������O,�.g?�O��X�+�vDF�B΁��f<�,bIy/�* ��M6�U��K��_��֤���m�}گ_�FVI�Ih�%���]�ŏSd8Qi�-xI_HT�@��WVh�/�ɉ�KЏ9%9I��$@q-Q�,I�I�e4-Q�<�&�M�#IXZ!�N�Q�)Q,�:,@��,��!�������/ ����@i�0�v��!����ecc�Q��B��3d7�~�ڸ�hrM���UK��~��`��C�a,0�����v,�}v�~x$pY�|��Ұ�Q�(K�r��	����Ө���R+i���S"�����n��9�r��cҋ~A+k�NA���yџ8}C-38�<�������C��`C�Y韢LÄ�u4y Lv &���(��U��zl��*����\��)W�,j�������I�~ռ^�5z���;R.�l@��y"��s�\\b�!ѫZb��q���C\����R�K6�19DIcۚ���P]����72LpkY�ǔ�y?w+�\^�d�(�oB�ĔJ�fu^����6T������;z�����T�h���U�@��T=�Q���"�G|���U!=x���u�����!�����Q������xB3'o�����a|�LG$�^���qP�
�b��.@}��VNͶR��ŀLq��o�qu��Ȅ�,C�l&��0�ar�|K�d�������ͣl�2�JPN��N����[���W�kYkt;^nV�v_��:M���(j1��i�HV�'���[y��2V�ԭ�2�>?Q��aA����,�{"m\Oґ]u����3Ӈe�\޻a���~%
���(�bR�q?�u1�`�C�h5FGW��?BVD��_'-R!�[�{��K���SS��?�5�L��l�]����<	 :űE8��M(���x,�m{5���`r�q<�a\�%]��t��a=o������et�����n��as��܉����,���A����ķ����ў��U8�lR��Qt)e�+ݡ���WLG䩈���a�ogf�X����"-����,����Q��\R�`��mEF�s$�P@�z�2����S�˄�d���ۍȀ��T���� �&��d�<��H�Zw1����`��;x�m�cq7u=:]��Y������t��f��4���Ӷ˛kF����C��W	���v��HdV0v\p�;6�d��F�Մ�1�_)T�n�سt��۠��߫y����Ô�-��}U&�獳�M�����vg���>��f��S�d1 7�S�cE�su�=�Tݻ�&)S˥�&.�?�z�WB�K�S	�5�V�ʽ!pF�}wU�����u��A�\�_��h�C����g�
`}]���!}�`ZBaݮ���'�y4\�0G���� �_ ih�Ϩ�!i��������#�m�'Bes��#8v�Ǡ�����m�mQd嫧!��k� �E����y]L�����˕��K��;F���`��u	J6:T���cڿg�������ot�+��=�ף-�"B�B� �ϰ�--���` F'̕L Z��O#��5��~�:�R�e��Y��R�5�߹�z�8.�]?�v��� �|�(�	�O��?�<c���c��Ѿ3j8�q�e�f3��t���&��8��g*��Y9P�nħ�f�p��y�=��^KӐT�?���W���N���4�� +��j��{�U�s'�.~�;-r
�x�q�N����'_�Q�mg���aq��٠���_�^r�6L�跳�[T�N�IH��������� ���AG�����=�5WK��j�&kIK�A���?}�6ė���P�n���]@F�dJ!����QU��/�Q��Uw���V��\V]_˄?�Y<H����I��&(|H=R�,�s4�����T�_��v ��T:U�=��;��m�=�>;�����
��F�J��s��l#,����b#$�M#S8}bp��i�ř(b�D�1&�K�#��1��D�{Fnx>�Q��KO�/��f�7�V�JSbٕ���V���}z@�֡�!৲��ԅ�!<\X�&~��R!�,�\��\k���~��}}g4��i{�mlD��Mʲ��b83 xG�JsY������yr�fMz�Ga���J���J�D𰺳�9ũ�+��Q={8�����w���� ���X;����7�H���灊b�]�'s#�9_:d�)d�l�.ڑ֪΋�X����qￗ;�rٴ~"�(e9
��3�,����7B!V��3�xڿ�a��r8\��"	�R S��NR����k�琎���@4-�f��x�e��ޚ���ۛI^�߲r�`��a��H`V��P�Dr�Щ:`L����g�w�tW��5�N�(��	�L��q��mܭ�� ����QW��Y﵎��`���}԰)�l<���E�T�g��	mk�hN�� 9�T�I�F|hEj�[ѫ�n0�'�D�~��ߒ�@qX�;�H���6d��`�6^��y,V�V����E��rt��O����g*��U����X�kڱJ�	-a&�y��5:]G���(�s���-��ևW,!��K[�_�?��O5C��,�&����F�q���OQ�q: V�����C���40��y ��0z�S�KE��O��6�'�+ch��פu2����L8��h�;ף��1�������_�7z<�ûm܀�i�Ȫm9j̑Z�ù�aj�� -â��T�RW�r��b��mQYe1��bҥB�tD9�ϑ����,K�M��s%�l1]T��\`HN�U�QT��w���L�v+�m��(}�yW��[�����>�����˷ކY����e�Y�%ϔ�ő��-ʷ&d*�=�$�³�r�O�aF�=-+��)�Jo}�u�q��(ġ���l��7�b:�����|�t����!�Q���d��i��H���Uk>屧ʴ��v��zz�5$�q��UwD��beM�--���xOU6�'LXZ9����&�tpEC�b��i�ie���k�Po�ߨTI�d�|)�HT�m`^����O����:�A�Q�?W�^����S�J:=`�]'�N�G^��e���B,U�\���-�H��8T�J��N�o|_10�0�#\�<�*h���k�8Y=k�z��?zN����6���l�P��4�An�r	���i��H|���0͘�*kPs1���w`�jj��y���
ܖqŘe��5l�B֪�u�?m��w8f�T��W��N��c���*�Xc]#�^�@+�T���OU9(�\��D�h��X��Ev���P1x�Rї�̀:%I� �/2�:\.��i�'�j�7Q/��Q�N�$d����n{uL������5:�,L��뱑1�}�u���97��Sb�2î_G)O=�3)���B��$J`��c�C�h&�$&���Cs�gL"y�|�-K�$L��$����O�k��ى��<FgE&%�$����6�O�_iev���h�D(r臤h��7y��&����9� 'x��}.M����#_B40��P�J�G���m��'*�1g��;a�v ���׎�S�?�l9��Jt���X_�>�M�d�����P����͚d�T:EKh�~+�,Gc���!e�8��
��y���F�� ,�M�4���u�-dȕ���O9���(�ǅ�k#�.���у,eyEu��N8$�1 �gJ�ǰy7��a�p��y�JP��e析9�G�"N�h~y�mY�ώ�� dӸ��w>{��_�ƶy�<���j�
�����hBY�12��G��������JU�.g�f�Q��ă���B���IgP�:v��5U��  N\���=����rZJ��Of�L�~�=�9Ӓ�!a�k�d�*qTG��R�+�#Io����I�R��#f�Tg��>��]m|*W5tC�\��wf)ߟ�L:wy��:J/r\P�	�a����A�����j�Z���ɥ�H6j��7.eR1�r�oK�0�Lxj`э������Y(n.=�a�.��}B��E>��)���ޓN��N������s��L����ӹ�9�,i��s��y���B��j�rT�IR�sM��T�6 �����*��A�����D/UV���JNɦ�ߡ���<'�A�14~i�&A�woe�j��Ȑ��$�S�����LH%,3�Y����]1k������b4��qV�i)��[��*�I�b�Ua���Ƙ"4���p����Q��U����k�AE���술���H�kg��h)����Qko_Gëaˤ[+a����O���$��F��mɾO���<�J��=J�Hk~�"��+�^��;��U�?�?����5I�ŌU�̾�s7p��a�0�7V�˅8�@C��/-jm����!|��ilg잼��h�ɦ����ȥ�k;�`I�� �N7x�����.��_��(q�u~g� ��J*A�w�G�d�O�ĺ�WT��;U���[9M��D����fҶ�&�%S�ǎh?&Y�bC�{.W3��g�]�h���q��H�a��ju&d�-
���F ��FL�����R�u��臔��u@�$�("��!8�L���%J�W��W� ���=4���P#�c9Z��N�ʧm/��V��s51ǐ{����Ĕ��@]�wY��v]��%�
�����]k`J~�A��L�e
�=�;N���u�l�"=�eT龇C�稌�������mKಖ���p�`�o�k{����}k�uj1!�
�6���B�����)��R<���K���'���Խy�P�0�FgKGs��ö��}ŝO�Й��h�aV��ǖ �X{��87�'^�}��J��pd��7�ތHbRϺp����@ 5��덚�"��K�K$2�#�4���k���E�����W�mP������k�9��&�p�n�l6�|#0�'�Mi�,k��+&��h5%�[@ݽ�Փ�x\9~����/܋�����x�AiR�b�jڼ��d<��>gW@�ȹ�svg�j�O�;Vq�(
��
!����&�@�y�3��K�{�E�N=�*�hV�a�U���G�� �B2�E��_��s.���)&�y֒AI��<�՟�>T!@�Ԗ�l|��J����#~	�p�k�'%HN�\'����V�қߟ��g9dZ�GjV���wo����m�R���p�|_�.;ËOz�]-���]����o{W&.�mn�����im�����iz�	9j>�bK�D�L��!�`~����V56�3��A�lݰ#�+����A�)ed�7;�h�0���4y�
{�`��+W;�d	�D��_�}<r�1u�՘"A2Re
��������#{�fg��M�8.ka5�z3*�
��H8M �:�c�c!_���vk��T���3�gn�6~�U�IStRD����N�})�N񇁡�= <��u��m�;�����_�6F����O�c��`�LL�.���_��������UG=��uö��d��A��mQ�ZVri���W�̹��RD-����^8Rո%������7��Y�(*Syu���H��/ԗ��܉��{3vn56�BFg���bN��&H0vpMaCh�.�F0�ݷ��Q%��F�؟v�W���Maw��7��:��B�]�B�>G51VB�Jҭ"�>Ҿ̙���"���m�Q��ص=.2n��aQ�Z�*�m���H'"kZ�\��UqII�����(�«@?f'J��K�D�Z*�����<��D��i�A�8���^��ᴸ���/2d q�k����姙�{�rX�v��S$��4�U�k�]+�����:).�!�&����i�8٘r���ؚ���P+Nɖ�!k�Ö��Gǚ�y�z4M�Zhp%:t�q�e3�� o+F�{�i�>�Y���S�)z=m�2s�Ew�l�|n���hp,�>	-��6ω�.��r�
�H�Tg�Gy��&T����� �^(��2.���YZ�UM���4b�����ٴKsOJ9��:��>�IF_Ĕ��*��q䦀:�́5��ƨ'̌����'������7����<���Ⱥ�C�ý�����k��1�=�?�U7��v��$E��͏����wV�����>���E�d;��]�xO���Ǡk�8�0n8�H�O`�n�����'Q�{���˺/}���O�q��ON��A�g�yߔ��N|��c�X��tt��M-�k:R,k����^<)���4{�0�Ȱ�w]G���	{�PЉM�>ư�	����<9,��Z�DL�}�W.���e0��l2��;��$Ԗ%�H�
�X+��k�jB?��(Q�Q�%+�Z�ʺ�?B��G�(�����]�T�^�z~X��n޿��j�q! ���P������l(Z1͘�ݫ]B�|�/��J1KQO��ЇpG���v���r��(��
�~��K���>���!'��R�QG�l�PsGm���2��H&w쿽�/���lpB] 6���%����`")������!����
{?���ܜ�x!��L�!�H�|q��^E��p\*&�q�5�5�����[s��+M* z��N7P��6�+G�A��Xb��Q/��C�Q��#�
�hu1;�Է��yR��/)C��:Hj2v	=*�k���x��}y�E����lw�����&!�)����C~Y�-]�szW�N|���Q�ԙ��ڳ��_�x٫�x$�\iE�Srh���o4�ܳB�7O@�0�Q�9����89Yo����Hf���V`���4����k�{cN���w�TX������qs�����Q�x^h|�$�L�zNF��2��nD�I/�����vF <b�P���uC����`��}�n�^��O�f'����H_�<�PI;�RP�8�� J.��[�<L�Q�� ���`-·��daq�@EEヾԵ���~���h%)��=c�@�E�$�
�Y"X��Ǌ�qלzÕ�� ���Ɯ��ndӌ�t`�d�L�
ZP��/�����tŤH3%�uٳ ] KO�I �
:^Ă� �R�c�8��5�BZh|�YM�%kkM0JI�r�Iw F��ͦ�J�2�f0�ZȐ��*��k1XQwq˸@"�-�Y��O����ݣ�	���ݔrSb9-����>SB���N����V++g���<Z-y�'MxۄF��|�|��(�Ŝlp�#� G��ٟ�5T7��k�y) ��3 4d�%�S��؀�͜�<�� +�R��o:ER�j��ɜ6�+�$8W^̲�2����7w��
�Eڛ��=ȊʡaA��-�[�G�|�k3k���]b����/� �xS?g��Wc�)m���J��`V����1�g�š�+/�.I�1F��I�Vn�qS\?����ߊ���~؀�K�ĝ���B���0�l�o��В�'E'^Yu�>��W�d�e>�̄�h+|w���
b���z{	qTx��	����=�h�DX\�z؍d��C�a%W3j���&��4�x��[��,݇M��5@
�2	���ő����f��ޠ�����J�ֽ���	$����5��h��a�� �ħ
�y4�����,ϨP��T[60�[6rj �}�l�,Af&�$o.(�?xl����{3@�"R���LC�:p�"K�ciЛHk�<�:\\�B�:ύ���d�c����[!3�	8��Y��,5���?n1l�w�ZRv�uE�?��w#���	ǹĽ�1چ��xL�fSы���,���1�D� ����	��}���f����n��^[cxU��~�|�Pw�z�w|-��DP��(r26���  �k��U�|-�]f�o�������^8C�g�p`���E��x-4���1�hBئ�U��`5� o��=�C<��$�Q���-pR��s�m��Q1����6��Hؼ|���:��$d�_�ϗj x�Fr�qS|M��`Z�Q���Oc^�4g՗%��p�Ϸ*d#��� &l�L�\:9���Q]���(������ʙ����^�VOh豄z�|�t+��(/r<t!a\�pI;�@��4����̯ĒB�#d}�bHnf�@�{xQA���.x�j��	o�%���Eav~�.zŁy.��ώ��s�N1��QH���<��DG�n��_�� *��̆xO*�L6(H�P���vdTU�K5U2	���9se����bō�8{������f����"��E�����EK��bz�������k��li�c���-8̻1F�du_H<��UN�Lp��G?b����`8�Tݱ3�J/;A����w�S���)/�u�18.
�� *����_ZEz�픧	�+�\��;�4�%}m�8���ya}2�4l	��5�V�\�?�5N�DfQ+9ߥؘޑ�t�lt��ۦ ��5=V,�X�� Sе�O.Po�\�H�7 �q����4��x<��t�z؅O�!%�Wo(�<KO?���^h<6�MN8�U��64��0�N�>�y�JS�����ʷ�6�8J/�HZ�F����W�5ʚ{�w�q�/B�\,AY{%N���G�I+*15���ro_�ܧ"M�_�uw!y�.�_R��	@��=O�3{�\�r���TD��M ӵ��#�Aa;E�y:�3�\��Ӳ���[]����Yk�d3a�y�k��>�� Wd�͢�W�Ja���OK��P��Hh�7�rF��'��$s��L�*bG~b���[N�U܄ҡ���cGh��f�u�o�4�=@�id�2�vRU6ҽ��G�Q�"��T�V�x����/X���;�2e7Ĺ�5��#�P���,t'�p1��	�S��_��`t����SX�ho)��{����N��{�������C�);D!S�E�C��Ԧ�E�)�=�@���3=Ri�1] �R�\�o��p�7�r��rD��gS�D�z���G�r��(��䩺j����F{��JU��=��t7s� �8v��� 7��0��D�n��p@yq�1�B{��H
�k7���2b�Q<��k:]�{��i��6�v�ےE���/R������=�����(Ԟ��M�vnC�O��H���SǄ^�\�;U�	��x�ux/��kM7t O�z��7� ��������:K8{�ظB�^�KS�۹"����7$٠܈*��a=U�W	@ٹ�̈ֆې��A2a���H-i�=�>��'�k���)��
;J��#�{mt��0�?l+^�:���nh#���SV��;E+�3Ɛ4��w����Pn����8���z)�-��Lău%�6;�Ε��O����WR�N��v�1:*]F�F,�g+���k
�����åƑ�A[��J�ī/�
>��C��d��P����k]��k?~�?�^�r�fS�bm��j����1@=f-3��YV���7�כI�o)v�p��8�o�Z��[��w�a�W�3r}��.N��E:�������=֡�!�#�R{�}�J^_E����,OQ�O�_�'�R����J"//�jp��j�*��f�[Oݙ�70�����{���<	?�5a��n�/B�a�������@��	��i�X���Q��7�%c�������YS�F����M���H����'�s��lMf�7f\�N��L�A�G
O�d ��:���1��YK{��G]J8����X�K�3�(�@�l��Z�0O/���'�C+�zG��C�����m�ȫ��>��Ll]���#�,!�P;�����ŹD�rVf���Ck˾B$Y�̑��}L�ͪzAn<��+v���\� 6Y���DZSPX�IJ4�c�R�-C��q�`uӟF I�� �L��v��8�y �)Sy�^�(���Z$�n�0!���ڧwʪT�u!w�����$s���2g`�!�<|9���A���B�q�OEI���Bԫ���$89�M�n�����|헜q���O�4��RE.�C�ɪc�f?��;R�F@F���}L-�T���g{
������#�Lv?j��ߐS�K�s+�{`M7h�-�nu���K~��xC@�PG�nRӎ��,�h�'=O��c�i�����}��&�a������S� ��� �=�_pR
3�����jyۧ�W>��?;��6�u�=���]t�f6���HYYn�2�F����#�O�Si^��bo��r�h�c��X1b~1]��k�}PؘL���S$�m���P{��J�_6d�欔
��7�C�r�b��s���B��y�q��g��е>�SV<O��!�&�p���KM�Wɺ���E��ɁF?F	������4Z�6v#2Y���;�Fk@ʋ��\���>[`uM�dA�_���p,
kt|�U����E�4F�|,������Oq-�����2�,B�;��Ùx\6B�A8Ҕc!�	ǫ�yR��gp��W��K������8?r��Z����7��W����yk�K5߾L��������3����<�a�:Hh��Y:�/[��X�{h1>�H^hs���+_A�j����[Gro7���E	�m�|1\��Dm�0�0�:��,�K+ G���G lX0�oZ5�����U&5��v`�MA�v�  �&��a��V,@v
ƿ? ��Qr�ʃp�0�������-��̕ွwG3R6�$�WS%��&K̷�Sx���9��^�g�&�.��r�ӧUf0�����I��?�dU��*�0�ڀ�1�`H��bVP��~5u�����m�����Qˍ� r���Ŋ� ��GjSHk$Yw@g�~�i�q[��|É�N�P�d:?
&��j�ɀ q����Da��³ǣ�G�sr�>�H%��ߴ��e͆�Z|���h�le �y��|w�#�X�v;.sԆ��n�O�|_���8��i{���Ip��M�xֈ�6���@�~�F/Jew�	�F�&E��yl2d�)��Añ2��!K[�'i��7�)�xx�m/�l�ч����{B��*�4�soP�k*pP>'ԉ�����~��6�m�3U�Ԃ6��_(j�lV&f��q�F��Kt����är.�x�ݞ9��jm�'���8W�7Y��ʎ_#�ͩm$�P۔SR�i��]M+��^�;�s����+y.V�~��n�yM\ς< �d�A{v��5�&�U:�M�	4�� �4b�K:�~`_�;Y��]H���'��ݹ�P�Zu�/�00�2�\(x�d��3�P||ƕv�aɁY䎶GReJ�	�@�j��p`�H�v%�d�R���m�8:g��D]>/d��ݥ]³7�xq��
�j������t<�EZ��Iu��ej��B����������J�+K���rΙ�f̊��='�a]8j�.T��L=l�?`�>�כ�Zg�$�_���nu���.��|�uǚ;�u�1��c��ʱv���� �ϗ͠�"�6@�������ˁ��6������R�	�^Dq/Leț�+Şs#r�,�g���@}�-' ����%���S���%�M\|��V����W�N��,a�#P��ЏRt5��`���ۖ/�=��ʋ�M�Y@��f`�zSࣸ�PYÀ=J6$^l�@A�f��c3_kJٖ�����|�i��h�&g������V�y�r,�����?ۊ�z�xK�4�Jo�e�c���װ��hW9�[*a�#8��+h(�}���LbD9�r�+���U��$�=^���c�=ע�t#��� �~�D'�)�j�Zk��'�a;�>���.iA�_�M�Dw����<�Ư�(!R�/֗��)^�4�O�֔�p�i.k�>T}��ڍN��ڴ`~�m��1r4fmU��7��i���+,��X�>�/�Q��+�T5�
�� ��V��D�&�HF;��D��bHs�jA������l˖��]xeL�����jU����0��r���g����i'Rӱ_��;�~�͆�� +)q���x��ו�W��]�6$�`4!t�3��n1ixA��6~���"�	�
ܥ����2i	�e�=���
,�� T��Xŕ��c��Lc�������bs��V �O���������D�� /� ����I%-��^ ��lq��f%c�n�u�\�����o���Pѩ��Dacč�qW#�1�p/�;�<bĒ�ǒ;^�k�&�UMbĪ�:a����&hCm��r���ō�9M�!����@�<�j�9���"�h�9�ܢ�)�6'!�3��y<�l��4��d�O�͛~� 
����`ur�eB�ʀ���p�(!E���<��c����p�@���+�a(�3޽9Z�`S�M͓��h�F�Y{�A`��R���h����#��w?�@r�'+�����<;�,�n�ؼ�1C]{���� K���8���oE'���I!z5I�v��J�e��\�4c��k��������z�,/�I��d�3y��� #2���ަ�;M�xq[&f���ir,B��Si4O/�c�$�gw�,������P1F)+�=�Z����ˇ�X�
�(&�Fʈ�$I�I�bAKM���俨~ �x�LU4�V`��N�8O��s١���S���qj/�uI1L�[�`b�ܿ����}I�B��e��.I�hJ�$�P��B1��R��e����o�F�	*�ڕ�|� [O"�|�G���7�"��uk3|*�qR��D�<OC²1%~���<��t�I:,d����K־{��X�	��>C� VK�0�6���
G�������^9�爄f4O>�%S9���LM�����&LZ0�n�=.�����/Gë, 4��G6|���d=# T�*���(����"p����2��Y��-����M��� eM����=��º�k�\U��r�%���m��W��h2S�����V�`%�9�B�w��N�F�
�4��<Ջx%d�f7���k�+v8�S�C&��#VC��ȀD�[��kv�1���� �Lܺ�ہo�hz/��ek�%�*�2C��O|�Z�c=�	�΃�eɴ6_k�$��3E���ڹϛ1t'�"�ڸ��Rd�~��OM�Wfd��?qdX��w��l�h�爧�s�s�>��W="���AWs������x��R=�.�8U.�5��O�NMA3_�9�,�b1w�} �f;��M���1g���*J�]|�H�醛�8g�xP��u8��5�aK���w��5�P�2�*��^���W������Qh����N����Yّ`�cW�ML)��-�w���fQ�hX�et�u�e#�x��0�q�k��=RK9�/#x�a�G������^׹ȓ�����^`?:f[5�[�A����m��yQr<�:�B{1�
�$@��V�(�ک2YkRh#��8*�a��
�.�; �-�iq2!�^m4DWFI������D��izW�$,[��E�Ӌ��h%ooi����:sM�%��u�)!ECb����,�#�z��D�J��>��B��G#��Z�0���w<I��>7�=�sϥ]��Cn�����'�r��c��ݞ�H� ��86�:|�ȷ!�k^�'	R1�>P��"��'�=� ��8��"�	G�c:��7��z�i���n�~��}0��hf�
S�����G�S��.Z`!?J����E�y�˵�~@���,Y����!���JS}�l�����\Q�"G�n?p?��X#uT3�F�ҥ�4�u��~������c�s��94Ʊ,m���j��ۃ�_5�u�`��Z[�o< �Oc�
'��F�fP����:q�?���E �Mv݉��W���y���>U�<����
��5���ֶ�vԺ*HGh`l/����e����G���otvM-+��}I�ϖ̨s����+��_�嬶�@A3>�Mi7?z0�W�Y6HP��0=�N�+BTR_�y��eR���;��`Of#ߖ�z)I��5o����T�'W(�����K'MU|Gw�� ��;�Ќz����u`���_��r���L��?�G�a�z{�W^ʶ!li������>��t�!`6�;�5I �^�����ʽez����R|3�j�(��(ETPisF�O�"Y�:���K����o�����^���$���遀�	�7uY�}�E6��X�m��7�@��Qn���A�A_o����v��h���=���ΐ�r�⮞����@A�4�b�����l��
�X�Y�Ϧ62e���I,R�w;P���
�c56�?�(�*��}҆O����{o�{nw9+Y*}���
,�R�y���Fj�{)�,t~賓��O���=�a*�܋,�o=4�F��nhG��B�T䞬����� I4y��
�F̿M��Uԩ��8 �>]JY%p�����s�o\IR��5���*J�kR�L�s��,�l>T�u���Sڻ6R�f}��w7�A�.�8���4z{�8�U�58�p�I���b�dY��0�k�yd��a]����N��'��.S"�VW߱X��}KR<s��<�(�>��H3��:dA�Â6$��S���v,�a��R3S؇��$�>�T@,�e*�����fc`�[�Z��OCkgu�e[n�4aj|&�dxض��au��yb��I��$"����H���/(,�;��5�(|k��Za��z��+t̨��^o�x�J3��;�a�g�í�P��=w�<�i
g�&���v��?P�瘬J�2/<N��(*�P�qO��P�=Q��fpÄ�F-AN�������4�YZ��P"f���>���MvS����kgq��Z`����"�|:�"}	5C|!rE���2f�N��ZQ��⢆�>�bʼ���唻P��a�ϭC���� �p��W����=���yyW�*���{2��a��ma� 5�V�"�8I�ub�(QEt�����Ǻ%Ɯ�nM]���C�`�DS�oF;:�d�O��NE�Y�@˴�����mðx��KJ\�M� �ލ/sx�L�^�%}*ӂ�j��� ��Z�s�������X+uZ��v$�Ѓ+�e�Η��B���o�z�P��?�JJL��E�1���l8K��J?��k�Y�q���e��diߏG�yM�TG�
�3��LU��ϭ���E���w1��sݳ@��t�b�{n�X����L)/3�Ԍ��I�%�~:?&W�	u�i-"�j��6�w{,M=�(��C�eWc�.�����E�ɷ�E��а�ʀ�$��2#��!$�e�Y��ǯ���F����֔���Ac�a�[�Ă/�@����s����rزH��|�؋�0��@H����Nt��5���4�d>'��L]��.`z�@�_�`K[�d��Ќ�	L�sl��k5���>�q��<=R4O,��%纷�<�Zd��<�M~ɲ�֯
�-���tC!���i�����phYҜ\�;z�e<}�Z�Q�N� _"#�������S��Y]}�AF;���/vD'n�*�0lZ���//�=%�C4��d�n��(��W#������lD;Ur�ƍy9H�3�Vq�Ġ�/�#J�ɚ(_r�#o��P�H�:@�2T�U�)f o��7 �y�!�s7����U����J��Z�m����p(��)m��a��e*74�7��,���'K!_��?>�[k�,�`EI���,������ݙ��c��߃�~�,���C��v����o⬽������y��
uj[4��7d4t�1�����W�,CĠ��T� ��!F�L�Sv�4O��ѸRt8cc�S΄����|��z�М�Lٻ@�+]����D�j=�YB��=*'�g<ue����vɳ^�,@9�QH�'���1��&�}�C�h�`�~y�������G�)L�(e(���q�m���Ş�&�O$���B��$��c�b`=�e��K�h+��v������b#~�^�i��T�z0���#L��O"S��N�x�7�m�|B�ZR��,�W�	�T�W��و�L���:���`�;�!أ��TUL���E|z/�E����k��M����}�KT�ՏvZ�'�+1%��ЅF!��"����d�/'�6�X
�����й2���pG;�g��QX²iG��RF�ܲ �ee)�m�]�B�͊��N\�(i�܃*�!�:~cp����M1�*]0b:NQ����B��BU�v`��RF�a'�bTLg9K��#{u���A�zP��)['Q�4%;���]t���*���r�z*O:����ΎC���х�R� �ԕ͞@��\�D�M��iX�tdE�ë��S��z�a�o�Ĭ�t%d��3��u/�hv2^�>u��Wm�t|*nC/ho�b�6�<��S}v5�����i�r<J3�-���E]�Z�h��e"ӌBY7E8�Ϝ���m�VU��	e�g�g�<B <bhvş�� Η���bZ}G'��7�~ש�*�T���p�?��
/�p+������~O7#à�{0�}��r�2�Ɯ84���!��p�8�"��Fq����NW�a����9�j�	q�į���t4�(�ԀID������@��`Y�r�p%�$��P��,�����A8*�k�5�S���k:�~�xR���U;�>�惊>��BZ�M:~lY$����c��_Z����-�K�:Y�਑"z?qTd��/�=�MB��DJ�����	_%�{����ГHii6��_��bY���(O�-��8�;LHh�cΫ��}yh�'�bN�_-�6�j.��:���뀨�%�M��\�,
g�5_�ǅ���	z��[�P���<�#t�	D+��>tٚi����8w�F]KBf[�r`!�V=�R��U��k�R�7?����[g��W���Sf��'�Mj��焮㴞b+,�sl �."�O;};�˪��[�]It'+^�j�#�J&��O-�#x6���c�� ��d��k1w�S�Ȥ?�܇."�3�K�������}^Π"�D�r�G�L.�هr�G�m'��C�N�Q��c���-L��G��ђHd�x�����U|��5;��_U�>�0'�5S�*w�4�����Neݰ.�__���t`��d���I0,��F���O���ڥG"�5����
����$��~P;~Li?��YÝ`�c,Ѫ)�|Q|�Ч�Bf.L�������D��Vb�J;�.�x�X�f�6m@k&+�u��cw �}��Z���4�z��X��0�l�.��'�[<�P����1�$؈�����+֯���`��uАK!^�P�r�Q�L��V*%�B�A&�!|�0�����kM�D|i�-��ߪy��,�Уb�z-��pj�]p� �$�\G����.b����Q��sp�]?�����r�ٌ~L�ߧA]\��y`�F�&;�d��X;Z�b�����!B#ʥ�:�w5�>�$Г[�U�u�4�h���&S��{��[�vm�N;�}'�T�t�-Ƽ_)�?�$ ��1�t���\J�dC��߂�T�i<�ґ���W+ݺ�	
þ�Nw[���q������} /��U/� ������d�$�;(K��,��	�Mv�ϔ�eӶ6�lW4�w���@��\��S��6X~��~�VGȵAM��1C1�o�����i�/䀔�}�Zn��kC�p��o��l���Nz�_�VQ�tw@���!�3XP��C�kHpK��K��oЇdF���\���IɎ�Y��\X�;�h��4#maÿ�Ϫ�<��)~���XsX�%ɟ��c��#�����A<��tX���q�l�� �qw��N�k5.I�M
O����<;�kwIi��ֿ�*RK�q=�Ӎ�qtc�!l��kv���G�"Q�1���H�HDpt�VX;l��/��1���w�k+��q@�P��8�� �����rd��G�Ϳ�'�J}�a�Jx��j���hN?ZK�y,9AlD���5,ʴ��K���*0^U�W��_顖��dX�������U���t�=�8;M�M0��t�{85{�:H>��f�4n��A{����~����޶�o���`�K�d�9??�?JpG?�H�>�5C�9m�؆p
/�?cJL9�Z{�����O����� Z�t����LR7M��i$"e�}'�n�����,��G�"h�)���G�0��%�����lX:v~�����e�5 ��S˕�I�@�iQ���r�8���ݭ(�{3z-�n���S�Gj�_P��R{�C@�0L�Υ�!0�w µw�b���:�Y20\�����[�{��w�洿�����Q��{Ve_��/5���s��~�|�R�Hp��B�\�U�6q7b?����|�;_;P����<o�]���
�}�;�������b.�h�Bap*�c����*�Z/���M�aM��!3ˊ0_១M���<ScG�����sBe 2PlS���w.�.Q{��z�����@t�+�J���(��eئ��h��8�$,OO�0|�v��O�p8�֧6����:�="z������]NWV���d��t{°��*�j��Չ�;���$���(.څZO���Vp���D��g�K��fN�J���M�϶[�<s�Y�~n��B�i=�!='�����������s����Gk=���=�3�5�Z�����y��}��Ǳ�Ԍ�!��;�{QuH�Wq��;U��#w�˗�Vc�P�DS��2D�Z��#�e!� 7�P����)7���Aț��Vb����[����M���7�pd��H���Ԩ!�`���L<�?P�J{ ��=��
h��ɒR��b4u+��9��շ��l��,��dg�9�GGc��F���]"X��=�g�)�y����d�c������p��m��4XV��k ~�#�]6@A����|ᘧ� �hݤ��t+�A!,��--U>��p���dMj�#b�}L̎ʌ�Li���p�U9%p�;���#�s$~���z�[��v"��޼5)�Um��A�s+T��x�G����	K�yo?�s�dя	����,�bW���3�h%��V!�o�sˍ�O�on�zX�"U���y�x��ܩ���ZZ���>��\�Xz肃�|�K���"�{vV0��L���$5�<��u��hL`v։5X��V�y�%�T=fBw�+m-.gٕ/�_y�ɶI���n�����̜����A�m��s�b�eC��fI�GrT��V����;YwOl7Ҋ6i���t�7+��f��-��������h��>oj9��enLh7�䔉���]�B^-�0���[$(��Vs3a�X��D����'-�ə��Z����!;����⒕$�����%�M���Jz]��m��A��a`c��C������c�-Ē� L��q��گ��Z�� 
��7y���h�ؒf�:t���j����h�٣(i���
�0�r2�qѼy}�ߝUz��9��k`Ŵa��5jٚOu�O�-�4��"=ة�ʯw�'��]uH���"�͓� ��H�?[�+J��PR�>��<��� ��q*c�)w0����������b���*�۳������|����hg��@��,[���r��H� ��}	٤%�&rNqI�?zB�8c���WBH*N�+��	�D̽b���౷�	�㇊�FG���j_��>�4x���4�c*WqO&譈����k�d�����g?2 �(�&f Ui��LYD�*�W��:z�F�Cy�"cu��	��i��3�����0�E©=>�	1Iվ$j��6���"̼m$�e_H�n�������ʊ��-�}�8�gd"Z�-N�WuU�Ml�6����B���}ݢ�I>]��ZMQ�jF���B�V��x�NBV�`O>P_`�nY�G�Ѯ��C�L�Md8G+��&��m4��,�ȿbER#h�8�2m�w�ۙ��� Q>�췅����Pn���uCS����[m�n<m�x �z��r;��4&zZ]�e��)�gQt�x��`6]�$X��|������m-���<*q���z���J��c�#��#���};l��������0!A��ϳ~!McJ0�6#MM<�;ѥ�EA5O�LF^�>�Wz�pts@�S�A���z�EY��Cx�a��fuF`ol���~��;"Q*,�`�<�3nTI]��b[z-	t�V�$������8�^1z��7W�d-�Ǧ�_���}�>�"�:/��8Ē�d=DP�b�\����?����U������D���,�z�=�X�ޭ�mr���h>����.�V�C/e����<����E�Q����E>��u��%1ӕ��7�+Prp
�P�}=�������7p^��G�gΚ��y1hO��U}�!v�u��ʇ'����?�`� }�t���W��d�Ͼ4jIC�Y��+
ߜ]�W݊7���0������jѓ=�A1�(W~����[R~|`����'�#���[K-oZcrA�P{/(a|�V#��]	�@��3Ň^�+u�&�ȋ�����WyK?x��`���6}gD��V��>��PW����	�F"��+(|`��j�YH�^����ܸ�9~:�r�m����AsES~+�%	�Ps�#E]��t(r��Q��#�Ⱦ�u'��ك�L
�n�����me�i�E����=���
��v�
Jৌ�*^�u@��:�;��p�u�/�s,Y-+i3��D^�_ɽ��a�eު�+�,��&t��l1��<1>P��j�n�ǂ���&i�W��aZ߶Ra��ŉ)6c�^ё/R����]�Qʙ0y�pz0����L�6������|�r�UI(e��*��͉zV���8�24>�u�.����!�- Js{��]�8L�'�J��<C�2}g����	O�K�U�1��]T7����hm�K�C�A�	����Si  ���9"5�2��YL��;���`�)N�����������,J�`?:��1�y��!���h�u2!H�.Ÿ��jŽ���C�&�"�����C��Y72�K�"�%��l/�׮�.n�\D��f�� �h�3g;���������-)ۨN��9�[�kFm���?㝿!��k=�e�L���+mZxH=�����0[�خY���
h�_i���桪��Ϡ�K\үc�} �QXDr�p+���L�35lO�A�������T_1~�"��x$�5��K����.���<R�F����?�I���[���Ec~��G�~m���C<Ǥ�f%�,K�z/`���ڈ�`GX����$����F 8����Q2��)��.z��hL��]��B�����G��I?��:���r�4ެs�s?{����%����01ձxkV]�9�6EG��xp�V����]|��[�2b�H�,Pl+���F�ٷ�fg��.�b�����_���Λz�u�w^o��5�����"�1����Y>�Z�Mc�V�ݖC8�(a���JȈ�$Z�ڻ�??�T$?�6�x����= ��>�g>��#���>�ڱY�W]���1�/��|�Ŏ�A7��fq�m�;{<�r�S0u�4 �����\Vڂ�CTW�L!��캿����1��yl�~r�.����
"�>�����-��0���Ν:�y��`Y#�	L���j���;~q�(��ֳ�%ۀʻ��:�b����6ӼΪ�ir%)��u$E�|o�s��nI�\�H����҉���vNQ4�̎�]�bٗ+����vުD���x�Wqwԏ�O�Y+���/=CR�Y�\j�v��D����!f�0�\�]z�،Z+�M������w9��c�y������c]�9���x*�h����γ�Uw�R&��O��!g�8���Ҁ�a�> ��=Hm:g�.�c)˿MŇ��t3T�>	N��_�uu�� ��T�m��o�?���k
�qx�`$ll�Y�E;�{3�Cz]����R}�Z�$�r��1	�:(e�@�X����w%'m]uAp�f] �>�|�'�{ڃ�A�I����<Z�(+7h��Yd`M��gctm�?Y։oi�۪����(2w�^�'�N3�;�7Dϓ���!�A�s�����?i�J'��pC�1A�X�^_�C:���񁿕�xP�ʳ1�Fݛ5�Lx�;b�|?��;�J$(ډ�<��Z���WF�8�,���#S3pPT� X�t@��1^�&d���4���'�
 �c�>g5��8�~�O�������k�Oy���l��{8�}B�rZ�K��P�ť�́��rY��􏸯KpD]���O�q��u��U�L�yh�����ʮ(`_��$«b�	$�+�>8܄�I� ��{(oM{WpÌعV�ù�_^�6��]��_�A���LyK��� U���6)5$���s)Z s]�o$�Jz��""��0D%a����zD�G�V�z4w��s�W\��������&?�
����(�*-"x[Q���m��(7 hv>m����WԴ�D�Nԗ�
`��,�3(죛��������g�
�>�^��E'�k�pmU�/:۹�f�nmzD���bp��m�s���n�̼S%��ƀ������A9���l�����@��������V/�0�n�g�⚯�� �^����#�4?��'�V�z�5�����O��b����5����i���=��"\�=�ރ�����7o��, W�98 	���щ?���'dQ`kx,l�c��\E��ʮHn�G���-��=-�C�� J+��	]�����]�sʿ��i�b����q�nJ���Y噒}�Ze��G�;��C˰s�����ӵ5�W㶢�^�	���ql�;��8�'��/w��K�a˛���ƔB;��Ɗ��8?X�=x�-�Y�R�f����>iO4��n�p���]'5*g$u�5I}?���k�gkų�ؘ'녊�ͬ�$�-
·�F�d�7d�B���@)�4�an(I!*��	y�yM�^�h6�Z�9d�Ⱦ�]�x\b�)�gݦt*M+ڕ s�b��eO.��E<r?���rO�W�I��d	^ļWEH�p���7���a RZGkBnEԧ�,�#I��o�Q+������҅��Bm�v��>� ��C��`�@�p�~���`8���y�v��k�����u�&�f��}���j�M�	�Nd�W����r~�y��{F4�wD�0�}�P++�����!Я����[��.����<���A��֭��u��'G�q�O$R�n!I�Q'R^WJ� ֨d|�s�5W=��=�c|<4�۠-���<j�|1޿��b��%�L��,"�̅G�{�c��a��C��:J�GK��6��S]��*�K)���8%�}/_fy?I��;�a3�¿����%�S�� @��*H�<q�J.�"��Ā@�x��V^F�������MpBJ0���T�=ނ��_M.+qf��V���'N�s�֪�pMuhc��ڌ�s��Qϟ9�׬����ŹZǌsE�-��?�E�0z�:*�!�jI��}`��Un��<x����v�B��cڧ58���c=9��e~$��(i��3����'S�55���b�o��4}Ȩ�b��%7d��O����h�s �6@�5P���2��"I�Ԁ�����l�I8���A�&�/.H���9�W�y��+?�y^�Г���O����R��B�x���b%�k�V��5a��"8.���J�P��x޾960#�EpG:�D�x���lZ�{kf|��o� �s�3GF�%���f�b��7�&�DY��c���sm����,�ǁg��!\,�
_��R*��N���i�J�
^*���^ܽ\3/�bE���tW2	uQNK���z�T)|iBQ��GF��JZnEJ�W�v��=N �U�L�P���e�(����y��>�d=��cW��t�{{��?�l��^nC�<%NT���P�M��V;�*`�0��84ei�{������R3ؚ�3�RX/M� � 3CݗӪ�aR�+E�R2Bہd�V�u>��{݋$Fe�@5�*�����v����
;8Z�9#FO*g0�ޛn�B�:����.�t�}��Z!���`��3c�B��F��w%D&�9�.��,B�r�W����tM��f�,�kn�=m�d
iG�*:5 �(W ��(�����WXt3��Դ�tĹc�v7ڴ���Q��ܶ86>�>��e�5D8I����^I��u��A{�0�,-�q��
�qǁ>4테�� U����k�G9H�Vy��(I. ���6~k�j����;L�g*��i��!5)W�M͢.#w��z�W�qV�����}�_���3cW���$��X�ڷe����Т��d&5ڙ���DA'��@d����"��|؁�������x�:P<:�L�֗)}\�rI,Ú�͞�j���������'->�Bް�AɈ��<ZV؋�"�7\O`ށ:,H��D�@6=�4 �����e�4_�떓�%Yӑ�!�B�c�I0/t�f"EJV.�ߺ6"�
"1��N~�/��KA�A�Ϭ�ŦA���O�v��/vC�s������	=��x���b�"���Ki��{Az��qA	晘O����e�D�a[������%�$Q����£s,\��f��[��X�J
5Gꭢ�����4����G'rUI�X�|&�|�9��tL��(y��
���=�>�Ó��������3z����j����s{Ɉ�I�`��v9|UR ���чT�H�ja��R��P���۝��Ql�o�����.���D�(�_��ӞE�؏��� +�-U�h��a�1�x����TY��j��W��'o%�kvm&�m���V�k�L�����}E�ѐ.����A�`�|�j}p /��ff��(L���f��xQc�����֥@;'��ۭ�3G� ���l����#��3��x��Z�KG�FiБi>�GmO��e��V�U��@ȓ�\65s�w>94<)�s����CE��<�N�/CrA���K��Ŝ5r����pd�-�;&��{:�`P=���?Y�4ɓ�W�5�ǥƴ?a�=�>�$xP@�ߟGJ0r�<ۜI(t�8�c����J�:̋���`
�f�5�.�0z^�ZqAe�\:5J��]W�QKƹ����=��pJ޿�9���ˇנk�ǝ�M�0uӍ0�T'~xZ{����P�`w���g!��J�rOyVa���ݑ��+�,4��2`}V�`�MV�;�!A'��th!$TU,ʸ�/3�U�����n�%=$�K;����pV�9捳I������E���Y�MДUڷ*�uJK��R�ޯo�<��.0qQ����2�s��i��Y˜�Ԟ��v������m��*��B欦��'U�*�(jRJj�33p�Z�J3������0�C�w��k}(���/�A�N̉�.�;(R?.�L�x�u�a=ܠ�����6�eM�i��vT�B/m���-?耳��Sc�4v�	?�l\"�!3?�n��&�۬�.Vc��7�L�J�-@�^0S�R �P؇�ć��������ސSO�,5"?�?��E.D���51&��[g�`|	�G��nd���Y�R?�5�p��'n*��ץR���:AOK�WR
���zؕ��}�H��i���f
��ې-�R}�����*p6#�����{c�bIZ�o�\]PF�t5U&�/���0�J ������T�j�(����v<5����S����2��$N��/T?��)�̔�mO,�-��Z�w��N᯼F�EZ��c����>���;����Aj!J`����y��>Ε�ꌑ��IC�X1�ٱ�%��S��S�P;(����o+h���U(FsQ�so[l��}���F=���C��[k�?k���j�!e�J���:�����>�7��Y�w�HA��>G�w �Ȟ���(*}(��#�v�"��%��m�6��v���'��a�B����ed{�#��
�Y����=�7�wD,c/�I��xp�� q�wA�b���HR/8�,�D�,�ݩ��V��7𡋎t�U��wpn�v%P�6 �s�=��k	7��V	huv�X'ǘ6f#D��](���7���8��\w8�J�
�jmH���$�\Q&�!�mJ�W����c��s�m�P�"�f��}�e�m�9[��M)7xhN�E�_�U�f�OS������_�1RM��:Ӓ�.KCͅ(^���	U��D[ȩ0^C����2���dT���q��V����b��le����� _f���{��a���Q�E�����S��KhC�]�3��0p�9
)��a١�h��:�Ɓ��8Da���+��,��Q�{�M�`q����u^�k0�Ș�
�f�G���r폂��q��6�%Y7{�Q�-p5�T<������&m���H�O��e~ͯn֖��C�F^B��dy�m���v��c~D1;���pa�O���zu������||j ��:w�q:m&�����:
[��'�/��)mˈG*�lrKJ]"	���=�R����+\$����J݇2i#��3��wCr�z�P���y�![��TPW'(ί�e�l��+o/�5�<_:Y�R��2̀{�k�7q`C��V' ��$��~���� ̌��i�q;��'�v�a�����N#	���L9wJ�j�Q���@��sb�#ᩙ��3 ���1���.Q;��3j���� <=x(����b���m,�����1�H��GO3L>9w�8D.r-c�I��b2u�����cŞ�3V��I��	A
&�2)+��3qĽkI�d�����������nYW	�oE�2�L[PV����!?8(�-ꔛ�fA<�!Uf�g�dbf�����|Mb��v�W|ȓ}���z��M��؛jB��Ioͅ��y����;\~���UHz�?6,`(e���}�o���U�j

����ƨט#�kؓP�l�=%��i��u�����h�j?�r�~�����GM�BP ��L4��LƳķ�Jp��?�_�W�z�o��D�6��*Ɖ5O���b8�s_�ܳӣBs�Qq�㳬6=�Xcwp������RBϓK򿻅�j����l��;|lڧw�\�2�����ig����_�UF�z"�zm�ަKn�O'h��%��n��c*�DG�֋T0�	 5�� c�)��=�QMx���"^œ�[�=1wY�'��+��P�q�w��e ��'9�ina,�<A�
�B�hW�QM(K��������M7�e���s�qU�I��d�-�N�ݗ���Z+�;^�x�kG��8?�Q���O)jG�t��}���%5����؇Y�#iˡ���1زИX6�S�a���Kjj��r|M��߰�<��(�fҲ�
y#���P�@hI�wd�j�}�<�2�'�ب����e�vg��?��?鐭�H`9)��c6@~1�qPuo�����a7e�)���]�U{`T���
������������<���U�G�݇碡��`h�U�UT���q��`bz���Pl��&��������+c���J��~��>��Э��k�э0'�A�A�.x�z�R-�ύ�h��t~�|5P�e#�%3sg ���I"�:z$��D]�j��b����)wkT��>�$_� �6�>�
��Z�{ /Ž'e�[�Gn����yo���8���JA�`t���f�z�a�Y �p���e�)|�`�("!�р��&:x�>ݠ��PHx����6�:���|��� �n}'�-�8���R��M��wZ�h�̣�/�{�BI���^cL���H�!�t�G�ٔ{+B�+q�{m���;n�c8�<I"!K$7�f<mο��1� �˹��{	���9�jEn�򏂝L	G}|���ꅳ�.�]%��-K�e����f�~�|�r��D�2io�Y�Ua^�na�R��b J�2����3Ы�IlG�G�(��8_7�G�����E����F��u8="0���PD����4-�>�&���bu�"��7��-[X��+�"�q����J/��ɤa�!#��̲�
��~ٻL��Fc�t�S�yz@nB��bw4���$�p*�"g���c[$YP|�8�I�^F�����a��%��r�W?N<������W��E(�sK6�R�S0Z���VGZ��'~0�n�5�@a����zF}����p�̑ �m�y8�%���i_`�R׎��w�:�C�����	�1*̄�U���n���>�����Љ]v ��)>KX,��ԤZ���B4�b7Rc&z�ީL	)�Ȣh� .��x�0|��A���=(&�~�"��$Ȏ��D�?�	�`�.Y8���Ձ/��^�rb�=l]C�+�iHבL+��/▰��\I��SϾaۯ����n�f����J��l�T�,e�J��_�&E�""nWl<�6�R!>5Q���ek�A�]��<5��Ws!�h���_J��=��k�6���Qq�#P��P.�4_�,ғ���w��~�+��N䢁� t��+ƞ��|����b�`�	M�9]��>�� T���e�~�g�L�Cd?��'�#�x�"�;�i�K~�y-��7�/s1�#-��Ԏ^J��tΓ@]^.��S�X|���n��,���'o`�?�vv?�%mٙ0d@����s���H�a���Z|�B����.�r؁����RF1��$�����΋+�)ln+�mTb�}7+ii�|@Ŭ�[-�	��!��6�~�h3^�d@�ɵ�#s�\4jjp:�u��Al=�q� W�$�ϯ�᫫f|�'��.����.�E�g��h56Q���M9{@�Z�ϩ.��^�\�3{��[8�D!�&�����f�*~ 8 TC<G�\h��XXK�� �����3163�x�BFb�=�Yw�6ޥ2���)�:3���k�$d���%���E�s�l�8�����V��,��ԑ�T�0mb���n�Al���_�ˀ<���S�IB�[���=��M
��T�;F�v���-�<�t�+$�T�!9�Z�Q�842[��<��^Ё'l.�$�O�$,�>�ݯ��oe�N�7��4��[�K	#L�hY�o���S��V�TJ�RGn�$K��f��?�.��ʖ�9���B�̅�� �!(��`0L)��nE�����&(ki 	S �\&��)<1����7I=����WȘ7�Xi�jB�%��݂n����\�QG�]�M:^�bP���=�`'/���F�tߎ��i�sL��#Vty�CEi�����;��ހyzlO#��ͅ�*q���#�(�H�8�\�T�Na	鸍|�l޻����M`��u-G��W�m��3�3�ה����_5#4�\�n[�V?����7UGIA��~,�%��]¨#�/YҞ# {I�A��R�}��D��0�q���ݟfV��G��g��x��˵ɉ��XX{�2 y(pn��=1x}'i�ND<@\u;n���e�as�O�ZNZw�:8�aI��<�qpz�)��]���K���?Mmu�ӽI,��e���J8���A��B.5� ��?OP�D��w�	3V���g�8���6)�5O ρ �Q�Z�%
����_�u��u>|z���MW�`��5��E�)5���&n�	���Y�Q���� :`��AS�s���!Ɇ�]'�~;;�oM�ot�p>#-
�v�����-���P�T�<��E	�<dX����_�6~�;@V�M̓ƍ�
�,��_�5U��a� �n�9;H�����Lp�q�ʘ�j��ǥ�1���sT	�P#�e#�V�q^���	&�R4ݓ��S�h��[��'�HMSu��AәM�R* v�OQ����14�,[�X�~xn�`{�RO��:w�}y��-�C-��䬝W:��ƽ��"�s|�uH��㦑�L������aݼ�aYH�<U����Zq��@�L�����}tn���B$��i���ډ6�
v��'(Yi��V� �)�����?�s�0��v
�:Ŋ�f� .��Fr��	�_���s�3])����7��O6��F�)G"j��yD��3iH�����܆FrH��qo=7v��|iI˲��5b�_�Zv/T�A?�k���H��(��;)۹Z;�EVQ�