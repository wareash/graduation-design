��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jåا{�\�u�?߷�dn@6�zf���F�ѭ�hU)F�4��A�Þ�
<��XK{f;�F܎�9)a�_����1����r�����ij������HVl�޳!���쭁V~R��aX�������5"�I��mK�����K ɨ�a0�}� ��RN`
0f���c�M����cf��ü�G��>���!v����Ⱦ-�D�h��[5�%BC�4=��p�T�)���̿t?���8�������ܩ��S<N�a�lߐ�'3�\K�xr���1I>��H[T`����r8'Z�.�NnS�T�|��p=><�k� ���m׽�@1ggt4����*ه�?�4$�@��M�͘
d�!/r�d��u���`zg{��Q
�Xg��brdZf�5�D.r�����Z��J�r���v��tE����(�i���k��������#��Y��d��d���.h`IT�h�}����3��?+x�u��A�)j��ٿ����2�6��m���J?�U<U�� ��T���6B�Q#V��%mj4q����#;���uc�D-��]"��`��,B2\�v��AI�*e�ċvڀ�4�����Ӏ���v����ipǈ�}4�YfB�W� ���w��=�Av��K�e�[�S9�T�@A3'�c����w��@7.��K�O{#�|��qfh�<$�h� �Ռ���;�]��C��,��\DV"�E���� �D�xe�_�!�^��OM������m�WV����6�H���j��i�!���̷�L��që?�!�+�%>���(nC4��աu�n�·��}..UA����VC�i&�V�Nm�PJ��?b�\�p�����cB��T5άne���d�R��e�E27�M473N��J�8A��������z��9>L��N;���I��rw�Q�[��6V��	f��CN�ʻ�Yg}�i�Ԏ\co�Wo-��`�g|�#F��ҙ4���r������s�;h����mt���KW��}|��1]�3�+�gM�	������H>1 m���t����Liɒr|6�s�#��@%#a�hD���CGe3���L�.�Xu�Ҋ�	����ácg��Zc�f�W�z�3���"��������x��wE�ʺ��H�KGd����.�ԓ?D�M�3��C4i�A��g]�Iv��V�)x��߭:�^�y�n��o^��!.�=۵kJ>����jtF�p���M���|����E�#9���3n���hN(jL�ss�9�v��r)���|�[��b�;ԁ�`d4�&-��^vS��͎��o�]7Y�Jw�Z�?x��<fW�ᒟ�5��ut�Hj�D�`Lq�ƚ�z�9�u`:7��Y��t�j3���*�f�lm���N��n'���W�5�!ZƷ�L{��i� ���/���e�UL§�����	c	���x�_�I���9�(�X�z���z�$�%����
w�W��׃d����Y��TZ�i���
���%�MK��Dl^A	ֱ�Б�?N�=�-���xn��d>�]�#�?=�q�b�d{�C+�k��?���4Y���8��#�Ό�M���,�4(ҏ V�,�Ts4���gE"k�e���*�1Q[x@���K� y��64�B`���nL�?y�����J�޻i�{v������0_n2��A�{1��Lc��V����Gr�=��,w�u^�x�O0�;]���oE�����O�ݤ���\]@j�_���4u���Ҧ� 1�n ���Ӭ09|o<ۖ�u�&"w�$(��R6OLm�|�,=�>I�����O2�M1�����Al!�	��4\�m��Wl<���룢�f��cE���ܥÆ�k��H�Ԩ8R2x&��#:���\i���-��Ǐ�m)�s�r��UI+�Vr��י�����*\�=�] A������~�!������t\�����Fܻ;18���hk)YiJCMz$c��}�\�iЁH;�X��.�h0�Ņ�:p��1FH^�� j?bٓ�������=��1'�`��� �����sF�'�s������NKl��^U�=�	�\m�/��q�qN���r?���u�!*�d���o̽��+�X��W��M�E��L_��i_}qfK����G�!k���8�*ގ'Z,6�E&k�v���G�=OU�:\�ˍ�z���]P������3�
���'@��ʋ�4w�Έ����J��+o�latES��mǞ�xO����-�S3���C��{P�6,ҭ��6�F�C���h��( ��2σBJq[��ix�"]7��7�Qvj_+~�}�JPU�ba�<�)��@%P�I|���[��`Ο�
������эDe�EE�`��gV�	);�O�m�z���:�p����3���٣�4OЎH� ��Ο����J8�>�CNS~E#��8TX����V��#���V��Wmw�y:���E�Fs�cX�1!-�5��){��B�'�A�R�Z)����"�w|%��)[��hU����3�Ȑ�������'gN���@}YO[����|l�	8��$�r��ѧ�c�M1�M�$G�^��ANo3lƘ&]�L��ڋ���$�	ˆ(w��Բ�Ѷ�uY�=m���(��"d�e~�	CD�;�B�-qY*8�:���5ё���M��B��x��CvaH�<ky�~W�m��{q�B�נB$dН��S��\Gر�\��P�5��2��f`*�_�6iw���>�Z��*�43[��h�D;K�i=z6!6�HǼN���n0]��T%f���U�08i�LV,�2�UGL33Uo0i&R���S����ADy&�Ұ�=������^RFS]�a���6�7�V5OјV� ��{��/8�z0�4�������=	�S6Os������/ ���t���n'� a�� ٩�Xl�RDj�'iH�K���/����̨�<�x��mW�d��K��A�arr���p�s
�.��.��4��Eݼ�MJꪧ��%��P�/7���&�
t�2�d����E<7G�Dbu�o�sB/���t�Z �z���*��:AO�����O���d�|ڇέ�vz�������}�$Ӡ6��@b�S�y��X�K�e`�W3[&���h	 $��5�xLÓ��>����饉О��x��n�����Bʡ��4��k/���\BGl� ��1�� 0Vl��
�$m���0ƶ�B��mx�����ၝ�8'���/��%��K^h�\��a{5<Y�i*qy�;G��(D��~�	�f��r��f� ��o�Rh��H^��_0M� �;bSg]A�_�bΉ�6�-��g�a6�z&�ѳǎ8u΋k3>�~C'W�6�g���J�E��l!��Å���ܪ�R�&7�<f����}}�Qi�zM|jZ�$c��%����.�X�ϙaC��R&7i^S���3>�9����X>b�*`h�l���p�k.ʀ���| /؇�A��0^Ng~���V5��c���v]�����A�����V�:�YS:>�Kq�����y�s��U/1��bIZ��'�!���Qs'�����M�7k=�����|/%+.�<�����_z����d��o��� I�x�?��`�=��QC .A<O��R9�[����7���qF���ZN n�|�E̓g��k����KC�{��g��ҝ�6�Pf3���:�}��g��J���M�V��F��f��LF�1o��>-�8ݹd���
. N�{�����V��s�A����qZj��� N�-&r��Y�Լ����CT��
{CT�X��wC5�6�7�����>0��癿6����z̴��H�o��r'�qK�ķ�GQf�)�b��+��6��$a��;��Ⱦ�'�F�}j�s��^7'��"+�.��\�=i��q�Yh]7q��$U�A��aMv�.>�U�5���9�EM�
L�������b3OA�������Ë̪P��@^���zrM���}{V�����	�4!�?�乕]HV��� T^�G<Pf+"A��J�?i9&¸�.@w�����l�Y(q�D�E�� �z�3Ly�����B�D���sPk�5S=A��L�>��oX�K�R?�u�)F����C�\�9�0�O��}2fS��|��9�ҡ�hc��-`�@���c<�	��0N���9���BJ�-�g+B8��Q��U����S�~5zem$8m reOS.��e�kv��ʴ4_����a��AUx�T���j[	���/O�X�`��z	 x��ֱ�J߅3u%�<#U��
y�z�#g`�^מ{D�]�b�<�c:���nlD�n�$�o����d�B�
���Q��+�<t�oD/'��izo�}@� �� 9�#%T�#��Aٶs������&�l���ov)ƾ3?��d�0_O�#'�nT89�jWS@t���[�'���]$j�O_�ez֦t�Jc�zD�=���k��Y���'B�ʖ��Qlim4�nCf���Z���Q
4�9|2��U�&�\SNQ)&{�nZ)pn&�si�݉�Y��b�7�&�z�ȴ����y��B��u,�*�쭷QC�q���W>���I��M��|����U�g�����'�]B0��(L�2`σ2���OZ�����|�Ba��Ɵj+�W�O ���ǩ�^���siI�����3@�~j�*"�1�Orjl�y8+v����]	 ϨC�
Qt��LA!>�zH0�� ���T����YZ�����e #.�a��4,z����RE����K��ձ�[w���ʸ�lBg�xI/��q�m��[������I�Ww��8�=�.��J����:KT�@�AO�B8OQ��q�,���Ke�Dׁ��S�
�1�WJ3ЯJ��U�cf�3jc����F��[��!^_�.�*��R�x�D�g��b��ĹȻ�H���)���HX���B�=�h�(8ږ�d��`dR�F�IQ���16�������pƲ��kcP9 �<J�8��9N��:�<@�>6"\�S�����{�bǐ:��	{���C���j��bAJ��&.��A��U#,��TT5O����;B���x6Wb0��3K���,��(b�v��.��n�Bjs5���e����,Ԝ����S�}Ƶ|�p����|�W��UG��Wl��+���3<n��kh���ڕ��+�6Yr>QR�B�M�srs�A�n��S�Yf���Ȣ����vc��#�\�+�Ť�#�&P&�͜>3�8e�R�M���a��ˠ^w��>�]='D�������%�S�L���>����a�_��"����6���^�;[���7r�^9?��z�@���+`:%r��0u��̚b��i}���M�� �u�K��șqJ�A�Y ^%��~�5W3�K�q8��*yЍ����y��J�_���&gg�:�.wN����A-Z���V�~)�F7��1���0$٧�(E��K{o\!*��#�)nN�V�,�����'�]�ސإ�4$͏2�se�̃�2��U�ͺ��6���=@I�������*8�y
����ł�,���-ĸ|�Mď�6��^db4�����`�}��SUW�v9�s�]�c<�,Ģ��2�]�n�q ���)24��S��2f����v�b�W���_����,���Q��A�Y�8ޯ��n��6��ke
�}�^���L��q��j�n�Bt�:_[z�C̻�Q�Q�[������Бk��I�z^NQAx�[ԇ�̍��k�JS,>�6�ہU��h��;��8���U��(&Aa�\1s� ���\��Գ	�?�ip���7O�v��1��FW��z�Vyp��
�lt)u�Í��W��'��O�,���i %꼙�^6z҈̲
z�++Io��.mY�`^@��-?D��մ��e�N7{���-�>��@��O{���wkT7A��h�r�OL��"J�S�u^��B����%��1� �����d�+m2�$d���ƒ@��DJ �X�w����`��&�,d�y�^ODM.�\���]k�ԩ�������b'SG �v�Z��+�}b�cL�6�>��"�O:�� �V\"��꣇J�[�^tZ�W����WV̔��?[?\�|�<Ѹ>I	%���w)�K���X3b���W�D�8R��}୬���O�������(��#�!:�?����N����1�p�_0��<P��tp���t�}Qivu�[F��W�UtLF��JwfwUz$�WH�c�mb���	5QD`]���\u�%�i�D`�����Gn�NDĚ�Y�~ݹ�;S�UX�6�7����x�=�4Bh��P��4��|#�1W���iل��P�o����پ����$�Ƈ��D�ገ���S�X�g+5M�����e��IF�}l�.��?M<wj�`˛J|�W�J3r�ܠ)L�}n��� �D��2 �|�F��}$��*rb��y+.�H��o�+��[�n
�b��r�j���ԙ���!�n�ګ�Nk��Xf<gf[�߰���OI��sVB7D�ۓ���obw>Q\�PC�^.ş{���a~&ny�V��|Tm���=G��[��x�̀0������m1jFɴ��r�!�h�
eL�,*d`���^�1��a�[0,�
�s�Q��z��^��o\M�4��h�H�i�tN����r�ϧ[����\!Qj���ڵw/m��,\�@��&An�cޠ�]#5wJ�jlyt?+���!��em�8Ǜ�IM��
J�I�J~��p�.�Xߐ�a��������l�K�{������ (<�r?<�[����O��B-��#�.=ϳ�·��s5�Hwn,*�~O���[��0-�ٝ�GRB�Ǯ�e�^��16���}8K�3�H"���g�H��b壨x)�8R裹=���D���2��sJe�k�7r(j4���$�!Pa'rr���6IEI룬V|���8+8cvK�K����K��9�d�PG��K��yv��H5�8��OG�Њ�:�q��RZ���O2�r�$��x�7�c�(T���קZ��T#Xm�a�yKkU���DH��}:הAK
�r�b1}
.F�Ip�K�������o��RiHz�H���82ҿ��Py7�>*I�F���m��7V�鶬����g����kͻ��7�4�E�����B�N�b����Aǡ�Mv�\f;�����c"�)vxNاla������ ����+٫�t��������c��况c&Q�f'<�ˋސ3lDכ�1=eY~ص4c��4���
>��Fn|�*� b�-[�1�O����C��I9�C�1JF��-g{�!35����RBL���O�D0{�t	:1p9�e�)ܑ,7��Ggd����V���[�cP�<�G��F&z(� ~�ˤ`�y���b���D�82Xl�L����amDyK����O��\Z��<�p�+���Pu)�6֔�ltI��+�A�{j�Q�D��8���b�w��#�!��?�-�I�; ��ʴ��b�(��3}�ܵc��%��V�6_���fw.�۽3�+�/R������^��(4���,�I�9rQ"~lI�n�U����"f-Ĩ�A�*�`���Keo*z+(�7��*�����j�vgCL�α�蕦ڕ ��<_��ف/}*C�Q��I�84��^ȂǶq��ͳ����-��<ɏu�OPs[��^�qH:����C��ng�!�5�<�?��P¬c*���Ƌ`lOdқ����9O@_`&����X9���* �p�0>��Nբ.������ �ޮ�^�3�N���Xay����4 O�D~�pzr@����fB`�8Ѕ\���f�-jr�C���U�n���hh�A�i�jy:���_� s0��&\�r?��|�!�� ���w-s�P>OK���EÍ7_!ƏM��U��b*��A G�����ɽ)�G��(��D��<8̖4�^�Y�X܊'�<��G3�*�V$�)��}H蘳��ި�j@�I:b�	[kIoG�0���rM�-�1@'�=�qb����d�(r~E5D?��ь��|@���ݦ�����d$%B�	tg/��w��UR�'��v��S�6�DtW&��B��ѳh�����0�椩�"}�!�6��3������x`A�X��K!��r�6��u$�M���K�pBR�Sa��٪h�O69v0z�y𦠷8��P���"�X�W�o�(�F��I��Q�+�p��ܑSb��B�����~�*��̝!�s���)2Q%n�LQ@+��%�)|�>��5Z�/�~;���"�5:�h�
�*�G[�7rj�c8fE�?�,������K!8�{�\S�M������ɽB#t]fv�n˿���*?xi�ü��rq�b��Պ�T�W��"Pr�������Q�7�A�̀EP�ދ���B���GSu�Z�*i��E4��w�NI�).� OR�����M���%��5�m�������`|�$rѼ��*�j=5->�W���t���&+0�����;�[�Are�O�*���^u��';3�/C�/q��N-�ݺ��똾z;Ўo�h�ɓ����n^۳��[y��<��F�hya#�D-���*DH��m�a�Q1��)��D����:��~z4fԐ|�,C�i:��D���	�AW떃��z�O�n~��Z��m��V���s�e�(]�<�7�O����/�I�`���w�B-ߤp:��w{P��;0�r�5�+ u�H]�>�JI��P5i���>-NA��{Pm�}K!�����D*kV�o,���M����c�8��9* �H|�5;I o�k�������������`�7��X�Hoh��� �L.�4l��_�\@�d
��BFGki�����C��?��!�±�q�^Zs���)�����ޱ��y[4X ����)�ȍK��ɣ!��$��`ʉ=�|�#�e7H.j��;;���0��|Ɗ�r�P�-mun���n�00v��[	��Q��t�5H�9�P�7��م�*��3cY�<��)�+9G�2�ơ���'�Z�{Ɵ��q}6�Ly7I�詎 ����g9���3>���t�D�}ZY��;A\�9=-������HgF��r�0Z5Y�]����=�j��cO=p9���G���(�P_U���v��hP�9��P�zf�9� ~�s�Nq�F�3�T�Ӯ��Ij��{���]�g����a���2^Y��w�A�N�!�$C�:�"n�`_����`���{ā����Ǌ�J]v��Nv֬"H�������~�Z
<3R��O�B2���J����8&吝�|_[|�����9���XC�Gz�l{Q��Pb}�܄�d~�$��� i���S ����De�
E��N��f�2!1��C��=��Lt�܋!)~+,�����[�{&����2JQ��[(!���BJP����ӵW0��p�f����7vBC�zp��sN��R�7F�N�������m��wJ5}�`B�������%���n�}�*(u�J��y=&�O\��u�*`>s�c��oF�&����Oc��%"TE�{ �T����3�!�����	�0<���VL���X�N'%EE���v�Cjk��?#��{��b��PaiVI�}�ᨰ��z{١���=��sq�y��_��C�(������ $S�F�b�܂�M�Z�1xVܓ^L�[{ ;$iW*�Vj�s��r�~(~���Z���0;�A�3����h%L4��$�;�z��bu�O�
�{}��_�kޠ���������{���Tc�!�y��$m�k._i������ov�N�g���`3:*�g�[���p�R��K�E
v�J���J�q�}��@�X��S�`��F��o:L�ŧ��y���&s~Q�J���lX�X�*(?������*B<�+���ːc9�e���'����B'�2��_KU[�0�jLM[�z��oڃ]�C��`d��Q50t�}�Fl��DJ�-�����t���,V�ILq���Nn�<�\�#/d�&�9ó3<l�^���C/LT��)!Jhr�f��7�Uɇ�9�8"��f\����Qp�=2��!ӭm������Ǉ�!�Uc���0�{�7$�T�R[�Tܩ;LGe���45��s,m�&NgC����������to5y��z�z����/(��2Wl�4W@B3�Z��x����"Hw����_���a�����=��!*&v�h/�x�`�j�D�:���Y��o(0�8�X1�Ե��;��<��0��=+�6Y�<�c���	�Gj[qk�����Y2z9Ť�8��8�t�sF���]y�3����eН:���8�zr���,�A��,��ޯ�|-\��!ZXE��Q{���օւ���#}O��.�܂��%�eٖ�"y�$�P?Ot�(��m:ӯ�C��۹��)�n(q9�}Ȥ��t[�}��m� ΂��1���e��L��yCTF,�D���s�Z�DE��l����Z)Î9��N �K��J�v��R��hof"xM3Ynf�3�:��Y
���Z(��Ŝr>�*rhW���P�+WߴU�\�W���T�Nj�~�L��F-�;�M�CsK�/�4�76��D.�L��bo6\`O�j�hD�6UN<r�9EQ=DC�����@6��^��'�I4ٹd�xGE���,�aIH
�Y%����f��H����<iG�"
�zgֲ�mEpW�f���q�"(���K6�ʫL�ԯ!z�dY�C�s��3uw��r�bw��`�-����nq`�I�W&��5	���}v}�����D���A��=<����a�q����'��pQ���(�V��{��C$��HC�:����a�����ױ��䢭2���:od��3+�Ȥd���<�g[D���}�$���y��
�A5u��&�r%�%ೃ�h�/A@��U��3�<�[��|\��-PEH���3-E��6���+WD�U�O�)�7�����5��~ ��O*��Q^���D{�]Yq�D2y&5��?��-Tv�կ�� �;m>����p-��v�ɉ�rDZ�R*e·��2~��d0{�/)7���+EgU����q����c�{�C����3�5��&�&�W,q�K���?tL��v1Q��K1
�h�C.�7^��PJ�f*:x��$d����ԁcͰ E���y��Q��CEG��L�n ��c\WWI��
�|�!�d��t�x��W��G���"�Jq�Ƙ��;�jL�rO�&�"�����m����:����k�S_���b�͟j��Vq�I�@	�Y��������
EFI���\��2�ygXO����.��<直L��'�^�[1��eǼc,oWbځ�I�8���h)�4���Z&�D���ga��dͬڌp�J�,΂�f���:�*�Y�M��Ց�B�ߪ�{�$���wQ,6�'�~��������Df-5���f�k�9	ɠr����VyI�%�:����������:�� (=nI߳s�P?�r�K6��L,Re���o��WYN�팿y��?��$��g�	��\�����
�d1����:Ѷ����s��w|' ���qj�U�E5�2�T�q��豖U�1Y��q�����>왧���J^��r,�pR��Hza!���Gqz�5��!�.ڽ�q���������E7yp@/��_�M���Zn���qY����[�C	3�<��xM�F�נ���U��D��V�#u�ؤS�m`���&����m�g�e<���u�'�kV q��)��A�ޅ�a�v���X�d|`D���6�7i�μr�D�#��~���죾^*j�d<U�" ����wF�����X�N�'�S�9X�m	����!�\�n���aD�/@U�@t���/8������3�Q��7U�:�#K�`|�M����Fa֥�w���N��U�=k^�4H�	P�З��
r��)�Z��%�]Ͷ��\W�|����KL��G����L���Ԛ&���e
� �+b�a�m����r]�֑��]�s���m�wJ6��N��.��B�k�	�U�BYx��<��R;D��N�7�a�� �d�Bx�<*�V��1��48�V�Gr�O`����'���z>�� �0�A"0 ���>��5ͣ�wpI�y��:��[�WtXhV����.Cܡ��ء3������|k7`�|���C�� ��)����4jhH>A��JE��o�þ����<�%���f��MXEvRo#$ۋ�����~�V���Ù�6,���:��8���U��ACe����e�c�Ĕ|�_��.��d���s;�c����C�-�̈����m�ww�2�|�N�'�e�vQn�\���:4�vh��c��a�Ek��$A����E��7�tA" ��ߑ����ǞE��;��
 ��A�
۫i+6��7p
�i.����"]��J�S~a\z����5�"c=�INS|���̑(c��V3�O#�8����,�+��l�bGAd���$Q�tEʋ��@.�!�0B�Q��A���\�I9dPN�7O&1�x�`ۢG����t󔀄B{%Y���-�x��O��>����M+�EFzK:N���o�����k��۴��Z���\�	av�c���uc�J[���rϑ)}�NE���N1B-T0$j�j��>��M��0��)��^��ڢ��ǚ~������-А��͟+�/��[B �KѦ��t�߶h��:����� ��=355��'T"T-�ʅ�-'
�.�k�1�.�*<����3�7���-��<6;7z�ʅ��wq|��-"+ɍOL;�[�z{G� ~=%��I��8h	B<��F}r|g���s`��S
�W�}@��ɯ"���#v[�b���}���e��ʇ�aگ"�C���r��l@�T�nʛ���M�S!��;m#�bd�=ml�<�d����%̼V�?��ԼZ�#��G hk1�?��X���]�/I.�� ������|�Jyv�n5�K�/jc�)է��:w�����t��<鯶V��Wt�_2y4ȇxFYѡ�� �7�5��b�R��8����E��������ǂ |���Edӫ��ej�ː�6(�<����J)A�F�8����G�ո6�S��c"q�51i���^>O�\��\�+L�-w�0RWEI�#Bl5��y�T�s���!�ձ��t~����^�)7{����Ya%�:Y��L�鼰֣(��I�bl�	7}��l6���"�����X����A�r�uO�@���3r�׈�� [ƫ7'xQ'qM��h�Ӊݧ�Z�t�||�,�f�{�p=P���M�`vE�/`�p{��Կ�`x�����
/n���[�����&�G�}��4� ^�{u���I���<��oV?	���Y���Q�2!�b�aD*�⟸Lr��_z�@'A2~!���D����8_���ͫs�=eE���Wm��}���hL���,�MK�x�.L��&�T#�l:�8\;-��kN4�KɆ�L��PŕfeH㴮��k�� �KN��].�mR�Ļ@��=��~㢛T�d��fk���C�N%�)ї{�d.= ���=��t>�����)�őbB+�>;��DVu�~o}�?��Լ��<��n�V�t�l^�Bw�a��>�ـyN���n�S�M��ϟ�R�t��C��سQ�^�>[Q��S��6&noƦ�m��\��B�5혠F��v�e�p�k�!�bA�[rs�=��^	��uB�j��� W�h��6�lK�Zͼ�ȡ���7����&����鬀�ǘ���,-�C�Z��-�^�tx���e܉���R�Kon8�Y�EťǗ�	~X:B���A�ƲkPW.��S�DA`;�Q��α�8PT���=�5s�{F{rT	�ܞ�P�;cf�'c���R�iͬw�6�I8���(9W��
|����L#���p.��.�t/Ώm���[�'<u�Qd>���hyJ��{Օ��a�݂���e�_�����ҏ9y �첻�St�	o^F��ϭSA��D��x=e�&l��QY�m�&�ڂ[*��0��w�l�k0CY���2���_��L;y�T��#���~�s�,���R���Vݣ�����J���V�-�|T�ȇ��hOo��M
~�Nm�#*H��7�Sʎ��~�7�sg�9��v��4�^�K����Y3�A�Neˤ��J����Π��ԭ�<�g"/�vCz�W|�Kb�PCq����81}S���I��sP1��-���`s	��/�����&b�/�Bh�z�����Q	þ�3�:�H�r��!��Q�q���c~0/�V��os2#��������kt^m|�����}�5#��ӽ�ZH|��@X�8lͯ{"C���Q�Y��f�u[�n�˴Ϗ$��6+�B9��1�)`i4�U��������Z�����:O�yR7���?l7��G\\�ሧb���� 63�"jq]�D ��vб�{9�M��i���2`�e�ᚣT M�$)y}����STN��cS���_��W�Qn9`׬ű{U����{{P.O��������'�%2啜���� ���ܔ9������6@�'����7��$G�o��$e*�()�vh��8_RAj�}�A�砌���̕S,C���5�����uK'��N��dpN[=�n9pݽ�����Ҝ�6��M�<���"y����0!�D�g���sSZ��ѷ�R~~GO��9��a�z�Ce{����z9G�GXnR�=�@�
-P��`�\��s��ؗ�O��j9��l3h�r�߷��qs�H�Ř�a&���lwr�N=��� πc�O'M�a��Tt��6nz{��@펞{�m�D�Ұ�kѱh��i��5Һ�Ns3��
���r8�T��Ճj�Kt�x�?To"���IzE���<�m�f�(){���p��1S�����?��>�[�f=�>�{�`7��3Q	e�.y���`'��Ԯ�;������7���O�fyU�&�bC�^+o��S
�=#.���ry
aǎ�R��
����¯�t@�B}ȳ^��ft�\�Pɪ��F؈��Z����£9f�m��EA{�����z�&]��uY�!������.�4��{������Q��$k�8?��W��ߕ��19o�%��u��$���?*�2ZB�*�/8��)�X�b��Ҋ��J	ʧ����Hb�g�v5�]@�*�v���:Ġa�:�����+�E�_x|��|e��bL��GT��^�$TT����c��$��ް��7�/<��=&	��#H(4�꧓�KkoARU����Fr�Z���z&�ڸp9�ܑq�{ر�6h�͡0^��a$;J�)���mY�N^<s��k*N��[] �,a�zv�,��k]��<� �4�1Y�����f0�c���qf�R�� =#�w��,�&x}O�'�}�)>lʨ3�ܫ:���yo��3����4�-�P�Kv�CAF������T�N�ƽ����Ñb`!%�H����0m��rr5\إ���M^���^'a��ط�slfk�<a�{#�A��� ��\�c��l�=F�$���=�ژ͎��#f�/��:�@:�����k�Ή�Ҭw?�z��aD��W��N��F����)G����YRW�R�[�>!��e�`F�iB�V��1|�=���? ؼ[��1*�̸��4{G��r����m~��w�W2��gf�;�_�d|N�E��h溂���dj��V���Bk=f��_�i�=ƾ����;���9���E�J��(1����)��a	��V�dU5��c��<>d ��"�Z�£�'G��&�"�;G������~����nA-��z{��H��K�
֋��5X�;�LJ	~C�qnu�̉�q
j�Zķ�/��U��������	��Qe�*���x�m���|}�������:UP�n�ߕ�m��[�x�z@8�U4�45���"���'k��O懶����R�2T�������Ly�H��o�O��?�V��g*UJ��?�����<#5��1�xEW��糟�}��7�9)�*�����$�ܽܩU��1n�!P"�,���`�Q1���%��J�ol���*+������M��H� a�0fM��x��
�zQ﹉���*�=�TH~����M0�^T&�f,֙�m[�� �1�~����"*�
Ʉ���49��fl���/8Z�d�92���n�%�`�FK�@�Wad��v6i�)�yi�nH(C�Cn@�Õ��fgDH����&�J��8�%^x����R�z��B�w��c���\���P�_n�)s���]�j��>0I_Gd$�.M�GƆ��\��W���R|�X������:6�?���*�]��=�#%�=UQwf�*
P`�/A$}n֫��{���{[�:��M���R����o-Tș���A Hd����t��1�*�&�@f���Ilje޸gt/��M��=����I. �=�z3�1?r�@V�97	'�]m@S4O�
.i�[�6b �G�n{�xg$�k	�-Ԫ+3�γ���Ϟә���&�MD�J!������5�����jv@ǘ�mǯ\��R�NYae��\~��hm�3�!�;�iVa��k���Lfz��T�pȝ�J���,�!���G�tV��+Q��h�X�Ȣ���B�q�6DV�u�6�I�Fs�ٔ?c�����G�
4<j���[�����bk���JIe ��M6�z�����p�n|��_\���RG����񴪜vHY�[my�t��M��v�2��x$,Nn�p,��D�3"�����NM�7a�9lD�|튈x�h��� ��ҝ���k���l�%�Ֆ�������0�W��HX��l`���>f�)�iC��u���2���mO����/���x��cx�%����W�x��Kޗb?�.���5/�������Ѩ��I�pO�"��)�� �!�{���da_��h�si`�u'I���
�C�v��1*S�gb����<a|F��[��:���
�T�?~�0촴��ȫ�U3vL���
�{�K��9��ǣ���_�ʌ8)�`։�k�����E�K>�x4P<�#�K�K7��	Ű6�O�I���D�TI��9��⸚\�E��^?dW���n7�(\ǣ�� gw�Ξ�[�4��֛�g\Lz�J�7���E�]���7Ԛ��@�D�T�	yBxP�X�����
1��1��N�X����n��K��:�e�˟ή�*ń؍�w�e�hu�:� �SM)j���mξ�X��n9�DA��q�&�0?++���9z� v�G�"z� �(~d��F��P�G����;���*<�p}��WF���u	��6ߺ��OLҨx��n��(r�ȫ�V��_?̱n�&�cR�4�R���O��G?�̏Y����7�|F5�%�lcku�=^�з ��a�k�rD���p�#����Z~����-�T�ĸ��>g@��3�E�~Æޞx2-Z���p#�`+��GЊ-(�98�\�IW|6[�3�sO{���<��=�H�B8���tV���i鸘��d;�-�?��|��N����۾9:U�Jm���@�޻g� u��!���3�e����YW��:\��@ͼ�J_	Ϟ����C��Z��3?m�	�#��r\�}_�E:�FB������(��d�R�25��#�*���X}_����Z� s�$̉�@gt��,�&�
�1�O�42�]\��~T����}���p�{$�d��KЗo2��;��ӯ�EdFLORY�-��ɋ�I�w�5)]��A�Oz4H;=���x>P���)�m(�e!�� ���2���8_�W'�-��$4)�����\�8���H��zJ�E� V~M���^A�Y�oT쒏����/��{�j��Q�v�@L�̒-/W{�m��X|OC@�x�T�9�&k�4Ҁ�??�&ޤ�������+�j����)AB&�C���|O4�c|XL�$�=R�8��<)����Y�oA�W�Ǜ?�1&꩛�B1��P!�a�KX�'X�#_�@D�������d����� ���E��^�����v��tm�>��n��<�Dq��<�A���K�*v��K:������&��@H;ݤH������P^���:�%���W(�/������l�:��eUWN���j�^u����_�)��z����@c�ӿ�K��*[�]q�"A!��JK���'���_Dl�':� ��d`��}�g�*Sur�l"�ā�.�L�\5��:��a�����S���<���Px��(��Ž"R�M���- �ɷB����N����F���l 	�� E��ٙq���~5�9�o�������
f�-3Y�T�?,���;.�Q$L���(kh���o��?B�j����uv�HӒP!?3u��3J�~�p��z�i�}R�cV�/�~J6ѵ����@I�����N����-���pb�汓gt�vQ�	��W�.Ґ�t�����ڿ�lZ�o���%����Qu>PB�>>HJdQ/������r����uݶ��DQ3Q7�׾޼�'����`��i�kC�>s{'vk>\sfi��)������"qb���
Y��z`���+�ً��Z�Ă�`��e Z�z���]y�t ��q��~�X�����\iz������)�jP�s9h�!��*�J�=4K����	�Ǻ���eLlD]a���L�Ht���ҧ�4=S�����MY�����0]5����x���,V�>��2�i�0o$������B�� ���aew���Lh�=�UM#B ���lAW *�cI&\9��W�;����h�&^�K��HJ�?#���<�����į��g>�\/J�*���gK�7�7��<h7���D�e�KT��� �qU��kIT� &���N��� ����>�-�a� ~0e͍1;%GjU��Z݋v�+|��?���;C&S�n^��oo�
�\k%{9m'6u�5�C���t#Y�=~斮\:����yzb*/�D��Wnff1ū��W��gw��)������X�<�ۂ���Z�[�h�1���{9����^���:��ER����^��,���������Yj-�>nރ�'��!���
�Ki��t��y�C�Ë�^�~w���������:��K�g�`1��7!�Ϳy{Pw`	����!�\Um�X��}�y(f��~��Ǹt��H�M���@NtØhk'S�ᡠ%8�〛Y�1�N�\ߧix��Ǜ�lE�S�Lg=����qb��B)��KEL����D�wf[���E��R6h_��J�����t.N���\�q"�"�s.��ͣ-1�"<q�� Z�:�ޜ0�u�_�����ڱ�ıWͤ�ر�2����zbj;t�l�$V3ȔlX�V�J>(έ��4kZ���[��C����!*�v_�Ika���$I�D���}$�-c�#�CǙQ-\8��ߨMv�q���� ;�����+Y��2�Q�xE��V�g62�^Qch��� D�����N��l����˵hA_��eHٞ �k ��(2@���, 5#80�od�^��pw:~���䜁<K�����cm�PV!��?"�*��`I�~%y��k��k�?�5qC�O0��Ӑ�������L85WFI�гq��:{�JB�ǚGAd�O�b%V
D��=�g�V�h2�#]����w������!7v�����evRL3	�/4hVo{%��rsUR *<��>gs�x=�z�Ё�"" ހǤ���K3�ߑ�:$��Xe��_�)�R$/RΨ�#,(�A��*xݔ��){:<N7���1�\<�I����r��@��ؓ1���:��)��x����$��h��k��fԦ͢#2�*Өi����i�r�^Y*%o�@u	�m�9�R���D��mXv��'D��ӁSi{�_�_�I+�wo�w��>�,X�����!&,b`�a���%f�^[8㈺݇��Sg�ԑ�0-'A7�<��(#�Ӈ���aޢ�{@҅�InRЛ1��٨���Ҽ�YR_�$�y����,٠��~����4�Y#� m�O!��l��+�/�>=�D�A��k��[���տ%��h��=�yD]���Wx��ܔx���,y3�?g�j�6�t���%'�ң��~�����/* ֢�����//Ty6"��us��Bn�y(j^��xE!��+S8���D�Pst��*�����b��cP������'�Fc��+w �-6�uz�\r��.;�c�ǂjC�&���mq(����y��>P��PrP+�Ċ�|�\�U�I6�Ry�� UOjy����FX&obͼ��o�����I��%�V����
ʂe�F��Q���_6"[,��rijX/%�V��N����q?���ov���ex�e�s/r�x8��vZިf
W8�'F:~9ml�ተ.F�Aڭ�K"�1DAm`k�Ҳ&�D�W�bG~e|��S	s0���'���FpY�I<-<����<��P�j�}5=��_J���uSt�qٻ�6���d!=`�+8RGv��i�9G�c.��7�����a\2)���3'㭦���mЌ����F���#�����Y�x�y>�c�N���4'(�=m��l�a(D�L��-�%�k�_D�[��u�
E�^���r�R�Q"A]_su�g��a*wWr�:<v�n�t�GQ:�)�r�l�F�8�+Rsi���4����:\Q����:��NY� v8�;��{�}/Q�3�I✇.���L�(�R�% B��5�̿Z��TrT��uPqN��;]t�y��Wa�r�@�� �?Jy}��ی��+��~.��0ا��d|^Vx��9IU�@ނ�/4�9�=���r���f�v�I�h7�g�&����p��{C0T�_#?�ө����(�R�s#Y� F\�o��aY.����އ4i��C���2���,�2�
DK��8�U.��a	�q��4�nP��j�k���Jl�jp���'�Tn���� '޶�-WSө�	�V 0V`Dqk��m�Z��~�9����D,i.�ǲj��?��_������2��kA"�F�4ԅ��ףoTE�ۥ�|ؚ��X{Gy�<�;w����j�6�;�42ڳ|�@V�3�t�J�'�pRE����������o��N��Q��p䴘<�*��kӘ�R�����,���� �2~֩@£4��O7!0y�̰�s��8>�*g 0�_�/�nl�9U���.��&Gƅ�����+uA�v�ax��қ�ǡ�ih����{��(��X8�*JUO���z������S����q�𰍙�eC���(��Ev���"^��?�i��+!oELy�
iy�l��r��a�L	�X�wn�W�n2�b%�Vdg�%)���n8<�ν����@o��3���Ɨ�^ �����z�P�mn���2鸭��3�'H����OG�#�BC�!@!%6���0���|�����	<|ex���j�$�%R��~Ȇ'�� ��A�dRp����r��7��wnՆ�/�\���!%#�~6B���J��n��Aɨ4Rv�]K��G X8�t=�p�ȕ[�|V.T��9�����aýi�j�C��0�!��8	C�w9Ԣ�V5����u��%�"�����_�,ڟ7l$�R��d�Vt� ��İ�+[���PH��+�e�Ch����6k��荀�=QhD3]ʐoT�S��v��ԁm4ߢ8M t�Hw	w9��܀ƲM����0S���V����U���V��+��F*�����#���er��'�E�	��0��=��rԤ�������]�;�Bk� FE����&(�w�T�+BS��&�d���qwY���r�sGT�
�+<rRr�g{��B"E{`ۂ���L~!vvF�h)t��� BJX�����M�5h:��4��(bU������!��i��L*��2ff��a���R�	 �����z�Q�2�*���>�HaUrl_8v�Uڠ���Z~�@�}	"�8S�Um��9��r��͹_�%/E�Q�����^@мx�����>՗'�)b�=���;�*`��&2( q����B+�\�m�V�些�����R�g'�G���R׶0n��T���H�X�.�j��t}c��l���f����>y��nQa�� 7�!�l>b�3vw^�E����Q�qq�F�n�H(ib`��>�'a���:e�3A��kQv���<\
wl
H���R���[��uc1ĜC��-��-�[�} ��7L�����zi�H��8\*�G���`-�hym�{�?r����B��u��!\�_B~Þ�
ÉB��w0΂�)R�q��������K���v69x&���;	݁��1�A~&�L�]����7���ml�@B9�(o$kdQ=�S�����hZ7���_���i�pI=\kmן��;��ܶØ[$�{����ymF�i���&�w*�|r>�S��:]��&q�����k[�%SW�$뀚��oE~�����U̓m��,:�ݰk-
'����~|�F"�?X��Ԍ�&cO��+���*��)��SAj���Y���~?��B���j��"FE]�4Z�������H���w���� I�tu*��=4���ݘM�.
BV����*M�5��e�w�uS�J+�Q�&�((��+r;�"��X��3���t���D��R�i�<�xXA�ޣ��YJ���8�߮.5�5�E:�!H6��}�g"�nب��\����~y/-��,�N�X�m$�X*?�'���K���+&�I�D�]޳�7��J��cT�M���m�ɗ-�?sQ�����;97���s��S-�4;�Ig�i�]��&���w���H��uv�ى�D�S��qȞ�b��$�d񁕪"��N�%*3�P�.����lY�͗A��C ���5~��<n��?�ojf��O;䇐w���%~mK-���"�c��CA,k�n�]��=�����\�۶1"&#۝�!�˗t�읶��������Z��-�^�n�F�j�)i�+Y��W]�"��u��^9���ט^�S��vp��J�,��S]�1�ACn�~��n�����՝{��0nz�;aL�l�?o7?}_>'C� .�8m�>�t��]��t񖘇#�mY���&�p�l����K˸�.�Z��-��)#�����x�o4+���yID�X`�/�IB�-�N��¡]��l�.��=�'�t;5�xV5�b�c�ؼaT��wBT\rޫk�i�i5Zrڂ�gF_�C�mڹA�I7��q*�Ey����:g�:O�=|��2���	�p����	���L�5�wɽ��i3������cى�'�9���#��<}�þc����8߽ѡ(�򎠷�^a���)��.�@r������T8o�c��O�5�*SP�:*��~�㻉9�9K@Z�j��:�?x���x.��M7�I�B��ƍ#�c{�������B�R��	�[r[�B7�T{�%͐�@���aqM�dU�RЀm� |�6u���fMg�"�xٷo�R��������Fv��!�5�|�s�Z/�w*�C�ֹ��%e�xމ�ς{�0�����eh�����C'��"ۥ������0kG�����!#4�F��pmB���}:U�N�i�'|��a��.�$������n���?��?���ƻ����wv��e���QN=�O�2#mp��:A�de��e�	�5g�&�%�}��˙k�H	�:d��o���,��{�
c���u;��]����Ô5f�	/I���i$s��J��^s��Ev�Z��Ԟ�,>�J(<����"��`M+��IJ�`�j�G��*^4?���\�s�(���>HE�fM�Jd[BQ/�H�0d�L#]�����2&mO�ju �N�d���\�9��-�y�d���t��%��Tϻ$�k��9��F^f|�T��8��|�-�N�4���\H�ȯ�MG��7blc$�����2h�l�h�J����B�:`��~�j� E˾5O���+{�"���b�kuazɥiU�ݹ���S�|J��t՞|0Vu4���3(�RN/7��F�cwr��m���3�;�j.t��*)x$��%ʫ�BW��'�	#u�=�[��Ա�z�Ș�SǪ'�e�C�����i���@�=��k͋U�m,HK���9�
1�}�:�̥�o"H2;���u��������S��9��.Q/�yѴQiR$W���HA��ւ�%���3j7��w��eL�����Ԇ.K<�Q@��=�l:wWZ3��%�U�8���Ȕ�@�	�kX�C��l�{r ��nx��rW�_���{W�5�DJ@~͂�!�fMv7��!�⳹�m�{�(�:)!(��X�*w��X_��/hӭG����+���8Z9��Y����%��U5�+�N75�y!�q?��;>b�}�{FG�!X���=�Ш�0"Zj�F���y£��#mEx��/�z���@���#в'�`�x�ZVr�@����ȢbV��ﳂ��|\N
��`���S�ȅ��2��0^vi�!ERw�+K�J�\���&'��ŚҨ�|�|G�I1�d@�]{:�~z�Q�J���Ѝc��QT�UP�ڨ�VK]kk�d�V�����Xw��c�[�\]C.�@]?��R٫)��\!��ԏ��E̝�l6�����O����#�3�T�%�;Y���i4��߄䰤�d���B��ْ �t.��O�%ټ�4��ZI����b8
p<أ�x8�:PX�sB�_>f�W�j_/'o��·Ɨ2��� �dg��X���u� ��X�I �iB⼖n��eMi���_~����W�X�X\.Z6����vuɹ�n����&��4Ͽ�hGc\Ҵxɣ祃o4�,��T��ƞE$-j0B~e��2�@>�z�Nyy7�}ŉ;�5!a	��ʓ1R��iJ/]�@����G(�#���S�j�+��>�d�s�dEJ$f^|�ɒ�,�<�^��d��^��$&���$�Q����y��2a�W�6���B�������>��I��j�U@����{�Y[��>;Dl!!�B]��Gt<��_IF]8��){�2	[�?����!N9�����:�="��;�vGA$E������N1�t����̶
�'wP���Ä6۬�Y�)L�B�����^��b�8B�����<P`�r{^���}nޞ�E]�L�N#��>ugN��?�a�]��z�֟���Rp�q�o�l��䠸�9gC>�O����}�+�L��Ό���E�}��a�rx�WhDaE�#�i�%V�2 ^��N�T�R��׽,�X���J!�_��)Ա�͂��$h�	c���ϛ�w�9�&�!kr�þ��[)�u� 뙬@idB !�`"p�Lr���^&:齙����ث!��j��"���~գ����[�E�ܴt����.!�͍����hfۈ������KQ����9�V0I�ݓ��f$���0wae"4>��~�[����4|r;��t1�<������� 3��>���WF�P�/� ���si����������~�bw�]&��k�6`�^��-c5x9�pKi�&ܪď G� �M��
/�Y��:�,��k�CǿA_{�k=w������Z}���hx�~	�v�P!�zT����5���������Z8�OF�7iz��l���J��qH�5��A葅@���%?D8!���J��2�6�:�D���)�!��3��H��zK#��/%0��8-.|y��_p@zG�T��@N+!ͣO��nK��w�^~��1~k,� ��I0�?��p)��7U)�f�J�U��JJ�i���mt�.��tm��Z�tw����Y��p{�`�L�������M�ڣ�������UIo�5Ɔ��J����>�?>9�Q�M�k ��|� ��0=��DIT!I$a�l�6g�^3���Sl� R��#ǆ��h��A:4�|MK���8Z�`<l�$�c ���w}�[�ٟjc�dB�v�-�A����&[|8���: "�ژCC�Ih'i���������'��R$!��M�d��Z~�����Gг�k��-�\�geҫG�[e��/���nVSI��¡���Em��UL�OK[S=��d�t,���xSwr
W��ںS&ϰi��m�s�c���v=�H� ���\��$LHa�"�! �X��ϖE�U�j�1����]�"�x2Qu��]|�q���q,zP��Z�*�_��j��|5?�v��Nv��ښ�:�o���+�Q�A}��%�9c%O�4^�1�������	�2Iߦ�<>�_��u� ���<�����m$��Uxr_� =����F9PF�Y� �;�Υ)��^�cѸK}�b�Q{5��5xP����@������� ��^'�?~��ShP1�N.�Bm[?h��R� 	���3-�y0�6Ŝ�bD*a�Ŕ���n�._�]{�]�iR��a��I��4��H�a)>y�
�8��M�SWNgo�
5�_�f�&0���6�c���@b��������;1�V��^�9�Өs���f�p�wrk�9r��h+U.V~�=�)��Ͻ�{�סo]��W��� �1�@~��8��TT0Z�е���Pc#=;e@��	ǰV�oi�c�G�X|��E��y_���޿
���a�}�mk.�����t�M�Oi�?J�M��L�Uf�{���{�N�E��� �2n��JY 9�Jm.u��W��9�q�{����� <a�㇑kC�E�kf�6��a�=����`��D�'>�����PP8CR�k��$�i�è�)�Etq2J���b]TU�s��/��bc1�+C\j���)�-�� ��7:����FS(�ٷ��%��S�m�qڔ"�l�I�Hl�g�|=Ɣ� =�b@��I�}t��u�I�R�0-|� ���%���CɰJk�<�R����t�f����0
ꖅ��]�G����+��U>iָAl����_ؙ)�^�F�|���㟮^�#��(�d�ߋ�I�`̴GI:O{�9`��˚�R���=�w��:|2���Z������.Yʔ�qu�E�k !�;�n>������*�zY����͆�*��NYcm��;~�]���Xϻ�����X IqAx�R/y���S���<��1�r+��v��6t6�9���{u�4�=��X�@5��ꆄ�!:v.�Ӓ9.
t�^I�%��v�vPOcZ�b�7�J!
�_�0}�D�<ɘ"[K�T���
����=�tq��W6�jɌ/l��ۿP�vj����R����]�t�����ie��L�����>o�ڧZ��Z����?�N�k�̄��p빥���b�����id�\d6�	˹.ߗ|;��3�^�	��\�]��ˍ��s>�����)JY�!G�x�����a�qmߠ���g�1v<�|L$h��«��%��n%�.��{�:��!sɲ�8�yY�OInh�]l���͞?d�p>U��:j��.y��z�`��-,�]x8�3� ��p��<.��sg/b���i�¡s:N��T��z8�
\�z��Q�{�=�>H���K3�H��ڶsn����� ���NE	��g;�/�H��T�so�������7r s�Z�����Ԕ�Ob�t��}$bk���(��_�gR`��UN��Ζ��F7=
=�+�:=h��x���Z����A樄��[�?\Ƭ������a\�f��G�S�ܷ7b����r��=Y�����=!�Bܳ����r�'Xx{��X/��:YNb�p󀻲T�Ƞ�Ċ��u�R��E>�\s�q͕J�I��eƣ�#����:��8�Cnؔ��ֿ.%:O&�V����Y����a�@c�S�WR;B����(45�>���N�]�5�K��7���h3�թ��cs����j�X
�	�������9�ʌ3Oz��[����<��XA:-M%�3@7��!����)=�� #?'N��*�1Q����&�xF$�5�R"�m��r�r�b���m��oRR�+7��x��C+�P�V�|��c>���hb�8����|��n�t���J��;����D��߳{�c�;|���K��B?�z�B�'G�9�pv��kt�l-ǖ�łS��yP���� c���%�3�<���Y,��j�w�#��F�"A��r���yٻJ�J�5�Ǡt+D�-~�-̐Ƌ��=����`��b��b b�8�dDy�-�ؘ/�cFOIܸH�6��N�����D�����Ł �%��+�Ɨ��dݲpec�#w�/,����=Ƞ̞�#_�j����9�]\��m3O{�ԫni_�n�g�FzzI=G�7S����O�-�@�I�;{1�����K�"ís3L#�k2�~=��������ǯ�i��;��
]�O��*(bb�^o _Xa1�5��΋��IUF0�)O�y�O���(8`��[,Y���z��3m��'��R�7�+����s1^"v3������ E�vm6��-i{��R�@�ϡx�����P%�C��{��Ρ}/sمh���}�QP��6ӏj�3���[�Ui��O:���B)�F�x�#�WEu-BP㶩m�Ã�g�7�PN�e��h�[�e	���U���VF�A���:�K�p��zF�dC�<8�I�C�O��k�Aש�s�f���gSX�_�~�l/dp�ً��������)xB��=jR��{2�MW�����AE��:�QE��,U$1�z�t�>�a�.����̺r���y��䗛iq�;��v6�������'�����%�y4��#���T�\���@��6�5��rc~�-bL��%�9�d����T#�Bc�ō	u�
�~�V�>}D��3���K�8��3�=d8�ۑ��%����{,���>贘��fZ#S�K����=��m�����G6G8� �]nT�X�+"�4��؝N3��R�u�����/jL�C��r��W�;��3Q�k:>�~ˏȿ1`��=І�Q�L݄�N�t̉�9�Ɇ��Hk$�SG�c�ENP� �JG��-Z#����7���-i-�[�#9}ȪF�f��f`�>�Y�H�%�gf8�Jרp�H])&O�Sp�aa�aG��QZ܂��в�q���9�MCP]?�z�=�v>n�'�t��B�����O�����g`���S?M��u�sց$��)'(�`7ZM���7�R�㲐�Y���-ߋ���t'=�Ԡ|�y��o���Pߌ4/� �A�|�hs�v��ޅ� ��,���b5����ĭ�>�ӄ��1��Pw�>?�Q���zj�"�����} 	���yV�m%x�?�0~��Y�sB>p$�DN�tG�]��	�È�I'�2�6�����Mdu�Hw
n���(��{��>1jc���	�\vo�庽֖��P����)mF@�[~%��6�l}���l&�:xf���ؒ�{4f[�d�μ�#��|SS��?i��$�კ�s���L�AG�$�4�vXk�{��k8��©X��{���|$�Rho�\�Z-��cx��ִ0�?���,%t�X�5RT*��AV�"�C����n�H�G� T����X�7m*�;��(���6֮���ʋ&���Xw�7�yD����+z\?Z���Y�83��Ls�K>��e��_^��;��/R(�}��݉�:�:��o����̣B�b4����S����h���o�a��	;�о�n9�K����II��e���p�Pk�g��1sy]�d����T�4��������T"rG{ܩ9����ɋ�CZ�����y��er�9�4��Ǌqp^�c�f���d�pѢ�Gd�.�K�M�:�~�|Ro���lj�uy�!	�¢v�{q<�/��#�w��7Q|����$���_\���?�ȅ��� �U���1����h�܈P�٭�wa�;bB3��D��BV�je��l�v�$<�l��+G �E֯8!��C���#��R� G��uM5#�"Y�w�H3.E%�<� ؞���!��l��_����F<V�/MN��<�ɰ,�_�B�2�zb����n�����	f 12���RKs?�v��k;�Ew����]%I|�)|�W�^lt菺Q�>��{��Xh`�=?���'>��L��iHWą� �o(�:�`���I��Y�)��x(�Z�z���2��^�\�H���S�+�_����@xhf��%	�����ީ�]�V\�n�7�r���c��תs�\ٽt��TR�~�!��JU��7��{�T��Ys5ۍ�_f�
��[�%�~2m�X�%�j	*�ū[��$�E1�`t������o����eU�W��������ByevRz�B��K��L�z��k1)��GsSg����ܧm�����',=2W#���&_����sM�� q��D�V�!·��$�	��Ww�-��̈́�#g-��@eBI�^��b��h<*
���,�!������+�ga((1|.��G�� �&�0#p�~�*��L��/P:��L�?�����iV�	�wLcҶ]��4��7�����|�e��I�K-��v (t���H�iv��_����#j��K�qlۥ�b�g�?���_�t>�P[�zt`#�����l��,����6��EI�}�s5@�ꠒ��*F��^:'�tB5:�FY���D+W8.$k��qM���6��޶Є�-��zB�`�^����zGN)w��\���tPHp#~�ʴ��`��p'���N
4����2���N��㢈��2T7�:�H2-u����ܮ��|1pMS�'�ۙ�+�Nxp�x+���l�_ߙ-�����4���������H�z�549�.Pq"�^�研kwCK�k��zt�+�ʥH(_���͑��=c��W�L��KJnc��{n)<����i�q$k5E�Cs;��\�fm�%�('��wZ#)���{T4֪@G��֍�i���
��; �}���ӗ�P��)<�@LE�3ҸOLmOЃҢ�|;��� �!�$1��.�S$lb�8�h�#нtoߕ�gx��Ļ��Q���ֽ���EsfD�q�V,�(i�{t��?Z��\j9�p&������ #��K��!{\�������چ ~-ݗm�0T�/kw�'��$��N�[�8qW<#�@���0��3u�è��wk�F�¬���/K��e��=#�ꤲ��d�%W���pdL������Ё��c���Y�w��XC-���ʄ�
�k�wY^	On�Eqa�UFA�ծs�@����ޠ+�Wr���&��eb\������ދ��<�
�w� ����	���:h��jͭ�B���H�;�b�>e�����ǮF� V�8�-���|
g��"P���ǩd7hY��1�.��mMbN�y���KE�_y��
d $#���E��~6o�+ �F���0;�cp��(�̐�g:�I�Yg��\������������S�t�vn^�)���6 �#��B�_�,�����A�a��-��� ��DH3�K�l3�!Y*��Q*����/i�8�ɟr�����[ �@�Y_����?ʣ��c�t�����Qݚ��@�C�\HM��1���x>���]L�[:�ԣ�?�h�k3ů	�$�2}����Ϛz!�^c����0p1�x��{욲a��w����ݮjf����w�U�ݺ�0o
t� b1d&s��wf�Qhi� #D��*�*kvû���IZ?�����]�O�:8N�^U�b�啞_��1;�5��D���e*�黨&�kVEp�8�+�J���S�׮Z��Ǘ@���K�V�:3�/�
��[#�9^�]��W'q��eKVU.Q =bd1���4I��F��%k*�� ���4�Ma��cd����S��Wwi?��ґ���X��J;sK��kM5��S.��^69�}������um��otd��w.��\���$8���S�q���Ͼ�-ŏ�L�)�0��ɔ�Xx�MB����܈y�Z�[�ϲ��;�,�H.A�yD�ZӠ�X��N2�^k�#�t��;���Am��yT%�W��y�Q� &t���Ǿ�H���x�Su�\��NW3�N�y(3v��Fd��R�,�et�������δ��
Q��~�*���!���^	RՖ��u��j�?�ɻ�l��1fV�i���l�z��l�cV��u�F2iIܚ.gNE��<؜Uc~J�G.*��?�=���n�u�0=�a�͌e�����̷�'�=�#~z��N +��DN�}8��26���I畄m�mX�H�.x�L�˙ǐ������Ĵ9�bA�Ñ�1eߵ��2;�J�(�n=uԣ��� *����tP�mu�y�~��,�dNw�I�m
��������������=4��u�@�c�A!���ۑ����J���^Eu��p��y�g�4�S�w�C�~�*���S���<	�^�M�)�E�ξV�����zxP���?$�R��r�H�n흀����e����3�#I��s�Cf0�B���_[�p�tHc!���e����dd����%�_��0�|]�s�4K�g�S�����g��]��$]�h2B�����N�X�E%�&��o9���s��Xcbۏh�>��[S�]LF����M�Oo��J:���,�L�n2;�mG9��5�u�З��	�g�M7�K�l���l�&���,-b�mhʁ$)�?�4�����L>�wJ�S b���v�l�>ح��[��FkO��ӎ���߲�%�@����]�5<��)m�[��̓@��"�/�!˿I٢�_*�P��G� �uU��2��PcO�G����
:N�=[���-
hQ��FC ����s�j^��O�H�hTȲ�=�й�Y����o-
�`�U�E�Mᓉ+� c�9���h�7�~O_���gx¬,�Fh�RJ�X��E��=M(��,�RP�K�� ��K&:�-?�����p���A��tf� )�̑G�����;/���[ˏȔ(Z<��А��q,K#*�� \:��"wZӲwү&��]Ux�3Ժ�k����}��M���:�Ȼ�!`�O�����;:#�ҙ�f���S�4�5����t !�!�E��c���E�E�R;�U-�4���Vr "��IzM�g�ĿEtؘ��	ޏ�/��~G�ßEj9����cen�-5��UI>l=N��SS��Z�n48�7^NR2�箭�R@u�/,���!��J����h�}{��:W�qih�V�L�;B�A4�T�
ںN�q��E��D��q(�f�E\��w�P��k*&B�~(�6GJT>�77�h&:�����0*���nG�-�kH�r�O�#^C{��^��䖙�1 ��_�EF�>�)Ш\lsu�������_|���]���'�/�&*�� �k3�j��'N�.��`�Fn��޲�ݷku~��܃K���@J�3v[]�CL�����n��+����,����σ⥜�s�?6��c .i�@�F����y6B!%�k�F���X[�R�� ה��!��m��=Py�Bߓ�k=Mf^DM>Gq��"�;h(�b��0��Q�V�)��J�S�	�-u%�|9UƸ��F)Q��gKK�@W�S����d���y��ME�/��j��BB2�7!��߅�S+��#�ky�\�T_\�%ö�L�nzYpwE�%T�0QUCf��UygyWL�w�e�FP^��Z��_���Ĳ���`�H}:�/�vuETкf`	�����W�j)��C��a�_gӢ�%�52BO�\�ݶg�WN�����?�4v8�bӧ�Ol���U�������聟��¼Z�WPf9{�Җ�����!Glq�F��B,i����KkUq���[XcG8��w<�h �H��Xwe��LE��ٿ@��8�Ԡ��J�-_�/����,f,� )�K��8"�tR��W�0�8(Rw������Mm��u޾Gz�ZlPX����Y���f*(w����X�AJժ�cI{�j#P(���:�����Y�Ǔ�I?"l/���<��_<~��h�/-��Jջ��&gsI��E�Be���W�B{L��ҳ=
�,�ED�"L8+�� 2�z��F9��$�A2���������aeE:�%2! ؎#����n��K��V�%ޒ�k����jl
u���/\�x��Zz-�f�F���!��G��޷�N�!�))��@h��!�.�l�*i����)9KdZ�W�i�ɯ�I�U��~����4���}�Űh��zg����ؠӔ��N��u&�L)���E���綉	.���ߛJ'#��j_�El�-��*X��x0E�*[�R��CJcR卂��������ʎ��S�/�۱�q~>���`�Z��IH-�&����Ş$t�2a�o�H^Y���l���dCaJ�ԓ�e'�h�֔>QBSֈ4�0>����9qsדC����Ԛn.�(⎪H����[������NYxu�|��#��^����{?X
�(��fLV0��+ip=��<��pR�E^ ��>��y�}T�0���j=�D�݇�u����S�I��ޑ���������m8�⮷Xy�F>ڲ(n���z���J�{0�-p�.gn�0����A�0�����Awq��Yt	�����~\��?���sL�0�r���wZN���ށbN�����'��}�!&VO��0�|��Y�b�Ř�u�m6�
�Di�*vx1�6�HD��.;v���a�i�̶�Pd�T@X�lэL���f�P������VΔ����>�(�y5��Ǡ�7�e��P<��-sn�O0A�������,ݲ�����_�s
��g��I�a.Њe�d���19�W��w����̽�5VB���2��e���J��a80��v�m��^��~�nMoݼ Ee��1��B� ��l�ִ̞�)�K�0*6���|�)�Z�t���r�{-�9��6� (���L����L�%�Z��m�U��JU�r�d��!A<lc��^��u������A���K ջ.�kUT���d�S7�
7����c�u>�ơ�(�/=��Ҋ�Iyk�c��kl6�|���&�b���#�������=�k�v�cƉ&��S>�/�A�R�qh�D�Z7\|a`٧�];�}���(��F�ܵ��'!]^69
��b�$D$˄�0��f��qb�T$f��Jg���pY�N������4sf�-�f%ݡ�W���)�����a�'W�B]�O�'�8�uU�'�F���>��ø���QCy���bu��O�O�@G���ؙA[��"�[~�� ��B����S��u&��7�4�n
��Qʎ'���no~����aM��r��u�E��+�K;Q��(�\��R���۹��YL�>�^q����K��?����������σZ�J������|�uQ��Cݡ��s���!KW�G�-�vU0Ju���]T����2��!#�}���0-�|Zh�3�u��d�1\��=�� �xk�	��VQ;� Y�l:E���vȇ!=`������,V�z���H�����W(j���hD��+874�y����܏M���N��vJ���)E��_�D�Z��S{[бT��*tP�o9{��y����E��0T�{��
X��~J{�2�<~n9fUb7�O2��u�¡��ɭ��H5�3<�5.�^��VDR*"U��wQ�4�8��Q�z;b�ϧ�Q���zp@��dA�G�k'���lĶ�3%��2�ݞڔk��W[^�㌾X�0�&�e�w���7��(���W�<���u������Ah;OPŞ� ة�^:�#�-�5��(5&^�bow���Y1���s�݅z��������U��,��r�޴x��M�4�1�GX�x�МǴ��:�����	D����qQ�ѹ�ߌ�@ir��b�Dӎ4��yl#�ϕ��~�Z#��&:>�q�rxM�s���:���ŵ��Ge���w���� p|vu�/f:%FK&r�j�Ҧ������d5x(�R5��&�ul=�Й���!���h<�&`ύ�}ab�XV*徵�=q��"��C"*�7����}X�`�#Qvi�O3��'qnw����kѧ��o�>L�"��o��:�Ճp\��#j'0�Ǿ>�F��95I�������2�\S��71���\8��q��^�o;�Ū���3O�/�M8��ޙ3��!����Ooz��a��U)W�-v�	�[�Brd�T):���ؐ��h.q ,.�9\H�L�����k��+�V+�B�q����?��n�hﾰQQ�]����Vw�gj=" N�a ��1�݉��j�>�o���#Q��5�����U@4��pM0Z��V��k����r���$y)kM<R�[	��(4�!(����~쁤�Cx�����i�a�&��>Nv�Y�lưM��k���G����+�%�:�r"���i3oc��Teb�#�O_4Z��4��Z�����޼mx�)_�r����w^��N��u�9w���zB�~�lJ�X9�B�g,)�1&�Mk��E*u�iG���H5�K0��\a�?��sL�bP��0 k�/���(����2ŭ�mv�9����\��R����JՀg_�w� �9��~�������.�jF��,P0��eGH�gc)��z]��U���1Iи�m825Ȏ�A���8-�V��Q���L��0�	Y�����(����*�|rfa�!@��[��\�`�������
7x�;�2Ag��Q|A��{�N�h���[�k�yn����S��Ӗ����5���zR��f_�{�E�?u9��:<�-,����D<���A��ku��[H��N�_��2c��Aϸ5��f��>`�/	�j��$�2��ګ�h���׾+_)�ܠ�0�3����l���T`[�@�`�#qm9�>�<A�ySL������?��tK�b�"���Y���H�y̥�4\wFƆ����|bAF��yJ��s�%H�- �k�S8�,.q��f�kR�z�U�C[Ǫ���}�����q+�q<�>Cj�F�Ox�:
�Q\*�sO�?A��Q��]���C?���ųa�\-
��B�T�t�x׃��h��j&DRޚ��V�q���+��q�_."�U܁�-�3CX`�6���֦�=�p9L��v4�y�~�m���a�Si�X�]7�Y Ӻ�$G�����SY�A��}�F�~X�ܘ�3Fh��R;�3���F�E݊ڹQ\+��� ��eF��f�O�~�_>�&���ͯbg�x~�.���\~37�*
ˤj<�J��o�[���d
9Y�T�YU�L�"�@�UAs�ey��2A�ы2E�7���'���s�(�+��C$��8��B�z���ͳǥ��G&|�ף��L01�}k�;?f�q�F���W�$vzF"���;S��+�t�}�����$����&e�,j!q��2D;KW|��k $&Cy��i��~|�]T�������~���o��A�XF��(}Q{V�:&�ud�ńn_W�� z�h@�(�`S]�~N��(*�?f0#%�+r��G���}):*�Ù��0�a`��ё�F�*������l*��� �}�Y�5����|�\c�4*�>+�
|�����
�_�ޟ����,������(��ʲw��?���,-��_���Ë�FPy~hp�_f�i�â}�
�Ez<�5��*�RA����LzX����"�=ݽ�ZK��>���NU�+�����1���E�{�QV�p����|�c���)�!ն^�|k���k����	�$6w���/�#��SF'K1��<ad���h���Vg3Ŵ���V��Ml����;2�(zY#$Rޜ#��7�\G��B��Z��A/d,����`g����3��EKRB�����(0�_P.��@��'�k��ӂ�ޱ�gy��O��o�A���bG$���e!��������h��������3�cO����C�ڹ��zo��'`+�����!c����n.He ��x,檉*_ ��!��Ԃ%�;[q2��r6Ӵ�fS�g���o�ɥ�~���Mx�B��ft�K��>�3z:�Hʬ���;9;w�$��V"K����ߋ$zQ��>�/��9� J���v|b��F"D��BF���d�I�8"Hz�g�O��n�&�� 𾕂��wFB��?���Iɍ��Ђ"- �{V�Q�^�ǚ<����s��ZiR�6�E�L�&�_3\: ɂ��!�����2�+ �����Z���h'-�j	�|��K ��~���fG�ᰄ`V�4޲�[����.C��|��7z�� ��u+��l^н�3����݁W?&Q,C(����]�y7�J�D:#�T��U����CQEr��$�Ei���m?�5��J!w9p�lڗ��sj�e�⟊ ��I��%��Ը���h%�fQ!x�����BV�`y��Oq����fT����"8�tIZ},ʐ�����\n�'U(Ω3����������Ѥڨ@Aa~f������Ly�<������hR$G���,k�d��O7�ذC9SF��;�ﱟ�=1�F��@d�?�C�٦��mX�r�HrJ��M�H��ZJ��1�J/�����|^)�#��d�DX��w���ӊ/<��9ݔ�7 
`m��K�+�u�W�v��-D��u�щ���㯋3�I}�	���K���5��J8��c�0<��J��䢤�P�E;Cz����|���td�C
�s��4K��Ģ��+���d����eGC��:i��,�Ǣ>�����O�������[��`�أ�wg�N7-,,3X�8I�����M٦��r1-��b����6x��8�;E.�ַ'9]��<cŶ�9�{�jt8��Rh�g9�Ά��KC[?M��p?#���DH��|	�z���M1�:�N�bnU�BXv:��uKtsb �N�k*�S�	X)��B�P�=�"Zr�|���"C�)� ��f\f��c��{^X9F	�>2w���$Fzʏc��ۺ�b�P�ly�f�R͸��zV���I��/\`�ń�X(�d=)�or��l���7�+i��Cg6:Z;X<�'�2o�a4V�~�6��@���F?l"s-�sf0�O5sui²�/`������u��X�V~鰸���R�Q`�1r�g�a򝣔�����xt�.!'F;":����SCě��0�PMI�Î`�(��u5x�Z����[J��}Ȱ1v~�Bf�c\I�L5�wtLh�����p�mܫB�nr��1���vv�0�CK67�P@�Ѓ��XI�S��Q��ؔ�'�Ŋ��RЧ>e���� Ϯ��	,�,fJNKoKD���F�@p4f%�f�>�"
9�F�X�z�$���Z��q0m���I.>��)��]�mD����3�Un�߶B
ˮ
��mIc�UV9s_��.K�G׆:�0��uǶ���}��fd�.�1����w�0F6���ܨ������	y�ݜ�5�(�-� �;��p�ĶdfH���ЗE��c��Hc y�ZľH�A���1����5�A�O��h���v����H�4�$��O]�l~#�6�@Z,��฀��a���Z��8��'zv�IǬ�z�53���3��78v��O��n�j�A�V�]P�Soy�2���p��K�n���&�ov��C���bΉ��W�	�,�r\��@���t����\zw��r!j}��"���{ZLŔ�qo�A��uqQi����w�pI�GYYۑ�z���Y*�u_s=Nq!�'�Pt�-`$�!�=0�uav��!�ɍ(�9U�y���4�b�)z!�b�=�h�\3�z�Ӹc0��_�l�a��%��Vn� e'���+@0��,��N��dFy��l��յv�����Y�m���5�O�d9+i��\��b�4J�V���fr�Dk>��ětpq_���7W��� M�z���_�E�ÙPn&��9.�`G���ʚ��8`��)3.D�1����n!U� �[�JD�v����^9M#��6Fo�;���%�|w�Y��}`CS|�VJ�j*Ŋ��ly�b�[�{�Pp�[�Dl�=H��][:���]9������$�yP|�L=b��X��`��o���A ���B�>wr�:@xJ�)�BH}��$>[�9݃��W��w��q>ͧ2���NY�r6���
?X���/���^����*��6B��>���*>{p3�:��Yɗ":�x�:H�L��ַ�I5U��#���˯�eIs%��a/���wB�n/]"����Ȑ�����X�ZU=ݩk��@8�_��{��_^9Kg�y7='�hQ����KW C[
8#9�7��l�'s��b��C�c�i]�%��\C;--nAr�Z9*`��H��ʒ�
4���Wp��ߏ2�:?�+�ʄ-Kwp��zqzw��y���K@]P-j-'R�7����7ƵҐ����l\< u�a.HG��^�)��	{��/�����f�����HF��<3ў�Д�Z��\##+��Wj�����"�ꆋ�a����X*��M�c�h������X�}�3�i�y�k�%�a1��Q�f�?� �Ǌ�����%����f&�ä�G����˖��v<x�Mȇ}<D��&Й�*��,a#L���s-���ˑ|�}ޗд�_�:6!����|-�B�h�TD�b��Dڏ�S6Zhm�ee��F���)�C����z�q���ҡG08o�L�2Rm>t8���l�w��̃=h	��'��Gv �~�8��|�[(��n���4��2�a���)�m��(��E��A�=r��4=����R������iS�s�[�/,�~�=�#���*�NE65��-�S�W��p��~��>���t�=�N$l�Q���R�)W����N����6�哕 ?�wk����{ZH��s�-�о�@��t�#�=���@I��f�/@p?�g���Q���<�!����B߃ވX��Z]�B;������A���(�k}�Ռ��	iդ�<
����#�f�"��X"��$C���#������p8t��=�y34G�������ċ����s�+���Q��ڙO�<|��� |�d�S�#�<D�Ӓ~M �bk�1C[�ije��S���LT��Z�(�O�?�eJ0u!y�u*���I�l��� c�[O[�>sK\���2�|��3�����^=}�W@D�}%��J��:.Jv`9���4Vv��ھ��ɗ
�Ӻ�b?��S�v-6��맛����!CnL=Jd��E�`ekKӦ��cBiVF�~]��t���xF�G�B�XW�F+�uxȇ ��MAn��1����(��>�ܻ�B:�z�}X��ח0/�V�g5��P٠�V�������lv�}���@-����
6�Oknv�U�O��	E�tM'v�``�Z\d���V䱎���/��(�zN�[� 3:��زQ�Ly-Wg�'��~���;_p|~тڙ�^�Ÿ�����D�F��"	�� �02��)����#.BɣR��5�Wg[��=�긹�~��J2��X��`r�'���'��%|����duc�Q�>�H$�GA����Λ,l��a�;]GL�~?�Ge�G�QT��
g��T�Vz{�ͤ��6�%�X��P,59Y+|��.��3d*CI�pS�O��Bׄ=�Uq��9B��j�z%�m^��=�b!��i��=���0ZC޲��ko�4'
�4��z{9���������7;4a+�Ř�����$$�;����#w�������A��.�[�8����5���}?q�����qu���V�����"�M����<v���i/^|)/�pS��)c �7�l���$Y�:l�%ރ�Y������ه�&#������'��"Y*6ߐ���1Tg��h���B�_Ԙ��rh����!^͏�O�x�:a�;����G��+r�3�Y�銘Ne:��b�:&V0������2g�j���$W',c���6���ȣ����eL��;���7�pG���o�*��n#�8�ne�������ϸ�����oKM �vf�C}�Ke6���|�U�Eh1e�6��w����q��=�Mu�}�߂�T�j䏭5�h��mc��X�s���{��\)Ň�	f.�i�S�� �32�����
{��*�7)я}y�6-������I���+��j��λ������w�4�<�k{�5�@,ݸT��>�{�:0{^'��O�7�F�s�:��������7��8����qK�+�F����q�K�?��<��ls�$U/6G)~SW��l�x���>�wD����ন(��
wgk�n�K����]8_�����Z��K>����+0�e���*����s��� X�C<�t��L����"o�B�n��b�I���/q��,� ������d����������J2�ы��t��g��x��L=y �8$���|�a�4 �A��˥���V��nt��3�>/;���x��U$E�H��C㠒y�j�v1�HUA����蒷����;����am�C�'aR��9�jL��:=�t�V�O��Y��<-$&:vf�wA�
�D
�%���a��}ˬܑ�B�Czr�b/��>7�ko�/��-����v�}�.h���?�[Gҳ�\
S���%�Б�9�t	[6#A���F%ό�.�|�:��uDΪ�	��_�1l�j�HL6G_���������~����.��OZ� ��h:�y�{�5�� �o?%��I��*,�����X3����B��Ҫ�p�&a<�;]�g0%��|ztD��JP�$����|�Xi4��	$����H�/�nDd��cz<�:	$+��*Q�ZA�0��h���A��+��lN�5q��e��g��n��"pY��8fG��I*�Ku7o��/����z!�B�=��VeW��m����ͮ�4�d?�l��W,r|X:���?�q4z����K��8�XIhr��ф`��Au�w� 7��K�	����2��7����_��a�7��h��������m^/{�sI*���<����jf1`�K6���0�{��±W��1�E��{�V�|z��w�WJS�$�s�T�!Ɛ䀋�e��$Y^7&ޔL�K���PGH��U,Dw����پ�� �����awn�G��'�+�q�0G��%K=1�Z1�WAf�-�.s���SZy��X3�rv�j�P�?M�/�I���=w��u	��?���7x���Y=^���T��7c�h�X{L �{��X|���2=��ّ�n�Ь���﹮��9a��2��?��HT��R�����B
᭭h@�n�O�˓�|0�����Q ��t_P�[�3l������G�T	N��,�Nt�@�u��@��<,18�Pw�IB���7� ��H��ZΛ��i6���|����z5��	�@�h9I��5�@`?駪�Bw�֠@6ZhcIg+fo�u���<c׺�CA�o�yԘn�oC&�w��ǈ��Nn,�ps�4/W��/j��]��B�(B��"�nƟY�.��;��K��y{Bu-�'~��."���F�[ ����[Ux�d�P@}s�,?��X°��Y/�/��0��y,�e�����V:�	��u���}m�50 }X�����4���ͮt�����n����g���������'��xOx���Q/]s�V�jм[k��U�;�b�'ZD�y�ŴF���~̐E-���B���ő.�m�Q��QØ�u;�5�u������L�9�7��~��F���0�ݖ�]n��3���)d��|��Y����$��g�/:��H��ID8_���&�hfe��'�EV�7|�
5�+>�[�ȹ�&�~8P��
1�Ƿ��<�Ir�u�EX� �M��蹤�;p�HN�gX�W4R��	�Ww�o����SA:��%�M�_p�}������.�?1�As���M�g7-)���&��Wmߞ��0P��!�կ'C>rBn��<�@�_��j�O�!z��W$�&���$`�|�x�ǳ$HT�xx0��3�1ۓ��<��y���N$�ψ��,����,�Ls�6��Bp�>E�޿>��Ȝ���	=���9__�̫�����'��~$�8#���P�k�<k!�vy��+t��a��Br�QgY���w���i_��a.��n���K�+�Bc�*���1��J���_A�%����˹�3���t��Y�N�㼭�B���v�J֟��5�G���s% ?��"ݠmD���g���ƕ��@�5�z	�>F>�������tUU���H@��%��/��#(I��/q�^��O�Sv�s�/)�`V5�$Y��=k�������l�#��+�UJ+Q&�A�������5����є�?���Ćʦ3@�J������`x�j]x��ې��(֖�,�p,"�|�&����̴�F���ͨ�q��w�X�z%uC�n�2
�$�56�*�C��n�����1�u䙑�����Ϊ������vg����Vj�g]FW����R�^ٳ�$�bW�fu$<w�囖ЦT$��?8�C�r�زF`�8$z�h���xH4\�R���}Wku�g�W3��Lv��{&9;�����e��K��A�QT���P<*�s3��$�V�UU��������7&��'d'd�L7:�*F�:�S��mڻ�O�hyges��`ٲg��&`��r_k� o&g\���%F	NH�5�FP�Lv3w�#1��B���6$:�����Cļ~����9
�2ԋ{�L�.�Dp~e��}ǥ�m\2'u��}��u������Z`B㇄s���Y��|��3���gi��b�y���f��I���L��H��q��3C������9n��#�! �L`΋`��4�C�d�o��w�3��UΚ�ݮڒ�c늝�P���5"h�43�m��uvҽ�0W�1�bTd��3�I������8ҵ����JS^�U(+֝�iF����ַ�`�+���6-s�'S�a]8Ֆzl����s��5M@���� h�ă�T�<����ݑ?�}x^���ҹ�c��g廁�Ζ��}�"�o��O����'��P����R ���F�����ҵ�bd45��X�� ����Xg2����t�X�_��)rjj�����H~(�h�S�bQBKh��o��$<!�����`$�=o��-��F����`��}��3���_aBo����k�dcĘb�Z�wm���Oq��;{$gz�&B��N�${C��4�[���4x�-����Wa��p�l6�[X^�� ��7I"����U�c�;���]�Ѕ/���U�׆=
��ݢ�l�$�+/cj���T7W�;�<���b^�,�F:U�XOj�:����Ѓ<��/mq�&墠p{�_���W��2y%`�^Uʘ���5N�����6y��&�;0���񵳨{8�sA�߯j�kS=�s�A}�H�PYw���*"ݴQt�8�����M#H
�U�tAF���$;~����+0
�� ��$E��0�9�ow�V��¶PVZ.���V����!�(�%&$��Z[��*fE#o�ʇ%=c��l~~�e�~�����}�3�Ǟ�w"��*A7ش��v�M��:�E�1����B/:��ܑ���`e�ڗ��"J}�#V'[�nl����ʬ��ԕt�Z��Xv�+�O�=�	�B��>���[�[�q�l/tni�������7X�0��g3���uB}�ބ_�v\}� �Q#cL���L��j޸�#���u��{��z-"Yo��>`�T[��k(z-/�����;D�iX�-��4�1�kX>�)3ÅD�M>�Wd���ԑ]���r?��ּ�������b�S�
�xry��_>�B�4� ���� ��^� ���x�]���4F&	Jh?��8�,�y��W"�����Y��߁u��u���'|QВ�F�5L���],W9�ޢx7NHf��L;�һ�������˼ �:���1@"8�`�Za�)D�����xʍ6Y���BJ�r�-sjB�7���]��l��J���R�^���˞ֵ:N�`�����|��T>
�d�R8������[��������{3?��qy]���k1OD�~�ﯓ6c��La���^� �]��x�_3���Fq��7�ȕ��(�GAc�DD���6�)Uƚ�A�F"��Y���~�#MLt^^�y��Q�땊|!`�5`�����ɞo��#��O��m�
�%�	g�,R�����`q�t<�t�x�fS�0��r����מz�(���uCh�0��8��2��'�g�)�aZ 	��6�7��=�`���Q�u��<g��P������B �E�1��v��G��:Y�T������,�\b
\��Vw�B������G��53Hd��D�P]��P�j_�o
R
��(�������8
H���%"N�>@$q[]+�A^6���E�"E��sCʑn����4Y�����k*9I6�g��iO��*BJ�K�� ��`h�Ͳp��{����@;83��"hѥG���%�>ƛ�_;Mrs���������d�Z"N�O�V7���{6��OM"�N�m8���U\�Ty��v�6U�,�R^��,`b�)?����H'���LwGsA������ٷ���$>�)�5��P[�bŕ{�O�U��q`�ӓ��TC6�h��ۉ�d�v�BҔK�b�R�����	>�zF\��Pv�����J����=1D}��P�g��Z1�����)��^���h������P��L
�%̺���]�g�e����!��.W�����*Aڸ }�Y4��CQ�^��O2$�uY�R2�x�ɥ��F�$��P5n����z:��i
-����1fg[�	���������g��Z�HI#`��[�Hzxqͪ�ق4
����
P�G��ˏ�8C�F_�hF�?昸�+|���W�^�q�1�\�^���W|3��P��Wi�pHCz��lJ��(Ԥ��o�2�>[�#Kc����;>/�A2��W=A��9H����%z/gb@"4f(�T}�lH]ig��tpJD�:Z�rc��!9Z$T����^��'��L^�e#%���O.�^�|h��6�����TF�I�I�Q�m�CV�7i({��i��������{5M�R�`S[��|���QϏw�Z�]T.�f��}����F`��<Z�*+�9��F�ó�:�~&+�Ozp� �,7�%�<ϻp���"�4�f0��[)o�	9��*��Q�ݫ���$cw�fF��n���a��<j����X��&ή�1�ET2$m/$��(\L�k�T�uЃ���e�>��T��{��Z5��Zz����5�E���cY�ݹ؆�������3?v '��&xv�,�q�A��Õ�gZ������c8�=0��^ם��ϴ�k8l�Ptz�`e��ɛ!?�@�6_�6q�l���Q�=hs40|�.V�a��΅��K�u��r�gy�2�8�}���-��~�����D �S��|�#����>)@��:�U^��nti�FH�~۸	��������^.�e�0ϭ@��D����+\[и�ypj�4f~�ygh�9D�7�~aa^�^��"��zI�1Ba�"i��X�y������Ƕ�
q��
2r��8L�Պ=��+�t��$��Xb�a�?!֥�^5�Y��^�����KG�)3��l�0�7}��9c���,�Z�GuU�l�{\���Ƈø�����R*�"�_��ς(K!�e�/�n~^U�9�'��?v�.q�J�A��9�&�4�v*��������I��!E0��|�w�qL6��7�gm�Lсk{�Z�oN���/�W���͢��w=<�q����q���&^�s���4r�s`�w%����p�%'�ш���>Q�ƈIQƘ�v�W�)���%���{�#��ʬ�|7���$l��1���mc�]��r��QTSZ� E�*�Ѳ�sLG{�p+�.�sd5������ �F�@4�-�rcg����dS��x��<��`V�(��$J��j"G�����_�3fjѨg������J���j�	~Kj���h0�i�ƴ[���0]�>� �q�R�'E���r��_���3�e�^�, {	�RY?G�k��L�*E�I�˵���/�S͆�̕���>X���+�aZ��w��@�s��@�(�z�c]]��b�S>b��/
�$i&���Ve�z=��(�a��+Y�ʀ�F���b��s9������4�hVM�t�p�^Vn0��Q8��h7�D��!���,N^��=�q�[U��=$��$�kK
��_CAA^�B+���0Ib�v��}ԁgY�Y�&��"9�M������WO�O������l��	\$�1ᢌ�qt�g��+mQ�70�/�P�d踙��AVQB����#\Ҏ��-_tܸ�R.�dV�g�%��K�#�t���u
��zz�d�lѭ���[�8��}��g��������bR�i���)��(ʏn�>��t�0�C��A��F�7��F�2�ƍ&ИF�2}㑑���FB2/�^��,QI�3�zʼt�.���H�_z��ώ�<��)��n�,4A%�r",�%����]6ӡ!ҟ�F������? �h�.-��w��3m���.���7Z5��o�.`'�1��U�2�xm𳃯�8�g�:�>���7���Tɼ��2����fA�,�nc��@��E��)��%q�{��Z�����lR �tR9?{�V��Xt���v�92>����.�����&,a����¼��5�ϼՖ�ʓ��MyD�|���y�`��+�ͫ�T򞓉�.��c��dZPҐ����x�O?g(B�Bgk���i�а��6T�-�9�����O�
��c�jߛ.n��J�P&=��u.�'�\3��Q�C-�ֿ��qE�+�;k�!H�D<)(%�l,�)������ .���vq� ���X��l�x0>����^#�1r���8�!&×����%�O�8Wpܯ��'������QB�?��3�w4��<�0�Y��(i�y����U���
낒qr������ϲٲ��C`<F����<k\_�Ł%�+߃r��l��C6:hM'�Q�\8�5�Dd8�ـ��:����nf�����u�ݍE�g��Όs��n5����0L<@o�ݹ�{��	aYW)�kސ�/Ȝ�n&�˃�=�y���1�0�[էXС����p�"e��O����x��@�sQ!�$�@����0���m�.��;�Ӷ�?nH�Dɢ3�kuY�45�������&��l��`��Ѐce��fp����\5(k)�H,����{UE^�^a.eF�R���?�g�s�~LְN��F1��v;�*K���(�C落<��1/7���?�
B��i|�uf�wx;9�ub4�ПҒ�f�`'�l����Y����(e����.��2��e;�_�fh���ց������7mN��u"����5�{����-X��x��l�6��D�W��R9��l�hh�KY�N�Dx�x�<��zb�]�+���k(�GPd���Cv�H=��hT�x��Ed�H�m@+�	a|�=������ή_�,#	�����DO�mK��Uè؊$�6bٻ���^�uo��r[�(.Jx���Q�wOĕi�:Hp�2S��/i	Dg�0U0���m�4݀���(7�T>%�4l<�V���=������wb��	F�bS��<��x<UDn(*��9�s��'(i=��
Z{x�z��g�[	0$03}���= �q ՇcU������g�3A�D���K�ԝ��o�u`����?���R���Ӂ�����Q���0U�:�|�7�����woȫ��ā"�v��m��\�\�[%UL�t��@�M~�Gf+z���.��V�:�����wKg5�W�؇q�8$�أ�7��M�����7�&�Ǳ���br���.{x4'T�O�n����_�p(�����᷊������	��wE/Ho��:��� _�]����Z絤5��tb� �u�ՅX�8�X#��\���lq��o=KD?ҟ�n�7nzZ<1~R� ��[�����T����M��ɖ#���B�j���p7�k��E���H������r���������z/#����V��s�__}���]z��ဠ
���=z��\��Z��R>*�&7�a
��'��&|�E$ᩫ@W@�f�.EM=�t��K�:�S+3y���=L��Π:�����_�<Dò�H��B99qxf위nN� �JJ^(�s���wg��b�`� ^� H\��"���Y72��;�`��i�7�oD��5E4�^��OR��;f�GF�'e�7��)�vne�gˢ��Z� �;���6b$�>�xq��M/��h�f�=�H�WD&)��鈪 ��v	]J���	�#)�P��S��_��/'�熽%,�^��R�G�8�,�wo�_�K=�0�M=}����g��O{�L��� .s�-�pt�p����+��*Lg�}\s�6�����	?��ea��;5x�Ev��7�I���m�)v�����4&��[q]`�@�	2��r����	8U�Γ�>���y�W2IRs��$)D�՛CiG�s*�i���p�̲:VZ���ኞ�4z��`\��oDHUp��'҄/����p�n�$�/ѝ�L��%xI�L�{�W�l0��h�&�9�V��*ֺ�<Ce�����(�Y;HS�ב8��&E!R���昫(4?)*��8����cI�5�.;/z-=�!ħLb^c��f�C�z��8���}��7���؉���abˊ���?�����}9�]��<i���l��o���f�c�-���6Lr���+�{g;8J�-%���\n���=���� �0y�&#��Q�eh0y2.�b`�y�B�n �M�\���z��z���S�l��P��i��(��z�L�W/n�WL7�<R�-�l�xj��u����C����x@�f ÿT����� Fm�r̟^�wT0s�F��B��m�����<�uI#{$�A��H�E5���T{��Z�6�e8!bJAb��F۹��(0>ҭ�W���F��[2�����+K[xi�3�U�4�)>��H��q��֗!�@�5�;*u��|�Q��sD]oTL�szf�$;�� 3Wj낱��vV&���2���LgV��k����p쌠'��#x�e���v�,��o~�NT�����''��%�_��ט���H����W`�1iy;%��Rx5C���j�0��$G���Ѯx��X�m�������ig��, pL�O/
��tGx�C0�"��\3A�4��̾�ה�S�ԫl��lɹ�O�������"%��ƴo'>���!sֿ�3B�5�h�(&��ؐ�"�ўS��Rc��*x�lc�ƎCJ�1ʜx_�O/`*��g[̡yɴ"�r���m9>��{X�N���w�~�u�����y<k_V���M���@��wZ�On�zK?u���OH6���!���.�Q��$ǫ�%Z�wK��2�����Jk�6�S ���D�A���6����
�|xYN^�A�C��n��lz	p�R|�%9��O:�㔬�䛃d�K�ZQ���a�]�t�`F��*�GS�b��9�zW�EUMK���U�����ʮϖ����]Z���ة�M��ݐ�"�{�G��?�fsb� b��$<��-^���p�B���합oɔs�Ô��l�������ːͽ�}���[[��Z��� �r��g/]��>�mwckZ��>��ЖG�Ŏu�mZ�Ժ�
�\�	|;$��-�/ dD���v�߳��[B�{�0)o��̊�Gt��<��#�9�� 6�+�VΑ6K��uym����R�Y�IN��D����A�W��~��1���C�W��-YN*�E7����_.IоUn��iĦ�qg2g����@	�z�W{��B�첫H��C2T$
�"D3C�����m�cV*Hh�A՛N���3GJ�I��05�'́h��m	���i�U>�HD�Q�D������Pbe�JU�=���>]'��C�d�m�_V�����}�->F]l.Jj$5�PyP�{��V�Ǡ[�8砦���� &�7.�	f�Q�nN�3!(vF���I���Et+�m�k�}u���<!��R�m�f�5%�G�[��i���c����8VN�����/�����ʒ��m-�KX`3""���e��L	�2D�<�HO���Ō�g�°#Prַ����?"�J���k�̍�ϑ�|�$���;S_
\���I�zT��̮�5����:=u�S뙀0�U�z�su!S�:�8��>p*i���Ja���vA��nSeK��"]�i�?��]��à�7�ނ���81��-4�����r쫳�����PF*β��3�I�)��ږA�&LѓJz���)ÛT$�Ru��v5G����7P��rۍI����]��u���4�yi::�o6V����S�S/j�X�V��0����W��\�q�ji�u+>(�T�[3뉒�G�l5a���vZ���Q�>>����_��h	�"yf�$�h0/F� �ٕ�M�v-�1��Vns�e!:h�&���%�bW4ĕ�i�p�t?)�)�cߙ�bLh���w��ڡ4�JTx���}��$��D��+>3����Fy�>�����r%����Ij�z�2	�/z][�|�(�q�2��	A q�a1�FO����$�\LOPS��6������{��w��=7rk�Q��$02 ��j%#@OjaL"�~{�$���3ȶ�i��+���=����f����q���څ;!�Y3@2%�C��ǎ`-�}���gW��W�Ba��=6٦&����yg��Ldt��%��e�&]ۨ0>L��c��L�o��bC=&&OvG�u��WL���i;��T�^��B>(��9�R�t�ϦZ�:w��i&]�X�B���[mV��/��8cb)���-����sI60)rڳb�SAj;	�݇�ʟjAY�6�J�V��A��5{�N(>'���0����M�H�&�����kă�hr���h��O �)��p,�W
`!͝N���?�=�R#pó���M�>��إ�� p�j����!��>W��w�G�����ЍQ�N_�G��xHXQŁ�;3.�O�,o�*.$k����b?
T��T�#8V��	4#R&�.�)��(*�Nu���;iqq(
�#��r|!^����m]#�y����&����Ӽ���Y:#�5��K�E��bU��_����t�u�,qZ�,8�X�V���V�8�ʦ;!��҃��&�bW��4`	n{����1��s��s.��=2�{��y��#���T��ܶi�ܿT��-wK��ݝ���s\��
���ئ�GiN�(����BD�����Yȓ׺�.d���R��gL�AG��e�ʔFu�����6�D�{�t�l����h�O`��H����h��{��'�������=Y��E��:��|~�mRs�PG�T�
���LpLJ��u�v��L%8�"��j3��1�����|{�0m`@�����B�@���A.x���O�g�;��N�c+PJ9�b7�V�Zr��E�g��:�i��#^b{B�UQsu��h2E1�(*��mSj��5�x	Ye�#p�ys���[�����[��K<ph��ʔ�3*,Ux�"��΁�*���<�����������d�D���0�!Ք���e���Ί����:?
<�DH�O��Ƥ�X��׾3I{���|:��.!�S�cgl�w
-�����v~�g<�G�	VĈp��%���Fe?����K@�azw�h��7�4j =���GIU�+1C{�]�F߃�͇i�'�E�jE�枕�+�%�(���C1������9�*�����4�Uѻ��x���%��C~��Hȥ8�6F+odT?|��[O@\GȎ콰$ڋ�5��Ƕ^-Τ�=���~�Š�(3C��0�s��O�q��f�3���/���fnm�*�vi�_����Su����6���0Rع��a�|QJNE_Vq1{.CZ��IL=�@q3!�,����и�}i~e��E:W��1�h��>�� T�a��N�SKu}$?��a�d���}H�/|��<��D��P���8�1���Y�mf���CҰ=��b�����:���.\� T���=��B��4���L "^�N@F��ę)���\{r?g�W�O�#���"�[&����Zg��g��'>��%9������d�>��D�:��O�98���!Ĵ��;�q��-�+�ɓf�4>�t6� �?����Q�b=T �����I��'%�dmyLh������.&D�屢�4���i#�p:⮿��ŉ�����_�*�D?D����8�I���z~�_ئ�K���M%6O6+��4�]	�L	ҍ)w���{4�����4$���j���tX]D�~(����葉VbťH7�]8�Åh��.Y�^�(����x�48dhjT���.��4s=�!�;�"f�.n#W��'Y"%n�d���@�OR�����|z ?1�VNT��������=�ٍ�9ۤE�C��S/#�2�x�܅�rs+\����|���:vY5�K���VGMvj��~��Q�i
$w �#��	�ۦOS��%Eڦ�^��j���� 5��23�O��z��9I�*'�8�f��*�E��d<�"�i��}$�il;i^�$���?O���)�6_�>���X���)�
	�=����� /�E7�,l���2�Y����D��.�'��/�i�T��Ȩ�̦�U�V�L������C��/K+�}y��q[���"�rMn,�b]$CGY�����jZ���311x�<�zt�D��b���;�����n�����V�C ir�w�ۂ�(V�b�d�Xr,�C�X�"����hG �޹!���LEO��nQ6��a�u`��������0n����ّ�Ӡ��EU�#,.�C�WK~�;Um=�[�n����yP͟��ZM�*IBO��5�(}��e��w*;�� ��v�*�2��	Y(�����+5H�Iy�p;��O�|.�֝�����c��� ���4޽Jh�@Μv��S8�|�Q����gWM��K�f���W�b1���c�Y�c�.����]ݑg�\m��>�u�[ҏq��Cܵcɾ{p�T%���Gls�. 'B�t�/vຬ?Hk������v*86�3��>�b�{L���%/�o�d������Ǌk�*���~�q�=\��*MG*���(� ��9����u��R*����ߴU��V#�5�HG�����޶��	��/�����.�O�+^�9:�[h,`�D�<���IgJ[0�?��隭�M�-v�Ot�xG�ȫ��kk��,4��4l
�B�m�2���e���ԒW��d���;vS!%$v(�#��b!"�[#=��ҲSA�y�m�#|]����k�*yG����C��NB�
1�� "wE���Y��y�u����X(�e=s��s�gZ�OBy��-/ �OS*.��R�n(�i>(bѡg��m�н��ۉ`�^U�����b]?؃b��Z��R��a��>����N����
6�ɗ�'(���4�Ŵ뉅����)��u�-?�s�?(��k���#��O6�IK:qL
�Ϙ���q���,<��0߅�o-Q�4p���}���iýI��с~�96d!�mKDEnOK��Ō8�
���Ĺz�6��6.7+���d��/�M,�f�q��帶h����I`[Z���3 1UFkߊє�j��ʯ���#���H����C(9�����L�Ȓ�{O�Sq9ʔ5n mΜ�0�s��t�p�0g�Q��(nv�Tyw�X`��[����xUb�a�ƶ "�(�^�L�ǐAuxϼ��T+XY�@�t�g�X�Я*�۾G�+�p���d|2�+����,o�>`�p\&>��9R�����I�ﵖ\�%�۷zi��3$4��8�FP��(:��§��Cl!]0I�������qP�>v+"I8��^Ծ�����O-�>:B�9D�bN3�?���,1����ڋ�{���$����VH������FE�,aU,�s1�{|x�$����m+�sƗ;���ҋ��L4!�C]':�
o�I�g@x�Т�9���e=a�3u0�t��8	�V j(�%�F:ԋqc�0��oy�ҼF���"��*!=��������M_��J/�^,
�� )
%҈1��4�*��[�'�l���` �u�,a��G7 ���Q9��B!����>y~v ���6����@+�.����� �%uŬ�c% �͋�O|���I��l��
c���J�Yѣ�.�@�0�{ �9=~�	�b��4QU�w�ݻc�.P�9�s�_d�>�>��2���2���x׆G��zw����d��q�.)fw��'���v��O���33��l�ý�`�C����R�Eq/9�[�9��������|B��2��hGWvM��r����B:G�M��U<���
C�ޮ�l�/�'L�a����9��;�r����Ro���'}{'{�FX����/M�%�4�Wb�V�+Z���jp�?�����Y��WG�K�9`�u|�>�'5V����Wj�A4�,B���нc>����ּ���ʂ̷�Iw8�[r�t!�D;��i*�S�(�0� Ee�����w�]hK<���LKX ��[0����Rw�f���8;�F�u}�6@��/�"c��f]�@0�C�2����~��GT[j7*��jqoG{�Q*B�e�'w��y)fC�;��Zł0������P��3��<��Ig���;�y�M���{� ��bY�(���Zy�u��^}���z��ԧ���~ȒK�j��!��S�l�����nlkbm-i<}c���	���vU�r}1��� O`���}q�L��{o��
7�_�{��0c���5k�r.(�j9CUi��m�t(�@�1�v,��F� �4�~�9L^^���P�$.�����6�^�n$1Q?1	����$7�،�E��Y\jkK߯�Ljç-q�jDN��hc��ͬ����W���@�}��	Pɸ?���$���H\���W��Q�������N0�7� ״��|#���.T��S�mS�����:�X�MO�>kaڀ�Ҝ���2I��% -S|z2���`����$׼H�niHvq2�)�s�l�H�\��y�r(���hE�H�"��<N���m<��.�ҏ��+�rb���% �FSx�p7/�����ڿ	!�q.K@@�޴����J���Yt���|�L�ٶ��r,
-�
0ۉ���͂�*���e��:k��hN���_��0o�����9�2.VqF���!/|�>�ۍ����gS.��DX�*ܤ�=��5�r����X�rp��f�$M��l)D�͚�$!�<¢~0�����>|���%�B)#a�m�>�q�p�ϯO�]�����G";��9��B�j�A�� ���o�Ȗ�$YG=��0��%��������7V��Z�1� �!�x=�l��}hL|�����^$Z�<U�I��`5���Y��wr�vB��W>h��ْm�ޥ\M�^ �|M��>
�FH�����CŦ��V��J��0H�w��e��<j�cO�ZP��:�P��RZ��R�0c['(���o�<U�([�M�c���
PD�E��س�j�0.8r�!��U��m}h�]�*�`}9���I% �Y.�Ip,s��@��'{�9��9_��XjUz�;��*����qd��B�G;�}S��R*�.LU�Ŏ�`�L���$�1�Z8�@g�Cy�=���o���<�yYu���2-Н��Oix}Hhf� 	�~�F'��Y���L[n����ݦ�w�#2ؔ�}��c~~!����E����n���<`�v;�u�xFv�9Ű�4>���-`r@
�Ɍ~��)�!M�_��<�Z#`;9�4"Yjs"E�!
�f]��6��j�C�¥�u
��]�IJa�d�R���˧��+���^~��c���mpA�Ft4f�D��*�Tۿ��-��\�4�G�>8P�ڽJG��Ĥ��zz����Z2a�#>U���lq�_�\�N^�+����%�#��	�
�3n��"��x2��p%?y5��&ҳ�[�=�Ɂj��7v%�+��u�n�$�����y�1ӧn�
h����"���3�Ma�5k���m��CŁ�)iGG���u���"�J�vA^䥈.��f��)���i\����ڵ���/IM�M0 �d�|�mEQEl���Ӈ�$oͶ�X�#G*j�|��K�V��փ+SA/��Uq>�ӳ�`d#�^�$1o�R�MÈ�IV��j��ae�	O�~��A	�b�� ���c(���8��R2d@�tX���F�McH\fh�$֠C��V��%	��`��Xv��	�N�X�U�a���a�T�=��6EUA�3��ţQѩ:�9GL�x�`J?�* �����Qn�x�Q	4b'~j?�Uk�p9�G��Z�E���0�����m�QO���>�_�.��N(?����Ǳ �DB�oq���쁾c�>,nt�ϔO|�v����{��K��n� dOE��pU]�O��AVf��K�؎Ɵ%d��1�v��o �tB�Z")AJ.7��?zK4�}��_�(����n8� ��0���yd�%��\u�*K�]�ٮ4BH����������"~�:H�*�1h(/�-k�S��#9ޠ�~�d���ma?p�	ه�;�	P{P��htc��&����m5�X. x�\:�r-�ɭ�\`�ΡW;1�1�
���̩͉@��L��y�Ea81%��h7�&(�qY�.�.y�s�ԝ:U������G��m(om���(���}��L���?V}hf��!���Zі�M�뛵�n��*ŏ�_�~���㏶�Rb��P�FdQ&�a���̐D�,�&D�Y ��%~n�B�z"W��lMp�В�"u0��h.ݦzx�D)��/-����Y����E��b�[�t�Ĩ;�����B{�}C�iZS��	�h�%�%O�~�B�#$=��x�W^�e>��)7|顊��b~#;Y��:�ٱ�h5Vck"�ŷ�=D�>�<�\��V{�'@�U�즑���n¬p��e���6�>���yӕ���jWS����BZȹEذ*�%����I�^��v2�#��A���?ܓu=���+��Ab����夽��>���Ƌ�ج��ixs�f�����H)sϙ����[/&��J�� ��8��FO�w��œ�a@����3�!U�U��#��b�̔3Lg��[�+���rڔ"��<̯ͧj^,��E��Aa��Efap�������6�GtahO���|��)սDX>��"��I�Lo�B�� ��rK��L�c��Nu�~�̊��I��7�F��j���T�;/�aØ=�4���\Q��V2��U"s��}�='ӮP-s~�^��Dz9�RY�H,(rk�D�hPq}�KL{\�>�͌;O�X�Q��^�s��aR4�4�?��0����~��&�\��S,Y�C��	*P��l�;���ۓ�1&�S��W��.�S�FڑC���2����e לG>��l5�b����Vj5�M�2��/a�뛒���D��2�;����%1�/JL��<z��������6oRM�bٻ�D�e�14~G\� ����2��mc�����x��tx��Ǖ'c
q�FS,@U�Ӗ�S�  �\�?(GV���y:��K#6!���!��2O.�`�hTj����h68QC��x�I�^��:�|i��a����-��k[wOP�p��<����0�8`�
T�=�J��'+�҄��_QY�k�%��vJ���=�=_3W`�)�j���}d�E�f��*9�:����o|����-���Ԕ�wC ��O�|/�R��$�������e/iW�u���{���|����&��ޗ�$�� �9���J_��!�h1��[\��p�����E�?�G�P�:3Q]��j���1�a��	���v?���I�&{��[��������	��v
������	�U��S�MnhJe�"k�W&�;2 =W������zE�I�byV��п]�ܙ<�8��� ӿ��ڃ�'�;I�4���a������ e��D^�����"}͎�Bf�Ic��	1��WOy27P��w
G��-�6����zT��1���-P	�s:9 �@g�� '�
��CB ���������b{n��d6֦6�*#�^ɍ�)�ߤ�%��V�!�����fM����<�DN�D��+���=�ݡM��SE{�XF7(Au���X.�RkҐ7���9M
,�1�W���Hv�
��贤��Wn�F�;iyp��m�2�aJ���J��(��Y�~>]ޛ�X=}KJ뛐t�]���VE⻠P��� ��ETҞ������?j��;�s�����',L����]Ԛe��H���(����3�Fc�0�R�d5�����z}qc�$����q5�;zy��!�JM�����k�� ?�~{��;��ri�lp�]�,3E��m��ɰ���z���;8c�/�ݰ|Z���f:�>	�R�v���!�H�-F4��.�����{W�]�}^su��H�ן�Y���W�V��l���V��(Y�n3=S�t=�Vf�+�cN�F! ��G�U��}EY����X|3$��Q�'���m �H��I?�I;.�6�c�>@���<���>FRʙ�Y)ܞ���>���t�$���Ct�q7���Ľ�|��1?[O���	ӄ��
�����f^5p"� D�$w"7�;���C�f���ݷ�0@wyB�W7u�g���P��i�y��f�oPUR�k���
)b�U�myl�p�K��w[�/�����3P�p��5D���e�MV��b�?�B��a` �t�D ��;��NQ��d><��58������k�@С�+��j�	�Aw
���!4D=p����d	%03�%OU-����8}ހw�u��jz.z/X��+�i^V֚�P����^�\�׹N`k*��yBW;����3B���A����Qȝ��0����F���q���̢M}[^(���8M��3�4�n�q���4n�e��'%|��A;šrWѼ�U��vO�+i��ȍ|*�/���d��Y�M���n*�@�"�.�����u"@�XB@fo�?�Q'�L��_m�dY!��x��ᕬ�٣����W��o�f�5�gA�:Ǯ~$V�`�Pؠ��*A��yݍ�&��W!��N��g8�P��Cw�b��f�ո���(���>ɕÞ�ہ�4�u?�ჽ�����˦(�蜨ّHB}U8��>�*�G3�Z�`�J�P6��[d2��	0���\i@f_UP�%�$SZ��T8I�Sy)�Ql$�;S$܆%�8�uN �A�B��X��)�!��uT-Dp����	@x��qI�I<������# ���B�5��z����e��`���M$�k��6��Dv��EM:ɾ[yp-�# �\��6��4Q�)�v��gg���'@�J�
���̵��NF(����ߕ�q�S!zO�Ox1;n*���S��M����L��M4d����a�5*���9=.�@��¡�pң�|z��ꂀp������:m��O��yv0���?,�QL�yyo��[B8��XQ�g��'g�]톂a倌����&g��ɀ��[~Ih�\�m0>�6��A *��ʍ���d�+s�P_т�o���2���h(|��: ���zo��^�ͧ_b�������&���[��	�y�8	�vE餼�5�_� �>�E��uЏ
g��`V���c5���lVǢzU�%>����@���X���gB���X�܍�w=�I`��^դ�:�<�	P�(�I6�f<�!f�W�6X�wKO��X� kƵj52Jd�v!doi#SycO�]9f��,wD{\���o�@��>�\A1[�禆H�8� �0�&�*~c�V��,٣6R�鲆�����!��zd� �_\Z�W��g�`����E:�e��3߻���~�p�/��0G!� ǀ4�BA�8�hW�9,��v��I�_���ֹ��f����R0��W'¢����9ۯ��ʰ|0׀�E�}�+,
�->��4������_0�?j�F^}+d������.3Pd�x��jŕ�m'�~(��b��eWmQfxWC`)�����@�w���/�zCvo!�;j,}k��릒���v֡�LC�+;J_
Z�H��V�ZOa��X�o�>$�����4}��mtwك�k���CL�fI��ݺN:��Ԛ�	���ЪW�{��l/L��u��<����q�6&����Z6V,������۾�ps�*ě�liI;�� �V�2z9�m�wV���p��\"{Nػ�'o�f���'�m����;����ky���`z���Wt��2��ڔ�.&���.-�(5
o.x�E����ǼwO�It�Y�ߎ��N͒	0�0�"ĥZJ�d:�%�+��TL���Au��ƻ���=����W0s�O��ϝ��xo d�FgBh3=����BИ�}YF�>��F�vZU\hF��\M���Luν�:�?Ϭ���q�m�������w�*�l ����%h��<��̲���&zJG�Qa�4W�.:s"�R���-E���G7<���/.���l��7�vP}��I���Eٯ�X
fߌp5?{�E~	M����{MB�W0�T�x6�YU`��O1^>= 3N�b���k�&ɱ#R�/ϟ��Tn��fo��L�����#e�"�|����� L$n�C�1�?��_^�p@�L�����h'��x �o��_L)M����Du���H*b�[F֟�h2�~f���t�n>�����#"���{NlV	Ĝ��x�� �N�)��n���A��k�(�޻�5	�<Z����;���cC�K�_�e�cl�@�����:���y?dy��K~epѭ0J�)�_���M�Nn���T��bNV��'��ڳl_�
dkήm^&�l��%[_r�����|�%��B|C0L�o��Ќ�<�cJY�3�ؼ�$`�kS��2�7�����2���AF0��jYKCӡ8����9J
6a��D0	��I������dB�=T5��s��+���
$)��v(��x�a�a��I>����E��v1] z�I'�D3���P�8o�1�T��/�1�S۲(2�w�ն0��<�{�%\0g�X�����q���}�g�֧)�נJ��A0���>����"X2����O���1�ⶒ"��L���+��]�r41֧b���r8��:91�����TFX���|h<Z�9�ٍ��#5 ���T�5��c.�`��}#@���b�Vv0R���x��VH�� 5]��^=AL\B�2��mY���
y�0и_P���?2�mСP�"S.(ݙ��Kz����Z7N(�1@K��"�=��Z�_D��d3~,:�y2�_�Q�,9���ՍU�����0�.K���/���u�S�)���^�O7��"Π�vkA�+w�2�o��N���Z�s~{'[�I��j|�݆��8�D�,hGn�par;h������Mc=�"����ͳ9� �BH洸���o�iL�>�w�V�0��1 �ȨDIr1�	3�!��5�0�� ~a�<�����e�h(g���5�0S}��O�9�N"�6W�	�*ۘ8�
�ө��;��4��w↭=� l�ߚܠ�=�О^�F�~�JS���}�y ���Pf��=|ͻ�"�Ir��A��+(6�u���h��a��{yw�G��C}*,`f��S��Κ�4��$�S�Ӣ0�P<u��F��ފwџ�qR�ħ��pZ�A��5��lT��4M�����T���-�h���s���ɪ�S�u
V}`��{��)2�d
�`ݗ �-��R���a���]��7֕f��Z\��#*��򀎳��:���IF�>�V ϟ~�4а�I�S���l�jt��������]�n�]yya6��!s���,�:G�੓����L�bs~9f�
H�r��C�0.��;*��E3�]�!ؔ��d�����	q1r�<�4|s��&��-7��F��c�;u�����7�D4ё�I��C��`���)d4[K D�Q��>�^|�E�����5�A���J �*���v���9��50V.K%�)��{��)�<}�Ll������L����է(�����Ik��&�z��)�HP���݇G�A'V!��VP	}c������8���Ä� �u�	%U}T�3HK�XZW���G��Q[�T��N���4D�5w �J�:SW�#��5���ZA͛f7j�����4��z۞@m�R���X�-ӗ{�$�`�>�<_	L�?�6��0���̮rg�ga�C�Yk�Dn�o�ml|� ���Q��0T-;�ُ!���i:Dh�a�5������&G����Y�G��`4�2��T�X$��v�]��s�S�b�d�I�hB�w@լ�.��=G�F���
�9��A橅�`/��9r�� v�pE�9�1�YRW���u=��g�@�FC5��"l�̦T��c��R�0m%)z��Ĉ������f=�B̒;t`�X�M����\�%(}	������)�����UMTT��uGGK��R���8��z�lx �._r�0��OX#K^w�|��{��ŭ���!�x4J��Ğ�s�����sG���v�(�W��f%A�$P	r�r���8�Q���%-��M�I�:����d�a���$E�0�"�"=s�3��Vi�����4:�ի��m9`���|kN�2���F�a� �T��L��Z��(2�5���,wg:��ka����°l8:��-ѓ�����8����}{��GiB�l!��:!�����	v�Cnɬ
\�<�`�*s@�gٸ���ƹ����׹��������"�㠣��o��c��A�cB�	＋r�D%��p|΄��A�࣬n�y��\�E��	:2��2����<��}WL�7���#2f*�\�܇P��W�0�`g�5s��}o��̐��5&�wccD8��H�7q���������	ko2�͋vJ��W&�bw�4��eQk$"|T<��	 ��U��`���1��?�����!ϔN��-bq�&ƕ�jh�҃����;�ݠ���Y�5N�[R��lw���zN�aX��I�w>φ�'�,C��3mi��FD[�r��@W�U�v��h���36��\�qm�J����.�U	�N��ڵ�T?�ÅȀ��@�zf�=�X� 6�(���h�� ����ڞ#�G �Y��%I �eLDd#,��C`�@:J�Y����}��Ծ�Ƣb�8�E���H[�_���+mO"�Z�����}�'J�w7H��Og�+~w0I���.T����tMP'����u�4aG�y� ��_:Er��T�`�����v}����Uhc�y�P<����%��������j���O
�mv���Q���D� =��O�6K`B��і"��)C�z
G�v�:�f�����t>�n� ΍�N������+/��
9�����5�٫��
���}~���ZA /Ћ�M��|9Y㫑&���%o��f�^:^`�S��t 2eh�'� ����W���ט͞`Lb�_f&?a����|z�}��y��2J���z�|5�1����7C&�( ��^;
��1���&�Il�?0�Ҩg���C|�Aܾ��nb9�Z�1?W,&���(P~��`\��g�%JL�sk�Y�,�?��@�^2,���B�"��e��|`�q�Uh�QŦ�c��v5X�������wULdU��A��#�d�E_1���QV:�>����'NIH�8�ow���
�E�r�R$�����0���}8��[�9s j`��;��X6��զ���8�פ�T8�U�iyN�]�m��*yO�s8��(�~��z�]�Q�:=p/��2�OD\6�C���i�S����^ӎVi�����l;�c&n���l��<����-� �H��q������ F��Z�h�F�2�G�1ōF�r��S)˧a��މ�ȩ���(�t膳�؎:c쥳1~��:�t�i��aHϰ�_o�v'O��`�Ն΋A0���촺��� ��}]���@
l���Ht��dLQ��	�V7O5A��Ԓ<�,��qt�=7��
>�=:�`'�t�R� �*��-<������:E:P���J�Ӟl|pW������L���o��HT�jʻ4%t�;�v��L��	�g�-� ni$u�d�V��V�o)8�ٰ��XR���h�d������#�kY�mE�
]l&�)��z@�Xku/��c"/zn+,_c��r����W��}��K�"-�xkH��px�mY�
�� F-n���N�<�y�(��2dB�歩_.�]U]�gM�B~����*K�t7.C@��/1��J�e���;S���5��3������KUP[�r%+ã�݀�� )M����#��{P/��_��y�N$�B7�M<��!�N*��~�E^�L�.��-��˩������K�C{=ޡms=9F\C0y=�%T��2zW
�A�T�*��H�מ��n�rh_Ӂ�x�$��X}KBq
y�k+�R�U�(J�wL'yF-�E�D&3���Od�����oΥ��?�ŝ�DU��	$|�s�B$k<��C���pS��k�K�~{�i�* �����T���(��] ��S��]GjLŶ��ݖi��{:玞wI^���7I$a��lLW��O2��N�qYWy��D)p��*~���r�jCE~�|q𯍇E0jNM	�ܛA�w�4
��❿�}hbM�|Q��U�a�؈�I\�ooۄG��#y��a��'��[�[g�?;_�{W�ۼ|�Ò��T,A���`�� %v���f���0K�j�L���QxvcҀ�c��C`��49���'&]D�.�,�ݱF��u������Jڸug���Z�=ݣ�>>ĉ�-�3T����,������SA��0cp̯V6wsuĸJ�G;�7��'�>���ow+D�����t��MyO
�Gx�N�]��&Rk�;0���6:�^�c�/��pU�U0/6�%�-Yk%��k݋R}�ޑ��Ƶ85a@�[ĸ��()jOv&��C~1r�\��҄��:8;��z^��{����C�b�1���U������?j�ڛ_H��ڡ�`���Ú�1U/S係ְfDF$@5���@�# ��O��H��]m���4	�Gy/�`�0d��d����k���R���H���L�!��������Z���#����n��u]����R��%)���q34
�@�v8���(H"v���-���N|�*�~ɰB��)�b�����zd�!i��jC�p��Ӄ�����3�z�^�0݉~���8�Ƽ����q-��"���ĸt:�	�V�=�)#%�|�5�q���ƌS�ᴍ��с�H��:I=�V�]'[���z���,�!��m�w�u�jy'b0o��p+ۿ��u�3p#X["L���L�?]�9�q'���~�\����}=�ω�2�[Ge�K�D�Ĳy�7����?t"pąU�p9O!��
�����
�F���ېm��n��-bo��įR�`{3��^����I{��ojh������(��Go{�3GZ�CV�|� TN_a�4�B1��ǲ����`�t�(nGz���dK���M"X��Y���1;�+H�3�8�@>��BC����f/G����]E)�z���rhO-��C�c�
��H��Ǯ���B���B�}���X��!��*\����4����Ȉtt�4�H�u�8���o- �9�[b�.��a�R�գY����1T��'�AQ��`ol�%�.�>�]j����e�ރрc��y	W�[��c�g5�Z��<�������+�x������oy`���ϷζƀQ�)1B��XYtH���ӳ}`�4k+��z���ò4���NUR=�СM���揀�F�e�	{.���u�h�G�W���|�d'�`����o�{e���v;�p�[��GҰτ10�j�&^eE%�j�^�r����ma\_B�Ȅ�����&�V�m��D
������jO)�ࣳg���Ǣ��d�
���
d������E����iN�ǐe(��0���]'��xں��~淌"�V��#c�����oi?p�c >�V������q;��G(t����Y#I��&��=�0������'x�$�0=���!Гy�-��ـ��KP�F���J�|PU�8NVc;��$�k��9�o�C�������Z0r�p���.�}$|�y 7D¢��BP�B���p�����
�ۿ���o<"rڭX���H�M��ZEf���A�Y�!Z�j]��cUGY!�<���8�$�;N��/Ʉ�@%M���b�L*0^�E��й&g�ȫжýֈ��.h֗Z�t^
(�p��0�y�c��z��>;����u[���T�qC(�k����d���!x<٘��	�%�CU��G�ԩ��WDԊD�/ ��rk�{�X:$S��� V'�8&�Б�p��*��$�*��k�z���۽�J�)�t�)��|`�L�ȓ~]
�T�@%z!+�A���UfPV�B��{�n��������D���m�~^�=�i�&�"�(��T>.Xg^ˬ 	�3�-p��!5�6m�kȭ;�h����N�r�,g权��_�gWP��S��S�\نr�M��R�!��d�=����f�	��H>B9KK:wJ�uގ>���&"�#��{������z<ƭ�杓���"eOY�FP�|��)1c�	�X���X{����Af�@��mUܜ���r�|q�ě���oF}��wX"}	 Ԥ�2zVz�O��KI�@�?ʣA�-(:'�:���aAib�x׳�"�aoN��_�.�?�A�^z� H d��Ա�rv�XA;������5����9U�*��lL���U�� iƏV��Q+��P������f֛��X4�,���G}�������WU����Vf>�hf� �s=�7��$�����DI�E;\������a���
����k7XW���Q@Q,ϥ����@���^:�”#|�ȳ�?T�_��a�_^��n^�gQ	�S��I���W	)�1��.�{2�}����\ѣ���g���5�Ze' �B{�8��j�Ɋ�x�_�=�ñ�����eS��X���1��7b%��� �3K��*0�TRt#������� 2�����DF<s <λP�6�P�yy�*z,����<�z����#H���v�z��?�*��D|�Rp�v�&׿�����\�?L��Y�O�
k��+.�F��\Z�PeGH�SL �%Pq&�鿓�#�}f�h>��qn~���ة��E�Xldit"T������7�(��u�H�'�}cyYrFD<���y���X��@��zO�&���`~�mۃ�'$z'���n�w���GdQ������R^kQ�9Vm�`�x���C[η{���q34}e��=?�����kkZ�@����QY�Г(%��(?7D�{>��r�6,�Z	������]:d&Kѿv�"�������I�匈�A7?�F��i��$�r�|�o|�3����0\�$j1���	�1��k����;�T�� g����m�/��9_ZIi;u�=@�lݨ�����A�V�`����F�>����(�\8k��9f�?e���Xz�n/xM��|*ɭ��������ՋS�%�Cwm���$> Գ�j�lAL��'`b�w��:Xf��/��{H��_6@#��/7{O΅cWdP��X}��-��)������םߒ�i�G������U����	ueHB@��֩d�uT<#/4Aؘ�@h������č�u��x�������/N�^Ve��?�k�<&��;���Sy�?s�T�5^W�t|	LIWs�� 2�*���r���O*�ѲJ]y�?�H�c�m-��M6(����ژZ�-�-�IS��[-�D�ۈr'��K'��{{�~kZ���mj2�_7M�-�?�pQݾ��`��:�c�0џ�!!J�Φ豿S�!�l�P���pc&� ���̿�T&�uy��O�xy~:d+u~�="�j<;-�pϲ[�q؋ٙv�^������9&�$/d:G#�ݍ�4��s���oo�J �t�'��P	a��Rr\�������y�(� �4�'���AVM���N �`�#�1	�O��!�o#�B�����F���u�=a�����򹄒�&>���H
��<�����Xd����S�_\�&��RC�|�	:VfX?��u<ޤ:l8s%���(�
�稩 %��;E6�����Q��߀rp�eZ�w����m�Po?�b�n�y��2�n� �(�EƦ��H1�~�c�|�I��d��\�7�
(��ZD��uG���!賜��M��ѻ�R��H��CoӬ]umT#�ً,��D �=���R	�d�p��'�#n��!���*8ଁ������ G�:���/!��=���1��-�p&��F�;�1�"��)��i��WA��᠜��ò��`��|<�΢��Y���>9 ���S�&{A	�v�("��}�Q�7O"Ym���iZ(���q���(�w��:.�Ң	�LHkR�M<�֓��u/���k�);�:*nA��T�mp�Kx@>�;�h�!u����^_6��G=d�څ3j����nO��mE�*� ��j�k8��;~��� i,�����j����$9�����"j��u"�%y}�hk4~�����ch[� �"b�����v�P�T�(�:R�#L����#�x��	6!繁���m�v�4D���)Qcj�^l��$+�dh�9Fl�4</cj
�����5��kf@ñ�[Ʃ��^�[Z>������*�7��(�l��ߓ�n�~dǦ&;.ܧbN��w�����)�e��V8ڸP(ʟ�E��g��ҵ�3|�L�f��� qp]����Ki��b�O
?�<�_� މ���JG��I�m�������D�̎���5���.TRbe'���q,��I�h)��0��&
E�l��{���q!�v��3jhT���B����L�0���?�
����
�qVU9[�$���Ӛl�����rmIC��>C�������m�M6������_fW�����)-��%o���=�)�;\@�d����$}��~ɠ���9�]�t�z�l��c����h\B�xodF���X��ޏ���wΝ����2M��!�N�;g �|�A����w==�2fWEtX"��qS��`�C�����q%���?�H=�;=Pַ�6֭%ҍ�2�v��u�/��8�d�*b��*�m���Vu�ȓ�F#kQU~��o��D<�?-B�w���r�׷2����׌5(:��Wߎ��6Ej4��b\-<�ʭƟj�Ah�)�f�\��4_��0S6��R^�9/=|���e�2�d�@<s�g�!H�1V���N�DЂ+��v���q$����9w������1d��@X���	���\[�x��{Z~���#��>�%7��+�%�L�|Ǎ�h�����F"���f#�[e#�i��_M���C�������� ��Ƃ����܈������}��m�,?�SyӴX�Fq�:7�(��&%���ۉ;xvZ3q�WN*ɗ.F� m��4|s�,788�aF��qB�y�
�-���M��/�o[�*ׂo��fFW澄���v嚶���7ҬX*$�%�����X�_��@�9�\\�Y�G����
�Z�4`�vt�GC`s��|;#V��F��aࢦ��(���< `O�ӌ��\*Gq'���10�T,1`5Q���#��vAI"�C��)H.�6K��B�F�����m��H������/'ɰ�F��7�W���C��{'߳R�JC�T���I�g^��Vă`ο�,�KÅ�j���2s~Clp1?�D��/<q&)p�*ō�G	;��������?\�
J/�W�����e��~s���.K�>��9q��ɐ-���3�h�9�%���#Նn�#8���j�	U��L�m20���$�#iJc^Zy��z�/	*k���4Tp��`?o��b��؟�!��d���n߹6�7F���5��� �o���D�uXrD!��йu����P��b��%}o�H��h+G��\�}��X�{��^*t��	F��~εjPQt�A#�=����OY�2�=�E@�HE�e�s%}rH0�W���jD���s�5NýU�����t�V�0��T�"L�P.��o<|��p��Wym%�I�!�q�U#gy��AJ���|�:c�GT�t��X#�ʼB��2O;;�!�QM\�jS��yw� �۶�-�zc$"b!W��-XTj/�00j�:
����l�8�� /L�m}���'��;v������ƻ�+b �P��l}�!�Z6�2~N�P@+�᭟��+�$noќ�7�~N��L��xR�Z+-Y�ej�����3����/ �@~[H���V����!�p�Nx��!�2UH�mo����t^�E���W��$��_�GQ��3�È�
m���[�����%�^Q'(���ki��6!��jæ�`�~��ڐ�����D.��%��_����<�Þ7Ч���~��f�7�S��
��K�������B�'�u�"���E8i�+�ס��
L�E��Є���������O�5�GK"�g��v��/�f_���:��e�;��"h��^���.1Ri���A����F�F�!M� I�� u�M܍Q��A-i��S�_[��k!(��o�!�mdK8����l�18�ϖ~���T-�1�SRP���ܺ��?>�%�I�7Uui��D@<$�zL�2�j�}P0ڌYA�wt�{d�f�&%��Ӡ
�g<�m������Z~���o	4\�C!��'��v�,%�ڪ��r+���c�x�|B�#�
W[��?�]��7MG��bU�Y�V�w=�f����C�'53�~M�y���A�}�y_+��da��_R��q�@%�:��k��B���� éGOe��s(���� ח	ۦ0Yfh�P2E��eN�sW�lG�]����q���f�F�a���%��� Y�A�
�*��������|��} �� Ā>�wNu����wJ�0���`��5ա�E�AX�"RNw�MѼj��Š�ʞ��l�Ձ0��S\���Jk�m�pP�
��yB���������+f5��q6�FMb�q�/kI��,Zjռ4��xI��%Þ�#��o&x����_��1���S~�D�E��F8�� �\�����ϥN�L�1�akP�Eu0noW�'�,������)��Z��̣U�����T(Y���[��"-CƉY:XQ�p�U����.�r:��}��ޭ�6vc:XhU��.R���S�.Rn�Cv>�jq�W�+qT$6�ā��e{���aE@T��� ^x���cI%G��
�TQ�a:.2��	�U|��Ri��2LV����2�	�d�=1��1��5��7�S���3 �j�� ��Q�F�����
�8����3�U��gL�xf3R<�� O�s|�|�~�Ŕ����[ޜ�[P��ư�NQr�6m$�/�K��ƴh=���^���fnLWB���	�?����G9��U���#ˀ��-;�+��俬p�q������͎��77��:�O���Ɵkԑ1�!E%k�1O*�,0L#�s�3�T[�6��!��Y�g�(xϗf��2�� �-�/�g5ďs ��<`��^��r	��B�6续*�W���d�gUMѭ�����N(�;P�+$�7����������{X���fI�|n��(�JY~�N�xz�
=ټƟ�o*������K��{K��	"�5�@�&sm���,!�|���#B)����EP�=��1]��{2�2N":�e}���&-N��[�����[:IC9�!j*\Z������t��KK2ƾ`g�9P/L$��)	D�m�kbol�������M�Le Z�w�}Ui�UWQ�h�&o������S�@����x�,���U\�	�=?�k��Hp�3��<�xz�lT�<�ǒ��ZD���Ho���;���mC�,�m"�(cA��Y	���74�<�)��,=3&vX
&�qU��,w��D��fD��)� ]Z�l��cG$d,dxF���t�5�z��i�|ǂ�����/r^6���gfd�#4�J�פ������JXܸJ�P�]k����������f�d��ܒ>�yS����� ��.��6l-�A� �	-��f{ra�A���ռ�Oc���3�CZ۷얔v6w�wc]��1�?2��76�t��[ �������8�~?��ݵP�/��[�P���̑z�F�>{�z @ʃ,�Q�4Ԋ��K��f�_�=�l!S	�<�֭@�|v[�5ȳl�˺eS��-�/xwu��%�a��F��.���p��[Hs�!ɗf��)u� Z$d�F8~jf�4 ����h�{�(�(	NMFG"�1(V_ޟ��w8*��J�u�oe�~�İ�c���R5���,B(Xm����s�.3[*L}��m��`�Z�ʂVRT���)��R !��6�p^|r�Rt��ӠӳL�6jY��̭0��0�yB��I�-�4���ٚ�,��U���͚�g�b����="h*�R��z9��|��Ǔ�3E����M��S���S��H�ȯ�W�	>�%�C_u��r�K������C,Xe���s!ܴhw�����̳w������D��~�id�V}��f@C��~�$e����M�RLP�;�d��?�K��0_<��Q0v��l�!@���{"$M��1J�V���+��"Q�)��]�����{���B�3B�-$��#���)���X4��ҙ�I��G$�<���F�H$BJ�h��e���>f�n�kbG�{���F�_,�����B�����S�(�f�'r�ʓ�Pǝ�������y0W)x���vF)����t��l���c�V��ި�t�)���(u�{�����o�LL�-�qۧEQ��:��E�Y�^Z�C��"�]��?P2D�0s�o_V� K˂��Ikɰjlѩp��Xa�S��Ij�Ԏ��Ʋ2�$h�)�+[���7G�}J�6�������y6�-����X��~X�d����@��j��O^�G`-�_,]k%�,�,��~�&�bE�K�����~�� �.����序.��005���F�i�OIr��:�Y��[d�_a��J	k�����{B#����SS�ߜ�	�$�2j鬠���t���y�Z�� ]��ֳ�������]�p ���<��)ݱ��&=�'�|_���c�~�۷�=��	��e���0o�n�� "�[dN+2�����%W���}t�|�!vO�J [#��P.'���^C#�����hM1�Ԋ=����;(J	pg������0krUP?�������N|T��[2��`�O)�������i m��n�Zͬ0�y�Qm`�h�S��j�j��dڿ�� F�m8rL�]�
�� 	� ܂�=j�!6g��ߌ9���ξ�>�q��M�{;��/G�d��gF��gȃ|G����28���4���4��#����F'�n}�����z���<������P$`V(���-�3��9��(�4�8��W�IY7�@�3���F,~S�I^���o���P%e���sJ��@FbN�.��kX*s���lL]y�<��C�*n���3Pr��3F�?$^��9p�M=��#x��o��e��r���`��X�w͡��#lU#���ǏW)J����j��8M ��x�:f����:��������f;ӌ��D��us�Fj'W�[m�){CT���p�-������3>Z
sP�d�k���n�����|E��X�����_~v{��DI��%���x��z=
�u��s�4�3*��_%��f���ؓh҂�v
�������6�a4^,l��?��?��Z8yO�AK_.�;LY�ӿ<Y�}�:�Y�:�A2�} ��;�x�LE����A�H���k��-G����0���}WV��^�?����.6�I����М.K�{���T�P<u�Kze��ei<�",8���.���s=�0(�M>�Ol����z���o��]� )/�^J�l��h7o�K���y�YEָ��g"�����{i}Խ5,-�Bk�P���U̴������kH��׷^ �r߻ٝ���=j��;#��ա��vm�.8�:�vF^��j�Xm�pr��;�d&'��O�rB}���fs�Y*�>j�oƭ
[�³So _��GذzQ�N:e�ho�)�t���9]� H ��+>3e����.�M�e�$�z�*�ǊCȰJc��u����R�Y0'��x��Kw��v���˝����t1�̐L��pGC�{G%���1q?���֔Uۮdjhy�p�4O:>��L6L��4��[���&-�5�*��89"q1Y�}E?~�{�.�)�khmR�>��8]Ɣω�Q�J���?P���R�ʰUV`\A�]7,�i_�">.��]l���/]�A;�����a�N��4f	oU|l�Z��9�QHF/;X�1��A}5�(|V�+��8�%&�kN��[�+����F�j����~�Y1l�.xО��e&�Yz{+� ��<S����i�"�"
�{��ގH�Ur�WA�S�1�՚w���m�;����Z�i�:�s6�u�;�`��L�����(����I�z��9�SP�5u��2l?� ��L�Nˎ���+֩�_��xc�`(�$�Ѿ�+�i������V�\.�
6��@�:����*�r+QqA�����9��8
�[��?V�v}����p ���|9W &��̿���xEh�~#_=�BY���ߴ��'nJW.x�4���dڽ����wm��^&���ރ��L{?��%B��hO��5�)�Q:���r��;,�/���µ,����v����8�Q1/�KR�K<誝CFmН��s�*g��I���1i�I�I{�E���27}1�3����=���07\�M�����r#}�cPA��$�P0�����<0����ߝU"�[��޺�Uc�rZ	������\���9$�1%�E���ɻx�:�/*Pl_65I�ޱw��&��=����\|
!� �7gѨ�����kw���������č:����"!��'ԛ��W�]7�4���
M��b������jK#?ol�`�/L�y��t]"�B��$#u�SV­}�}�����xG�p(��'�@���۰����vƷ���*eFf��!)��*����*Q�̢��
��ۛC��4˝`������N�[��&(��ʸ�$�;�$�_�q�heZ��/�ށ9��#��Q� �x�:ʡ��d��qmHQ:B���kt�Q�䟮��:`��y�ܞ�d�T�!�����sk̆����B�M_)�7�>��{���*@eH/�^��|kd1�|<k�$M�K��#ld�+��'H�'���` �s�$�J�K�D�=#Hj#���c��z����l��#��U_��\���X� b�`_Eg(�IT3�Wc>�U#Xy2,QH �.��谷�Z,/��WV����vP$��㕞ec}
�x���6��Z�?������џ���),����2���0�����ʿ�8�.*��T[����/�\����͠��o�+�z��r^  �����{�.�\���I@�w�wL�8%Z��Ń]���@�t�u����*�4@��#ҧ�4�W�Kΰ-߱���]0 <�x���K�u���3`�XѧY��C$k'ڣ�P6%��t߇�N�Jh ��o����4����}����?h�B�ը͊U����&�h�H.9U�L���ג����*S���J�Jםe������{.`���-ԭ��C�af����_T���7�V���Xie�ζ)�0��#��az%�^ϖ���Jidc�������p̷>5@�����1���:s��-�V��F����0[�B��/MR3���od��Q'��w�4�$:Gw]`����FQ�ė����X	�9��_�����/X�yW'��� �2����qi ���X�4�fC\ӵ���fy�r�ܚ��n1�MX�g�O];A F���_��Ƀ"���te�u�V����ܺrex�X�'	�.������M�b-D���<��w���a�+aZ��P���L ��*�T�]���Ƨ�8�?WV���J�m+/[t&��)�!�t���̙n�=��^���=��\�TQb��������2��r���;�<���8#{���!>�D
[�hr%�����d�����e�l�X'܂���?��"� ��j��5'
���}���}���k��R�KҚ��B�ܿ�d�Ƕ"Q)�>�^���>e�����E�����MW�������m�Ʊ'o�SNN�y!"?b Q WP����z�W�|H�g
��6�#)BӨ5�LRdU��~3k��zG�����D�T*�����Z"I*��S:�Y�����F[|z¯���N��Y��i�] �'S�]7��,�k�*���戧TS�Vw��j�7�d+51!8GkctQ��b\ ����KN��4����X�_����~�w�;��2�Ҏ�Q0a;�UK�GW�_Cn-�{�7�)c��hԐ��A�8J�v�ɻ��Ŗ��e�Bf��Q$���t�u=M���3���L^�Rպ���J�~���ʴx��������	�����_��@������ ,54�Zρ��X#y��K�{U�LTtis�����ӏF�T x�E��-~�28��^��۞�-f�`�5y1X�LE>T�i���~G��"|�%��m�ͽp$�����o���]J��k�cc�i�=>t��z�q���Gx����\����w�r�����U����Sq��{�\�.�E�D�J��ڧ�J�:Ӥzj�����3Yf(�b������{�yϔ���&f?���[�r��wP��t������c��!�5�q�8L��	2�qCG�$����5M3{��ZX�%h�S�ڐ��$��mľ|U�Q��ؼw�qR�7����\�oe>3x��9bl�y�8�/N3�[e��*G�t7p�J�.�K�f���6_3oʷܿ,����y�����=���*	f�ի���/V򯈧qV��_��^�]P��<����_ ���l���S_��F ����t
Z1�P=}GZ��&Ma�=��%T?}B$���j.�Q����աZ��ϸ��=�w�4ޜ.tG�W+<�CV&�|ᕦQ��rx���fhw%R~UF9��s4�E��g#�E�d>��JSnZ�:����uP�H�1p�%�ߢc�jX0�kT(\�_v9�4QQ�L��?k����j�ˌ�H�erg!(���p��w��(�z��5�T�M����8/��%�o��R���j؍�i��a�~s"{j��3�Z�e��
��FuM��Α���?貃��K�2��}�������B5��d�X�!�s6$LN
�@"!�f�c��� ����%輆�8�$r9*M#Y� ���cg]�R�	�6G��h����0gB�������j]j;����%��=ͷ���H�w#��x߬�>�db�pv�ZZ��n��jr6��N��9�[l!���;�Q=��
��Kj�dd�&��n>�7�֙O��o�*'*	�[�`t_G����h�1�<��f��bxG��C�|���z�ױ�۽�� ��G)6�H�Ϳ���m�� ���aN�ʏ���]Z��h�A J�2���ڭF
#)���g�<�>��߉�c��=1J@Γ��E'��,l5;[k�kM��,e�%�z<�V�m�:J��I񎇍?����_�W�0E�l��Z?��GԸR�����3��{$���4M,��*�M�g���Cer�\�-'7������E���j�rC$�uy#�������h�����@�A\N]�t��~)�O����aF�n����a�Y���o}�#?�J�b�A��sl�rY�r��E���F�<���;	5���#9���_�RtS<���'����Fu��a*(QhEY��
��Ql�8���E2���Mf!y~���]^Yr�4"y��O9��#�P�AR�k#xZ�a܋����dA����@)rx��!�71x�����u���: cq�O��*W�R��]X ��fa&^�*�O!�xђZ�R���&|���!����k�&�}�47���'Q��/�w�GLQ�� ���]�H�å;^��gB�LqZ��uz܁]V��K9��A�TmU��TF�r@�I�*$���LG��g�;�\8h&�H�5��vU�|��Z14��;N��uD����>h�}W'�;	n�I�h]�]HT�'�����L"�F[�s���i�1[�6T
쫊C�z��ڶG�}��;��M�k&��S{#r���"�Ƞ�z~X�Z��j�@h*IX�6�x�8Y ���y���}���jhd��s�RX��:�dQ敪��}^�;}�p�/U�b_���A'݁:4*��)�h��>�Y-�H �R�v�+S�s{Z�M=��}!wQ��e>J*A�ػ�($dqF�]�A���R�e�S�N*l��Hކ��o�aF� ⚑����&�#����8�TXN�[�
����b�Ji��r����/�t5�?�h�9��kIYBW@��1�Q�h �h)����b���J�i�������wL�H�W�_�:���ʘt�?5�ɉ&a�v���~��<33]��NU�c���`��G@=NPfH8�?ћ�N����1C��G�J�dV_�o"K��;���s�'HQ"L�s��X6o��ZӾ���E��/,��X�.�).��`��7�_���d&�\�f����$���ϖ$�f��.00V5.X��x-j�{iA�ȋHS�3�S�XC��nZO�@P8�Sk�DE\�F��|6���?��8Y!��E(��-a �r�ᄺY��̂���99�Kb�J)@=�jC޷ch*T��7^�����xM�UrНK5�sq�T!��dH������<��������~~�u���LF�����lF����ᡸsYLl�pޯ���la�v���UW��4���b�{���X�PS�T)����;��*����)q�R;O�s)U4qc ����4���Kk�8˅kC^��j�A��U�:��x��`�����/��VE��U@�ju::�'I�9�Icz̓I���\��|�n]��)_H�T~��nol�b����~%�ho�Q���������\a �ffG�"<������Aƫ+��Eo�R��2[�ə1�>��T(���_�����֙V�?Z��l�Uz'ew1�e ��9r�o7��,��Xj�xo�8j�.\�j�KCʱ)WU�4�z����}�p#�fËl}�$2��+�0~�oA�>/��l��%�rJ5E����7�2Oc!_t%�+�iK�;�V+/$�����d%�L9{��kp��,�C�nd��e�ϼNN�L�H|E�	��O��Fz\*\�����ǖ{���Ϸo 7f_�| #�_�r�e$]Vاb.a��չ,���H*!�+SA��eTE�y��iM�L	po��U|�:ڡ&g�y��刬 zQ�^Z���=��շ�����8}`ز�b�IM��"��B�b�r޴+T��z�'�?��M2����g���@��
B���U���5`d��[J��R>91N��l��r�i���U&�38���v-3d����qB
3���T0��l���n	����{ ��0���-U���q(}%J��hD�.�C�-��̂�Vſx�U��2���h��-�.Mg_mH�A���� �n_o0�A����;�E��/��a*~��"H�{� 	P����W��-vn*`<���t�����ޏ��c�+�N�����J��jXYM��ĄU���/Zw�p?����܎�/-)�9���	��Y��8�y�����Y%��U�M��e/���!��%�4����.ٚ�_����lEa����Q=&g�B��K^u7�W�-:��s�>0z/��S����@��J �3��]t">U��[Ij��m�1،x�i��8y�0�׼
�g �hp�4@뮧�e��������W�B~P���iZ&�_�p\	�=��FQ�y4j�c��dٜ����wCl���uN�ۦ@=�ط4 '�ڤD��$��'�YqM�*8��+�����Rߙ�t�H�ҟx��<���
�Y��?u>��<��&�U�]���%t�.CaS<Wc�W���%x5p�?h�`nM�Xgd5���y���17��B�~��a��ǆ�Kh��Nr���>�:"��0G୺̤�����,�*���+�'��S��~�1-v��vSjHז���cS �Pj�J��t�b��� b1^d����[+�$�wj-Y�� ���OMwlRM�������
�YǳaIJ��7tvMv�1����9ႊ��Ԡ-4e\�}��-����O�g ����3w����}J1�Twxҵ"�6�� �J9��u��'
��;o&o�VU+w��-�;p_��=o;f�iy@���W�#)2�]h=E�.�m\�i�q�Z�X�1e�B�=ã�Æ1U\ޚcM�;*}�8�;��F@�����k�}p�̕�uҩ���2q���K���4� $n=h���Њ��P<\�aj~<�N0&�袻+�U����?-�b�N��7��g�[� 7�Gm�"?H��?m�mX.�V�
��?~�/���$��D���-�/���3�s	��ԟ/'���n��������J6���m�b9_Ytw��h����KO(���p-�kHc��q_nv�]R��A.��D��F�����U�|��O�p��Y8Z����Ё�.��Bjsq~�@�8ApﱺT�8##��V�0F���]��I�a�I�`����g���B��fv1�"�N�
���&U��_�/>�'�L跐�j}��dXJfꌉ���[��/1��I2U�0�35�!tӺ�\��"I�<I�6g�l`2����0$�W�-�D�SI���\�j�~��Wp�0��ӬiF$���y��Lq��z�����V*b�n�����p7r9��s"Y��CKl�_���NZ<N���_������P3n���4�Z��8��i�oS�u���T��ɤϧL������❈��i�+��'O{:�[L��7��&X,C�J�ED$}�f�a���X���V@�:�ˈp�?��IW�-��iu�+�24�ʧ��FzC�Xr���)�*;<��0jm��xg�@� �c�l���~bbi3���ҫ�g��ܠx.�?��$���� �H�C��)R����	H���,�m[z0�X��'o�.��,�ܡ�,��"<�������'����7v6E0�{���3�v��c�_@@��IG"��4g�>���>v��-l���s1�[.������ ��!���ژ��~�[*�b�+�81��x�0PiOX���}�ny�*6�z8�uQ�ۙc���[fA�|�(ٟ�T|�0��A����jh���ɏsb���T˵^$!�T-mG�[�<�]x�� �/6�5.j9��n=����h~��H�H�I��x�[�^GjO�};����s$,tپ�J��� WܫR��I�Ȫ?���MD$*�����?-6�F!�\��pb����a��Pj]㓔 ��A�h�!lqɦ����o�a[�M�l���!u�)Bn!R��L"i%��Ծ��&Z��53�˨VH�+�N����Ǿ����u���P�٨��|v�NO���B��G$�g��04�{rO���oI%�7�]�ر�ث�D	h��'���QwLG
�en��U~R�O,-+I��)[���!�]f�w�4c�y/��u+d{�����c��:��ܟ�M�lA�xR�C�("�	q'2C�44>	���d�M�B�>�EP K��[�����C�K�' �0f������\�޳��������j{V,�ӽ:{umΟ�`�Hw��5 �XW�kY$\�.��3gG�__�3����7�!�i�dZ�v�l��p����#�� �OMA�Eo��1��z��t�J�L)*���!�7��Eί˚�^U�������w��u2��F�P;���U�����b��~��kZS�x1@�
���k���Q�	; h���#8���]M��!������Ԑ�����ׅ:M#�~�[Tm��/e�������~����UA��H��):���z	���ǄTDlsT;���)�P�4�̗u�T�2�VǶ(����5��~�,-�bS#���Z�k�@$���	��9\�X�E��V|��5p�5�P!��b��-y�%�c;_�Y&�i��GP�3�݉�X�l�%��t�Y�d���UG�4+2ӛ'=�N�w�s�3�/��b1N����<ԣ�d��h9l��߅1�����/k��-:�dP���b	�`��-_=��2��v���4�>����ܓ` �eb�����y7�w�]��Ɗ�\TK܋ߵ^^Y���r�V���D�Cո�*B�P��Z�.�fys�O� "�妴Af�eON%�/�
�};�0^�q��[Q���E��X=�%��0�ɪ� �3����׍r0#f�V,o��Ɉ���h�zH3�$�~5�vm���KP�T{���J����N/�����D��;
<������pL��R�!>�>����A��v�F�ΰS����a���|� P�n�5$u��it��S`� ��'&8��x]�gj�el�ʝos�[�=x�d!�j��`>�
���~R@ �#���!�=>�:\m)�<~��/���[*��=��Dr.�X�Us�c���H�M�z]V5ҏV�ߔ2zX�ƌ�]���D��Z�#P��WMd[m��=7���47��L;Fd�R}F�X{��P�e�5f�t��LR%zB�Mk�o�]���koѰ�8����z5Ĭ����:�GV���������n��VA�������x�X�<R��S��Tj*taY��:��t��I���ᛖ�����2k8�	�.��%�����+��.a���:���ɞ� K`�P�bnTS��j��2Ɂ�l�Q'z�&���l��� `�m�1��8��6m�?Bu��~Ɵ��U`$��/M]M����r�M�ǯX���ې�d���m����ͺ�LɎ�7ɑ��
ӟ6��ZJI�.�h�#�P�^�6��]~0�����&�2�ᄽ��%�3�q�m�ABC�Y����8t=r4����,����}B��1���ek�,8~>Kw>��05⛽��F��2O�� YµŁ��i��Y��lF<���pR7n�HX��-b�g�>Δ��%,��C�7l�� 
�m mX:�U�f6��YkiF~�K<�|��&�����ۯ)�1�Q��O��6l�֖��Zٽ��7�T �ЛH�f�ѯ�.^���zbn���������NzݙM�:+b�L!�.���*���'?��7A,͎܃�UnL'0~ݏ�~����Z9fl��/)����HTQP@�p,+1�