��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jåا{�\�u�?߷�dn@6�zf��r������;��������W�a�ٲ�� ����k@o�^����44W���n�ү@2��������6��$kw� a��(A'��!�����*�������{���c�(	F�s�nHL����0>�̾leiA��i�3�����q
��Ӥ�nύ���zL�m�FǕ>'�b�s�I/�Nf�j���no�O.�1�Bw�f,���U��o��][v��i�4DO�O�:��GK3׍�XH
��#Z�|���k����M��~ǵ��?�-i5
L-NE�+��DYԌ�x�f����疀>8�l��db�����.t,��2?։&���Ĺ�&��W^�5�Ը��|�I9�hA?q�G
�(������;L�3��0�Sju0<\ڀ�pZ�[^gv�Q��/�̦SU<���v�	Re����9H:�i��N���,�7TiW{�w�\�G�~�PY��
�{Gxxs:[6z;�(b^�Pm��\�7�S��j�&oբ�D�E����\C$⽣�D|bLXv,�QbJA6�dGcz\$�#�cO:�:QUkQu1�D��n�A�ց��A3)���@�&�H�j�g�z`�����٧���@=��Xl޳�wss߭x5{X�L�l��yJ�;�����l5��u�����ד�v���:�ʥթ'�!��'�����:֨߭�.p+�W,4�M��@�폇���~)us��V�(4����ͦWc7L��o�pt
���1�%�qĎ��'����G·%^1w�kmGjAR��j���%�P��������E��O�F��SDO��J��ޟ������˺ܠ�z�m�4�u��N��nS��E,R-��hZ#���6���}���j q�7�_G:Lc�t�8��H3�:��HoPf�,Z����������5KB�z։��t�ú2;h��o�@������UѢ&��t�� �L@N�?�n!n���/O��=�*�>},5��Ǆ83��0�J|*�
��I'r�i���Z��ttP�Z&g� Tb4H�����@��ɤ崕�7XM}ʒ�.1�P�ڡ:��{�@�|�?�[T�=4j��:���O.���Z�� �x�x,��5	kٖ���m�\V�Tgk��������»#��T�"QP�mycJ�`v�����X�ei���R�_b�lu�/2�����i��^
����f��s�"K@3 �ŵ��Z+����Ӝ��"Kݏ��N-r��w�,��䝼8�2Y�������	��<l�*��6U�k�ś]u�$���~�SӃ�X�Y/�w�i/Z�(L��������p��.^H<�&`�R�փ�a�*��B]��o;��%�ʽ�hмs�
~��_���^ؤ�D��2��F�utS��j�����("�������?gc�z�>1�,�~ʫМ�TP�W��
蜰l�GkG��2�b)��z�M5L��B�����Xb��lu�eLzK=,Q�<6:�!�qB�����>�wr�~�t�q�����݈VܼgRe��=����VǨT)ҾR	��u2r3}-���
��F�_��c�Vos X���b��&%H��>���gې�_�c�,�	!}�x�ÿ�w�B�Ġ|�Ζ�m1�ZK�Ȗ&����A`���W�4���U���������&Ø��ā5u'���B�����/01�cH)6f��a�F����,���(A����o�v��y�*;�"��Y��}�m�ڷ����(Q����C��Q��As)Q`�8�z$TU�ϭ��6�m��J����KGA��_-�_"�cbNzS]�e�(���K����	�P��[T���A	OVT�S�`M��7��8��[\��,mwPT�b���)�������캙�Ր�>�CX\Z}��F_� N6�{p9-��E)�,����xa"�<�f��ɞʽ�Y��K�L��奨��[g�� �2rS�;K�+��ȯ�����ї��	��螼VB��*�#�t��^t��hs��)J�ϵ�9 ���q_��y�(�\�F���J^gY���8d�BO�+�N_K%��� �~�ܛ��禾<W�,�����4=�#w>g���\V�?�
n6Y��k��z9��-$�
8g P�Q��H��Ar�qC��Lأ9�ZcÇ���lP�G��;E&I+�Q��B��䝤�޿A��-W��爼�)����ǂU��e�ě�������oʃ��Ԯ�~������kl/�M(���%�ѷ^����c������W��G��/��kϏF�B���{��Tj)�г_�P<^���f���Fb�_��ݝ�I����ʻS��bh�M��DuE4)���<�*"Zm&����n�׀YA,��2�z�������d1̃��!{�0��jO�d��翬h���"�P�w����欕jW,&����<�92�&~�)�Fl��Xm�	/��R\��aj���>\���oY�)��Pi:����zT���:g�.�O`wq����JW��ˏ;K>}�oN�)�\��v���+�{�kWy>���a�j9��saM�+s�d�-�tVa��;=#�dbDgi�_I�0�>t%.Z�3�H=�VP������^��Q��`�;����m6�c�a�{��v?CRB�6��_ɞ{j� ���e�B!��RL0�>�8����������9haC��sA6c7�w�#��h3CO�Z0�	�0�S17x�V�_ߛw4�4���0@�Ő���+P�e�k��xe��<���{�����z���vO6�{�7�\e�ō���s鴎�� �ë�Wϐ��c�#?��4Һ{���avZ�Ub��:��-yF��l8u�qA�s�)BDS�1=�JSX�}'1`)@�����aX���sr%�u4�?Xe�<��=6�  vJu�O� yT�r_A��E����]O����.�$�d����$
=���A_��6��*�n{C��R���.�A�h��2uzuy�Qe���Q�H��_�����ğ��X����gg�{pڼ���m�(9�(h>W����Fʢ,������u>Z&:�\�:�����Cn�{˷��(g4�"I����$�����#�ӄ�m�P~*�i�����ip����D�b��K��=��J�������W�	��'ZWrL	N>�J��ԇ��ׂu����� �J3k6=��~��зN���3R?��u���l`"IC��L �||�lF��DS�,GI,G������6I�I�i�R��Z��j�	̲�SHw��
�'\�ؕ%��t�,��j��3�R?�}�V�%(nQT�Y�N��L�v���/�.]��壪�`����z��-��6�.%���05��U�r&���x(�(��XAt�Cş�ۢvѓ����%��qŢ��A^�-��=�1�Z5	�d�G4�˟�yC��j�b�4-({o���*s�F�	4��%w<`{g�ꪔl2��g��/w��rY���$���:G�P�
K�=;����٪�x/5Z�W�}�RC���K��Q�Q`+\�����۹t������g|@�gr�Ǎmn��"C���W���z�g$k��&C�Q+�2)/�1����qC�5���Vu�ː�p��d\���N�0�,Q΍��(�c���Ǎ�Ez��Cq�[�R�+�]����{>4�5y�0���o�ƚ$�
��2�����xF�[���	D����3�L"/U�>S��4�)��\9lp�!���qx�F��T�꜕F%e���]>]��`�;wGT�:��!�7��vpd�����_��ő�g�D�+�ou�Hw�2PNm��Ik��Y���>���oun�����I��`��`�׶v���-����~�0�slf'����H�mN��|�l�$�$��X�SM�0ׄˊ[F���j���� ���~s�)_Gzk�_�IC{��v�"d@6`7��ƥ`���:tF���A)�̓������"<�"�L@��IR�y��NK�@��%�(�π唟ή-�e��������4�Ů7�/�7xP�w�3K��j��"�j���eQS��ç��HY�R���7�݅�(�3��Y��$o�"��,�>LS�z����t�u���qf"��.����[��\+u�1eÊ����oY2}�
�ɈdP?X�{�oq�`PNe~8x�Ҍ�wΐ)b�,��;�
��u�z=���DY�.3�lv�^*,O-��1)�䆅x�B?�6�]ՅZ���}fÍ�l���%5���Y2x+�p��?�Ok��E�[�e���n��I��9']�Y�i��Ɵsx^�0�ޣ�N}���s,�)ђݥa��NI�/q��cOn�o@�(U��~�,O�˭q��[�����)����J������%*���r2j(�e,S� W��O��PZ+w_LT�^P��,���ӂ��Pi�����o�6\S�>ǐy���e�˹�:0u}��g��P�'_�)8UV*��$t�����+|����M���!]/ըl�e9��R@�#[ۊ�T_�?6D��o��|��;���x�	��V�S?Ui����Р�7;�g��f
!��I\��������1x�_��A���ˍ�*-	��Pv5!�c\r!��,�?�����ӂ;�R��C�'�p"o��j����x��Ъ����K�?
p�ʽ7Rph��ǟ�CT�z�(L\����6\Ԍ��p�OϏ�����P�G�N�R�5��jq���tMHc����Y�����W�*�<���8�`����"���5Wc�$U�!bi���jN𔝩mF�ס��P�}���2����و#���TC�U4������<nX��A	kl���A�<����2'O��NU��n��Ca��/
_���Ҝƿ,,Tk���Ӵ�u��>�\R�,��M|��1�Q�kFº#��	�3.�~�e�D�Q�2Z��n�ئ���@�<��N%�P��]����Mޭ�U���p�����Wc���S&OkQ/}�o_�1N�;���8�hwʗTL�&���O��ݲF�7 �
{r>��	���j��J�{P��.\e\�O�J�N�9Lx$�5��#�x�{����,?��ܟz�b�wr���k~X��-�z�P�LZ,|H���F~�y>�fr~_�'-n�ijb,a�<�k{,'#�=.��%��{�O�1�Y�>�7�V���Cg��1Z:w.��ϑa�7�t�䵩2��("�H�Q*íoXK��V�����0�i�x����9s5�Xr �i2�s����3�E=�<������M��.�.� ��oL��`����<&�D=T&�z=�p{y�yQjR_����u��|O�1b��C��#��*"�X��a��+j�*|�UE�6�yۙ�.���H�!�|ğ$��6z�M;�SP�˚�4\��mv���AP\2?�N>��� �835��i&%��l�����R�ׄ��"��v�B�,%����n�W	2]��Hԙ�x\ݱ�0]Ǝ��$ ��(,�m�KTW?�xj^hh������\p�y휑S����j��r��v~��ō�U�)<V�L�e�D�����h���.�(Gs���6�"�A6�gg���Ib�-��l-����7y�7|^2�Z1,���c�9��K�yd2`�T���iĒ{;TXA1�߀����Au�#�G�EI=G���ٸ~ޘ�_**�������4N��z�kZ#:G�je����[��hn����y'M<�Uy�d��s�n+V�c(�n��1��$.�T��ߨ�N��W�,C�V��:�d�4.���Y��r��P#D/�t�(Y�v�5�	l���_��L��R�Lq�X�"��y��B����V�g�ځ$,�� {oI|�MH�7V?S$x>c�e�{:L
��P� m���y��UV��?�k��5M�yE�ȉ�����k5�)}��1i���L��tf~Z�oH0�4�Vt��>�n�
(��6��a�'h&�<�ޣ�QE␫����<fzF^C��G�/��B�=1���=U;��*��������Y>�a���[QP