��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>,M�Kߤ訯.$W�7)���uٝwl׮Z�+#�Ɍ�1z�m��rj]����
�x{�!&�J��zy����·��e����)Sέ��lo[|�kgP;�U��tPs ��-���?�s��(�#0S��(=b��ߓ�"�YIl�xyҌ������=�c���r�u�OMU�C︴�N�U7�Q�V��o��O[����Һ�ؘlϬ�����L(�!��V H��QXDU^�hQ��M���J��*\�z$B��\5�>�' ���Q*���7|8Ѣ���9r�g���}sw��e�i�~{.vQ��"׼	�~����m�o8�<��[a�$������W),���TX�'KN�zS��?%]_ �.�)�Iw��ϕ�����J?u-'�Ow�8і�C'k�VCq$�3��z�����^���O��{Th��`��'���EW�B����(�l�/t�����ޕ��Sv������cE*��Y�\�ɷ�<Bњm� p�v�2��P�P��c��Z��˻G��O��з�	h��	�H��#
M̓��3������������۾n�Gn�|�]��/�p�h�����O��9��a%v��aN��(=�i�?��H�ic��M��NO�lm����,NhLj��@�M���7���񰈿�Pq��Klȇp�^Zy��G.����=��"�4{���wle`�\�!`Йj�8����j؍���&�gE8�#��37E��T���;)���4S-;���5��,�?=ޱ?�u�or��2BK�\��������3�ruyG��8��{��	=��q�~\��0�b]�e�!=8X?b����G>�j�Ee�Y6�P��TAU��yr�hs�f��F_�~ <�pk,��n���m�̈z���Z�f^?ir� o�����E ج՗�P�(����NVi������)�������j�?uu����<^��n�w��ߢ$������#�Ba���y�V��8�U�T�
��7�C��%�U<�G��+��=i~�ǌnr@�AYt�w�/�$f%�ݴ�^�K��!mb�:G�|w���IH���]���Л�e��y[+��W2�t�1uĒ��T��m�����2%�b�1pպ�{���
��VN�9 :�z��h]�U@$�,��bſ?��MA|t�Tyzz�}���^�W�#}���8�+S�C_D�6�C�G;}]D�5���P|s� f荢Vv^�4�Ҧ�]m�ާ�L�*>l2 �Z��K�8/���L��恆'�t�7Z-(9��4-▷���p���U|S��QtQu}��)��;�!��?z�NS�~����	���;�`0GZ�Zށ�V?�>!� O,w�U�'H) 	�kˑ��V�U��ZB���2s�G����,�0�d��B�'19>���XM�J����ϴ�l�$e�<TF�E�t
��p�d��IT��ξ5����΅�U�V�{�7 1V���-��44E�q�S���1V���%^A��;�'�8�(I<ň���R]3�M�{/C�d|꺼��s�E"wr�H��-K�XWs%6A_1`c#k��WB�Ӆk���Y*	s�?���G�pJ5��4��k�f=4��SF1������,����F�[Z�8W���9p���Ϭ��T6q���yp��j/=7�4�	��!=H�W�^��3P��� ��\��s�[�/4Q�K�t�/oC~�=.��?x��#_��`u�v-�\_��`yP�{��8p�F"r�5ze�Թ�x�v��1��*���6_[]��t(>zS.b4|�S=#Q���1u=��?>,^*�֫�;�(�7��^�t���:�<�>��7�3�y��\�sX1f&?!��:�ĝ��|,@�weVe�`���w��tL�(`�ݲo�f�@�o=v����/�:/wG�+t�]�����E��Ӷ�<��VPH8�r[��S>k�K�@?l��udd�Pog�C>n��G��N>4�� 9�xmPPb{��^C]�i�a���V�d*袯���8���ZV�l�? �Ƭ4��*j�2'0��8��h0��r�uz+0=1�ʫ�6
�����\������L���:>��}<�Y�Ɋ]li�fa��3 xHm73���T��I�ѓ�L�U6����э�B�/�3hd?�:��q�rb���l���v#�~7���8xE���S>�ޙ���k�/ǽkn��; � �T4�܋�^QW�]S�j�o��xXFC7�s[�ӛ� �L����2a8���q�kHfHIUUk�9�^�+f���=��<�=�q��-b�)���=|Ig&�M��|�!����U���{�̐f�i/Au�()YQ?�Q�*{�
Ӱo0�ʞ�Qj�����
a �WK�c�3q4���J��HoI�����.�w�f8�v67;�C_j��5~�i�! �9t�1���ɹ�m�_;��>xd/�A,�0�+{�H��q�sL��;p�1�s���,�y��.���K�/�Cj���ʄ/���!��q*���F����Yz����[�Z�V�l���>Â&���8y� ����O�Y��1]�����U������OӰ��̱�2�vۺ�� k\94ρ�^�nB�uy��`��b^"�kf����3�w��=�7Ĕ��G�V�oS ���~ؓi�.F���`�)��ܟu�5W�{:qC.�~ ,���J���R����5Ul���l�ف#��n�e��P�=D����A����u��	��Ċ.L��u�J���59�"`t �� �kҭ��7B�z���� ��epb��~�R���xW�B���#%&Api��%�b�}�dYS17�<��!*���f��C1<c�{�Ǭ���a5���Y� ��ء�'4C�Q�5^2/Q�6�M�B�J,�	x4��~�A��-ɤP2��ǘ�H��ȈI3ٓp��^��|�����Cg�kLu�׳��0��VO��A�ș:�U���L��e���V����h�G�8]��[{�47�*�j�z�y���Z5��#N�".A���~*MLo��lpy�s;���X��KR,=y�\��֓A�b��>1���j� t�㼞��`O��{�����K�y��]�>��8XeD��7-l�z�;p:!� ٗy
��"	������$����06����7���g�Q�~S8܃��8�U��7Ð1/�g�gֺ8p����M��� �C ���غנ<w�v2.��`
��Io�H~=��D���k^�*�+��v#��$���ɚ��Ã�0�TԼ=�%�<���������a���>�Hx���A�B���<�c���>�k�퍪�����P�_��q/�y�gz%��U칑�ݵCTWw����$.��'��`!1��q�ǡ M{RQF�6���b�� fK�s��
�MH��*�#�k{0l�z�̈́�\}���(?��c�d�_0�Z�񮟦�x;�t�1&����̈���S/�  G��a�n��<���ж�Z�g�e�4ȝ���U��,���ʩ!!1`�_��T�_�"҆��d=)m��)cd�H�����؎�1�#Wa@���3l]<���º��!�{��\V8ЊA0&>sJ�SUh���޽�0%�0��\�6���,� ��]��AM�H�()�a7�n���U���E/ ���\ף�Q����s}��H���b�@�,3@�W��y-"W�R��&��v�
��^�I ?����tI�"F�-@h�r�2gm.�X���H*W}|ߏ\���5ѪA�����-m�{^K$�p������`�V)�sr�"��$�~��ix�>�P+_ܬed���P�ң	�x@b�ٺ�K���n����Ɛ��������?c�nX�_�pyI����_��Ў��<~���qeĆ�������we���]^�b[��n{�ZY����EJ !D�W>���ԓNZy����HY_��V0���¨Ld��b.�N//R$<����N�C �Czi��WD�@ ���_o/fݯ�T��B~K{�ih:>^����n���/���Ӄ�	͵�x`^���{{���D��T�A#R8<�����g���t3�L �ti玵'mNQ$.e�*n���l�9����:orN�C��O1�uɠ��xR�LF���%�[]�ڮ���GRjb��7Ex��h/t@>��ܥiB��/�c��s��x+�#�J0Q�e��&��Rǯ���ܕ�y'׻����%1 %����Ȣ`O��b?@���9�D�rxp��$W�&�IVl�!]2�B���/�q�R٧]�P�+�D��e��Gi������y��1'���N�ECE��:=�y	���p�%�{j������|1W1`�́U J#��4u���N��,����k䳣nϭ��c���W~�t͆v}����-��NQqTV�P�tu�Ɗ����8�����%���4��@l�¡������dw�f�U�ѫ6.�1�;�5[o���}f�_Keu���*TR�^�c&=��$D�^�Λ���(��������o�[؋�g#	SL�g>̐��rN:�`%U^]"�<p�����&��,5O�jB!�99
	�4�j]��k�aOA����a-Z��T�"�m��0�T��53��󄢟d~����]�{O�3&�\�/z0'AG/CϹ�bҪ@���pGR.��(\o��w�}0M݈��w�Z�!�?�`��O���;�V���xf1ɂz"�ђ�.,.�"��=&��1�Nε/]w "f��wi�"�-Dƞ�T�����V8x��a<�'k��y;�MֺT�&vλ;��� ��E�.�"��b&��6�8NUt�2N5��O�Y�0���<c=��/G��B{��R̠��<G�Y�&S���6j߁�K���N!*,_�D���J��e�Y�kǻ8a�2�e�_�w����e��E˸�x��&�B������gA?>]��S�'�y=�$��ƥ
[.K�BE$�N-M�7�����7�'��t��<�=�E	�U�k�1���5/�1�Q>���y��`�T�����,{@�^~���娣M��Vx*)�����N�|g��a R>覭q`1�R}����c�����P��;�@�F0
���iTN������"�AAؤ�)88�b2�H{��i[���n@��D���le�Y5����C�x�y�����B�����"�^�m~^��i��k��K���Z�!ߝ�m%�iް�֍��b�'���N�|����n�N����J�4K"�;�����@Aڦd�`R�+5�>�%�2T�=�4��7-}�jY�K��~J����j ����,�����)߹�l&�o|�#I��s��ʭ��|aȊ��M�s�]J>9��5f��5���C����S���
�mj�M�laoU�.(5J�%�%C��.0D����Ts����[y#���@'ԝ�K$>���=|f�x1�H��k���,���7R��~EB(�[Ԭo;��>֝���0#sTDI2,�1'���h75h�)di�&��\�����|(�.�-��K��7N!s��1�v������e���,�t�<�Q��=�5�AטS3ω��k��@����S��n�|���]b84o��ܻ�S�G��G}?�WJ��GwP@�5>u|���L�d�b�I,��*��{��W׻a��ݘ�CnWo��@,�ҫh�����g
�%+	�A+���9H20O诺�a�-�I��QDE���yKnW��" T�i�!��]�D����Y{��F�����]}
�^]T�su�R�Q�`+�O?~.���o{l��m��&��a�y�` 
.N�VI��A���䴔�ã�3�O�[5P�Jֲ(�h��kaܐk��@)=ʅ��I�g���uW�k�33���ZȪY-[9��D�a�aaX�R8~��$�:�fm\]��}u(�ձ�� ߏ�4"֭k_����7U�?�\\~`q�}�"�\o+1���O����$0�uu�,�d@%n��
f� 㙂�j����쉓�??����-���HH�Xw�c+� p�D�3�;�0Q7�W���ks����0t.(.KO�8����e��fj��{ 覦���K<�;&��9|#��A�T�T�Q��[w�7���t��J�Cl��fA�����	?�.	v��Pؖ�2?>~k��w5��}�;�/.���^=<>=���Oo+�Hr���um���D���T���n�l�J�s�򦳺�����0Ŀ�䳷�i����;�lf`�����b�q�#QrI3U�̗4nH֖_~�[2�+`� '��N�0�yH�1Pa�b����M��	�W)3����TpNJ_r���ݎ�.��
�gg�rM�Ừ ���`���t��T����R�f���QX�S)���i`2�P���Č:%�}=�[��ڝ�	u
��,��x1�a��c6	
d�dlFV����K�$���j��sa�<<�`���
�2�߿�y�y\m���묤oŀ�2�'p��E�δ���tW����w�l䛈D,DR�d�p՞)%�s�*�z�1��ʔ�(ߑ>�Ռ�w��f�ÍP�P3���W��{�'�Hd&��Z��M/kT����	�r�i���;�	��\�%^r|u�`>��:��S��m�t��Y��M�ނ��-N�̈e�p�J���ʺ��,6���]�c�H�~��ˈ9�Ŧ��i��x�������2|nG��>�m�������I��R�yU�Z��X,����,慭�������wc�����v�����p������B��6ҥԎ}H��hS/(,r_Qn@d�玈21��^��:`���>0�0�<w�N|��?R>��?�T㕜��,ou�%����c�2��~k���nE�[����������!cb*���Y��&�)�W�&{=s���'W�^O;!u��jݛ�!V�V?���Ob��@ �Q�#H��l�Ö G[v�
�(�S���C�cf1��5ۍ��"L�g��'!c�x�5���d�*�������#U���!!��3�,k�P�gm7��Aa��<ҙsd���f�5��3S��X������>����)�6�"�
L}��'�񢆘vv�A�u"w�N��1��s��1눅�[��y��i�����C�b��Mi�aw�(��۟���D-�׍Ŝj`(����R�2���H���?������Atax����Gl`�;y!�)��Qѩ��(�dg�3��_�Hn��W���P����=�=�3�M���y���qZ�5���v(/޴�>{	M�q����ȫ�����3k�ϯ��ᄈ��.���[�^cE���Q�
��mI�ZKm��sy���f��,� �BO�"Ͽ۽�������� k�cx�^/f�����/�����h~�� � +��J��١�VX�2'(1/��%y�&{�J��NSV�G&T��v27��Эs�V@$x� �2�(p��ƞ�O$��I���ӄ�����	8ۣ��2��{pZu��W�9}6����86�e�dm�R\'bU4�u@TGVpJ�I$dK��0:c��_�㭔+��]�k��,XxW��7U�����ў�ފr�g�F��<+���#:o�J���:���1����-��!����������5��}攰1��=$��v�n3	���g����H�P�6��V��+�_h;s��ifC��)?��	�E6�	3葒I���ܲ��j��s�S�tX��ٞ�)�����@��I͇F�j�T�]O�ɐ948>�$l��.~S�Ѣ:�Ai�u�u��|N��$�/��:�j�#����.������|%9^�m�Lr�Ut��n���J~�8�`������^�.]��}�nXB�*�ք���s��ٲXpr+��1�C�9Q�������wԦM�'0�u��MB2�ߢ��1BZ����G��ʧ"@�2I�� \{�^P4s��C��s�����֭G��vǾj!�(��J��==?ozA-:���bc$�2$�6��.�@� ���Iw��5��kق	�uB�L@g"�P��t�����Q�e�,�j���S�����\(��?�@�#n�P7it=�ꓨK�������jt��]�q}�^#��g�*�9���(�`+�� �e�d����s���k�+�N�9�����QV�D?A��W�;0)�7�ξ��ƽ�pS)ILu�������(��α��� �[(��m�X3mK1'aΞ	F�d��w�s����)����� �興��W��*�Z�^�;,��$�'��[�Wi�  �J��	Ɲ�7Ҹ��ۋ����E�-��=y�
*N)��=�bD5Ɲ��[���������T~)���V��������Aߝ���CeyX�t1�'G���lg�>-��{�?d���*�c*�����Ys�v��F����
�;�b}P����	�4Pf�R��z���n��	���8����'��P�Ȧ���1+
mM��/Q_��������4 � ]Xb�N��	+�K���M>B���c��0��z0ؒ�o �؞¨Y�p��Z��Hwaf���*4*6G�/���/,�TEt�۾���7\0��7?Oښ��`�~ڳ0��1!^��YU�f�\�dEM��;����'��a+d���A��z��i��� ����؉3P׳���KV�������h�n �5��|n�65_�QURE#�oL�AH�&�|�j���i�Fg!��;7���0���Uݓ�M��0`	�� �)̺�z�cy��16�2(��a�QN��oa܇D�"
?/�{^..YRA�6�Ɇ'���H�C|&7�n�!l�.��}7�g0e�},����#XМ��u������iz�q�V}}d� ���ph��@����,#I2�b�rn�+X�����C�c�߯����^p�J�S�0���%e�:4���P�_s�lj|� �8qVqԝ�*W�ɛ�(/�B�C�M��g[YYn��3I#^Q�j��ܾ}��z��8jM�v��HY�D&�>��(���n�rU�[�律9/���K�X�  )WMd`�_e�"{��5�<Fc���#��v�[�O�m�k<^:j���ִOO劈�@FfB��ߖ�7r�˄d���μI�k���K��� ���D�m�$�yt�ځ/|*��^fb�U�o�n�y2��_���3cy�Ac�����,#���F���3
G�;�ʘ�#�|�j֠@���^�� �I��3�P�����0�R4�{��~�U9(Rǭ��h�;�s���ۂq�,�mQ9R/���x+���~��Hp�M���k��;�$u.ö�w�\:u�j���O5�2\��s�[��晬J����4Tq���)m:��V�@��n#l��^Z�cVh($tA��j��0��e>��=�8)��K�a]���/LeG�̵��V8&��4b��"D�X@��q�m:��Vyn�X������uL��i����#��v�S�A�$Y�͏��q�~�)�C�7��޻�^�.��4��v[NZ/V��W�o���Y�h�6���i��ެ��o獟����P'���ˤ��H�3��ӧ�����U���[��!x|� ŗ-��^�nb�N��# PY�y.�ë�,����&Bu��[D�(uR���e���Ճ�(V��B�ڂ���Rk�Xr3�u�.�1��D��9�Bݮ`\�0����4���`�Έ=f���ˣϽ1cq|M���&=�Q�T��#�߂<`�('��{.)M�7�p�����~_��0l@���Tc����7��l���Z2���L��$k(��"���2�ܭޥ��|25�N�_n-3�Q��*CpY�Z�9*J8X����-{�\�{����-/�z	��V?Q��H�c_�ǲl����K�8��Z*M�z��-�ɭ��s,Г�{������ѝ+�����b�Sոߏ�\A��ڪ##��+`?���z{f�!E`�*i������d����HbJ���P�1.'����o2���z�=l�ɉ���ͅ��*N���f9l;?�K� �w{Z����
;��\��%��4яG���X�G�.qm��S]��X
A��y��5�c0ź�T
v���zהUt	�0*��e_�I�ځ�h���s2�*�s�Ѫ+`�N�zd���ط�n3���8��5�W0/�q�hUw�����F���|w;���:].�Y���1CI�GSN�06����a��}��+�1�:5�˳\wgD��P�
�R��_��rS&=����[S0���z�]�)BZ��k�kD�@
A��Q���6,9��a��i�Bԇ���V1_ԇ&�do�I�3�v��K�8��mu�.�ͼ��{�� ��Ϙ1�3j�9�C�,�M�{���0-��H��郐��@���y#��AM�Kfd�|���޳Ր�
��8�yX�=~l���Uyz�}�sT�~��7�G�� ֐x9���`�D�oq�,M+����L�ݺ�����FA,��N�8�� +�4m�¢��,Fc�`Vz&��~�!2��[6�y�R��9��~�}�aƄ��и��f�i�r�r>����}	�zy.Č��!)�=�� �-��	Hgg�y�>-t��,#��q9t��ڢѴ7h�T���Sn��z��%�|�ѭ�{	{zD	n����
�F�`"ü�*���~��s�0���	�R���25> ]�v-���蚁)��ks�e���'hO�$�_h��[ļ�����o�b\��H4R�T���d�5U�F�IH�� �3�l	��ɉ���3����j\4��vU|)����/�4���!�����'�F�bSv ߝ��˞^IY��xQ~Hs웇R��r�͍��.�X8�����=�խ	YI~ �ŧ����NAP%�&����C����E��<攂�� Ő�':��=�_��P$�O+z!)�^���a2O��E�%򬇫�w�@��A�wݪ����O�K$?)w�	n[���O��$Y#9_�Ś>�e�
�íD�d%�O֬�NݳO	�N�$`������B\F��[϶h�"��2���2�,�}�]&��H���kh:|�@Η9m�������e����^