��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2���"WYj����i� �N�7A!�@<e�]N��?�jj�����W���a�q���#����MP�F�pdoF.8��+:���h1�ԭL��L��[j�1���߀/AP�0,r�F��x�N��>�RziB�M�\�P�ua��B�MɥBe�U�����v��+�R��|BC�:6u��8�B�����趟���*���I�lklry�.T����b��`����zF�v��o{�� ��)iE����[�Ix��L���0�𭇶�/2���e�P��;��D�f�
)2��du˷u�	��I�,���U6�d�#ǔ�.9�7��/�;�T�������5U�p���svl��o/3⧥�k8��4Ʋq�=y#��[/R�(�~�4D&v���^p�u,Z�1�O��&�ZmTgG|�,�
��>�1ݭ*`h������!/��tX=�6ϛ"�ق�̷��e1-� �`�������_��� p>��"n���4�^�����3�tGՎq�f��(.����R���E�<� 't�0�����B�F�
B�ڍw��������s $�ӭ�4��2��Qл��#�,���ٓ�A���(�Ly҈b`�b���W����ƅY����}G�<�'4 F�R�F)�X�NŲ+��6��1�iokGeP�� r��Hyp����d��{�������V�.��f4���4�� ܞJ|�b��J�öN��@�R�+/��t,yZ�&�h*ĉ�8�j��A!�?�?��߲4{�����w�8~��riS`yG|cׯ���)�ފ�F�m(��M�ة(��{\q�_�������C�g��b`�>?��p��D���8�((<��t�\"�#�rA��z׷�|��?+Q8w귕Aq���&�����d'��Q�raރ�v���b�,��R|)<�0"sF��Ic�3�b�ğ�W�%V01P}S���я��K^���r�1^	���Μ�= ��1���f�h����S�Q�M��k������6�;�>���C�@��f��L��\�󇀖6s��Y!�2�f��(_��(^�mgC�D}�`;���S�p5����լ��b�������)�t�}���T��9d_����$C��uw�p�^F:S�ԭخ���ʍQ��zhH���-(\0���YWcD6mO,��U>�2��dW<�b�:� B�Ȩ��&���)������d�
��M��|�^�dt��������'A�M�xK��)i���ʜ�Y�{�;�3��|H�H���İ�c����,Xm��d��́�8�o՞�?	W�A��.�G��9h�;Z��v�<4~��N����Xc�M5\M�gM���o�}g~G�7~�k0��<�ܯ4s��;�8���S�Z��B2Z9h�f�.�G �5�����+�q'R#9�݇H�޸qi4W�SQ�y>�D|�oըS��N�A�E�[�+	y���xM�<�>�\�V'U:�­���l�s���Ħ�IY"�P�����ǁNB�?����F��O�ÞA[cPALpۊ�F�,�d���+׫�N9� %& R�m��1!5~i-̮&ξ���YX(8����[#ܻ�F�kJi_�3�UtV�u��������2R#J׊]7
,������4A*�<���F~Z�������u���y.`V�7�P�~S�n��i*���I�Y;�6�Q�tK�͛bwvW3�v����XT�~[��).���ob�4���J��H�4n ���C� 3~w^D���5�nt�T���5a�-)2{7��s�-'L�_L^ -p��Z�T|�߻�"��"׸�CZ�g꺋e��&AO��-�!ї^���P�����]S��A�P���f�i蕮�^
O9Cj��@��#��X�i���`���NRcsĚG�
H��h�I��3^�گ;�l�*�O���((�����"�y������T0�	��
���@�.U������x��6�8r��K���!�dH��m'Id+J�H�Tci�����D^+��\�2��*@�ȶ�Z�D�<'S�LcR����w��xg�$\}��Pք�=����4-���5����&#C�����b�S�Q|^q��(��]� ���N�&�m����?�P0����8v2�E@Ɗ(��A8P�0.M�H�:^qz�����&;�j�҉��B��-"n?���3ci����x$"���QU��u�ʉ����)��DҺ��kK������������֮��J���.���q>����U�}����m+_�Z?�5r#��k��&��>��~-j�c�#j��E|�!ﯫ��j�-�o0��^N���dxB#mbO�L
���#lDC����ݗyAVe������ӑ�3i;�o4 �a72�N�Y�w��8n�F���q��mRY�MG�q�'��
2��Y��bPh�� Q�ɢ�}4SЅ�.��f��d�K_-P�Of`�f`���M4|�`0�=���	��iR?�g8ax�8��eު�B�b�p���M�A��x�bQ)�`�4gp1��ƺ��_��@�Ne�*H������xf��ןz����� �e���h�q	�N_`F�j�)N��5Ƒ
�Gis�/��Y�e�m#{��2ȩY�}�GLbŪ(�qh+��g�5r�W�t,J+��d��]]IJ��/���fI�Q��f7�e����a���g��^8ճ������F�7i����m��������H���>o�%�k��E�('O�b���?�Ĝ%���9Y<b�4U5%�� �v��z��hx�|�>.�<!,�D��e7�e�����H{Q�������G�6Xޝ^(��<*P�W��;��u�ht*IK�e��T����s���Hl�!�KN�ox?a���mR��/Q��%&�O嫞��o71�F�n��Gb�7p�q��=漳�{����r6d�56��TG��^�5�2���A��N�:��� `���/���y|��'�OH׼HB~� oS���,�a�����v�O9CjV�4���VaͲ���pc�%����QK����q��Z�u�O��0/|��S֋�� �,�2
j1-�������p @፨Ѷ��u�zο~�YSVF��Wa���'������y��<�B���ߞl��\�֦ -c��&s>���<�������?�q�dT�)1�����ߞ��c�V����`کǩ�2N�O��댓��|����J!w��e�
�`}�{|f�c��0�7nF�_��a�d�J�ȟk�2�}G�����Z�I��v�'�*�Rc��a�s�l(7�	�t(�� b_?ގ�h�X,�&��Ӂ�;����m����Q��[Q�A��x�^1s$��S�z��(� �V�0�kJ�Y%S���b�?�Z����["�L3��(a�X�H���x��Qb��(���1�;�)��XG��C�s�h�-�l���A���_,q=�yT�V�( �CL�00���[M��?z�Z��D��|��,c���&n��b8��DO�b��	���ٛ�������(b`'�6=�Eȭ��4��W���l��f�]ٓ�ZHh��yp�[�bl�1(���aȪ��L$��[+1�YI�4���Q0��͉��I��� RǶ@�rKiJj�Б������ڲ�2�<@Oِ���"~<y�������ޘx� 0�e|߿f��5vj��Bc��3�_��Rv!�e?�N1��vB��Gh�rM�����0a�e�@���<���`���'���:*0�w��$�(�����{�sT4�CM�~�$��� �͟h"$�6Y����Xª��;�S�n�[���Cy��6+�:rC��S՚��8pD��HP_�!���G���>=����~��=X��� �c#�S[�R��J��d���Ł�3��A����( ��.G<v��L9*^[���"2�o�\tb�TWp� �"����t2����,���5<@U_�Fl��WC�*/.]�nU,@d��}.T��5��M��D5��fv� b\�i�L�ZQ@�a����^Z"w���Ϊ��O:���i?�U����=�t���f,=|�R�;��@G�I�)�8�L�
�����%d>�g_�J���,�'=���Y�@C�knj��i*����Р�y�SF�9��sm�ф��A�����nr�@��߲y�{�/`"��u�%���9nb�#:�^�L�n��@.k3��z��(��r_w�{�4��z��ʪq¸jg&&���jz�lU)��7 ~�S�=6�~%�#I��^F���+P�c�5K�"i�d��.�����fS��b��n��$�;n����x����U��J���$���+�ɹ"���4[V�e,��!p/�(�|k�yC:Q�`Ӷ4���fw�ҕD����' �Z�U	�����bbtY���f]@�1p�|��|�9�zQT���a��q����\��܂ �Y͡讨:]zv��q�'eÇ��Ќ���8����%�_��Ծ)���	1�nyA�e���2P���ׅ��M�V]Fw�TB��c���,�h#��!��I������aI0�E+���n={�1u
�1z����0��B�U"2�%��WF }�ޖX��lI�(_.���Nr�U���%j<�`���IIV��̪f��w<R��\�����
�*sl�|����\�@P������¶��Gf�	�]Y��]�y��s�q�횰n�o�M���+�@�@��J�ط�����SLF�lV%��U���������oNq���i�5Yp���\<9���W�4�j|Q��p�Rv�K�e��աw�x��Rx��)�c��2"�V④M��.��`$6��#���^[���j��� ��,!KZ>7;���z�M�Gڌ��ЉQH�̍{�@�>�&�;)z��]��a�+4�!��@ul�����bo N�{�tz�#��(�I���zr��X%��crR3��c#�m�Y�ظ��؜� ��2��A�9k��
*�ҭ��B;ٟI���}�/��������߯��y-?n�E��a7��+����M(��>1�3Fv{#0��rا�4LV��r�:�[���^ �|wGŜ�4�ؤst��OSTj�v�M��%Qs�Ϝ2&X:�������ݚV4:=n��O�-�b�c2�`5��tL�$�
(�����*u���_��Z�N�G�ה92vv�å�?�|�*u���gSme��ڔ,1d*Ҭ��1f�Z�}x:���mo]0���M`"0_���V=��������𨲱�w~��z��K-W�f*�l�����&z�w)vjnc�VEDr.x�=�e;�S��q�wD�P����Хu��+�$n���w����X��R�%�a�,VGpt�`̅��~B������;iS�I�6��r��@*?z�_��0��8z��Lm�ְ�PI����K5�\WV�U��		��	��m�Ec֝��?ś�����:���#9'���"M�k������d�LG�k
�sR�5�E99��-�~�4��PS�f��Z��� �)Z���I檺��'����q����v���>
ٳ���i���NK߷��Q\�iI�.Ta�ՏqQQ�~�8��{�� ��ɧp*ȗ=8w�Vش6� 3�<�+)� ��T�h�M'���0�(}��:��r�	H�^D��MYj�pc �{�t����aߍ�[3\��;|]��s(U[��U�)}�u^I�����N�<t���yc�r1�`�5}���E;M��E����ˀ+�f��+�~�?7��m� �,��b^h~9}���Y������}?x�G]և�f�J�6�� *���@�G)����[d7�D�����.6--�����gOFd�5�T�$���	$<2���I�l�]���@X�;	\�*��끼@����(Q�s�>�c�mIR��Wy|�^�rZ��,���[��v��8�s��Ժ�#��V5�,����KmM��	T��k�ֳ�gǆ.��㶏?�^	�X�w�q��8P?x[��C2�?b��}����l6��|;h,�eK�,�-~~g'!!�̕J������_����u���}g��?&k&��hpZ��8� ��<m�ҝ�w\�k2��1B���r���H$(�Wik�N�E�w �+�)�4�� �_�H눔ֿ��%j��� �ʹ�$���˚F�ͨ�&�B)�N咅� ׉�pf��ݜl���b�cۤ�}j�d7�\D\�K�M��͒�-j� wp�|Pt�Ѽ�}ٹC��˱����_��;9J�5�-�S�Z�[x ?`���#A�.f�L�.�;�o�^����3�e��U���rF��z�`�"�#M���
LÜ��LO�q6X��>�x0Q7e�<<X����CK>���%��������7^܅Vh7Y��/.���
ʚJ��ϣ3B�A^l`��2��+�Y��~'�`��+�m7�.n2șE���N�4�������γ�O=
��av�On��6.�<�	�
���3�w
�m�^���m'
�m�\/3�>��2e-O�X�!���?�����m��L�簅@���� � ��F����IE$V�,�B|�5헄��\*tP\�)��T��~P/.���.��8�{#�ʚE���|��j�r�y�L�f����h�1*�i([�����>��~�����R��2��`��*�ҧ* I�*L_�z��@��}q���L*���֔�BS'{f%�yy����K�C�R������o��8� �����fi�:����c��a��S�_{�I-�qrp��<h^hv��|�`�m� �:j�s�HY(&������C�6���X[/��<�㧳�Z-��ߜ:M�u����|��g�P!�^H�>��F�~��$fS.�+v�U:�;����v��˴��IrC)k�9�MVM��=L�������yG��z��T�#.��B�Qf�L:W���ʕ"\�Nw��L������Z�B_3Qν��>�/R}�z}�K��q�7ws�������D�I�/��iYoHYYD��%몢(x�\��c�����0�7�ܑ�lN(q�Ԇъ�sO8���r>�E��?HͻUs؜G�څՑN�������2����m��ԩb?���=6��i_�ۮh\�H胸7��K�|�:�3�z�ŢJ0��Й��*mx�&��Ǽ�ɬ�
ԕ����$ C��Z8oz1&���>�n�օ�k+�uP���u�$'<)���9'\�D����F_nO� I��z�.��m�9_��nR�����!>��CA�<����v�m���KRܘ"�'DC�;8��5��㔽*��'ٽ/�= ���f?���U��-a�3>��~����ks��3g6EΒ�בO��0r�^N~�y��'�^K��O�`2�쾁�܂��z��g�!���If��E���tO�����@4�����f�'�����[��q�SP�	2�}�:Qg�
��H�Jf�*�C�����hb�:9ؑ����6�#��o�U�K�m�'x���ߖ���b_8̝�;��Ѧ-��]�\���[TY���7�.���/��c�$���c���c��]SKՊ�	+]��,��,���\s%���}g�3Tj4���H^�������
`�w�+t� ��j�7��\8����F��ԙ��*%�N�<r��9�-9�
�_�z��ě���s��$�(����� u���Ǐ�7�V��.��A�_�n�aQJ[ru��%L@��:��>Ӎ���������>/_��y ���H��qO� ��x���_$RlL��׻�䤳#c2�]�Ǔ�-��K��Ƥ�$�$�M-�5 ���s�)V�Ji�>�%�.�_��&�羠��ɪ��h��>t�n��]R���ddk������׭o�R!øc$U�yr�;��K�
)jO��!{�z��p��J��.��&�w9�ϠQ�]0~�v{dL��7b��[��4��pu^��B%���M��U�͗u/�l�P��Pq�!YO�C�=͛�O�Yf���ũ$��y�ĭ̟O��%�PS_�r��I�:�<��ӎ�n�9d|���=Պ��G�H2���g؍��9��V�d��!�*�.P�K��cc}�d�L R{
�g�i�@d��u��da2"2 �|=ĞH]&y�����,�ۅ�u�ꊠI���b{�a���:�����µv*�Q4D�F�S���r}Dӄ#�����q6�z�2���Z_��
�IU�r~��˨�z�,$��W��=c��Pd���!���P5�F�e$F·�ò8�*��3tC��Yzm#3o|����a����Ff�M���{u��/g��<5-]���u��l�~�%D�&�i�1;���tik�K,z��$#��)��,�D�1�Z=@���\U�W�	��Ј�ɪ>'~D��ָ}�<FO�ӣՇUxU8����[�9�dY��	��{J����dŪk�����*�F<�Pթ�Lɺ�R�t"a�� ?��/.���S�y�?bc�C��|Uo6ԧ��I�Z�l��13�|"��M)��L���aWԙ	;|��*��Z�"�����O�I+Nb�K:̦��42�w��97	���41�1.�p�^?!g"��#ܯ�L��^�a5� �3�j4�{��W�F����)�Qo1�t�_]���{��ʫ.F�>�����#�}�:�A�Ac4�2�k�ӜV4u�Vܴ�ap�D��b�7���<S�X����@�1��\�e3��}lv߭�|��H��X���Y�5��X9�/i*������!Aޙ<��EQ��N� ����K09\Ǥd=�������K�se���Bl���d�5��V A��iw�mT�����ҭL<AQ�ꆂ؅��W�-ä���Y4|A3C�v֭��ǸZ�qw΁���m���j�J��"�[
���Ɩ=�{K�`��dj�Ƨ��,�L--��QE���,�saȏm,�!���He|��b�� ��N2��򢠇�ޯb�KE��|�C
�À_�r0u���$裲Y�-g�t��ʔe\]�v�҂V'~Ÿ��E���sBS}eW��x�l�DųD�Oe����:�,��m��Yxd���>��u�O�����~�����K�t�OkܩEs��}M>Y~n8 �9�ԧP�J��ᒕQ����0�|uX��"޸HD��5|rPN��ԩέ *�!�����˹К&Sj�6q�k��y��*�$����)
,�A�˄ t(\M�0�Y��&K���\��-�:˚�
�W��9x�Ƶ9�%�[5]0 so�gf�
��b�/� ��D���gK�L��.>��`S�.��9���M:R��d$�'}C��'��Gɚc)yv������l����@���W,�P�Š�����:�t' ���4B�psf�*[9�b$������Y|L��H�Ix�V��H�x���L�� ��tIc�#qI)^�&���6|�O%��g�zA�����Z���D�o1Z�s�ٶ7���D�0�Vg���LE����W�3�7�Uֆ7`�����9���:U4��f�����#�Q�B����,Sc�#~bn�֒��p��t������D�D,u S_�Ų,�)��q�;/�Qk�XFש�嶀��H?�/���I3_}�d ����c�i_,�vt~A�5��q
��o�G݅�7�[ǥ����y�yd���!$nO�"?X2�Zr�Me�_�[��b�w��w�5�0��e�\L1��dK}��e�8l��7-�I,@%�E���ho+4����i�X��C��� Ш��x�ݜ�Ux� %G�1���ҟg��]2��W1G��;Q�|*e��|��N�{+LE���4t9��N8�UK��F��+!,WkG7��<[iD�*P�11�۹��Yݚw�?[����b�r�
�����k0W��n~z�4��\Z�KU����_i̟RV���{��\m�������[�ҡ����۲��zf�����龍Ѱ/�JkX�b�-���y���A˳~��R9��$��A:��P������J6.\�L־�\��FFU��B~�F��Ut��e-���!F��_y��|g����uu�`�r��]-hr�*�*�Ec�K�L�d>�2�r�C�3S�xs��ܯ�̴
�k����N�LW�?�Y��u��PB���%!�&\̩1o� �6oѳ:>:p�q�n�lUx�Z*)�~�S���s��Z�s�,ؒؿ^��#@mb:Sꡫ��Q���j��=ѱJ�xᚍ�ϱ���%U}�]��L�·*�@��yP�˂����MC����	e,���X.'Kg��Z�`�[�� p�ȣ<�	R�v{\w6b�A��W�`NR&�����1ЯC�
�=���~��B�=�} =T���;(�8h�,cït�l�!�%�IBP��[��@/p$܀}b�V�L@���E�A��[(3`
.�u|g�_��{�1��H����>��֥^��U;W}&�f�Z��iہ0��&�@C4�lw��H:�5�a��Z�jB��Kyx3ڃ=&�{KO���>�Q��� ����BG�d�Z14�5j�F���UG���s��b�t��[�;ӂ��N��CZ��(N/��r+���>��?�ޠ�lw�OA	�`��[#]vCi5��P�W�m�cG3�	�����"x��1,��)ƂS�y������L�N2�
�G+��m��P^�	)O�k�L��?�y�g6�KK{�v,a	���@�%�:���ؓ$Ay��#SYϡi�����{<٪�������Q��Єc�$/6�y�F���W���USE�^1`Ŋ��YTgr��!�2����o$5�D4�Myދ^=�w���
҉�mJbɆ�t�h��M��\䃓����`�`�A���i�R�	��c���q��n'���}Ȓ��.y�B��ݒ��������$YTL�XX��b�ץ�%BI�M�1ƞ򊻶�j!eN-,{���J�lB�U�\,�rϊvM�œ����D-�}y��$����cl�t�?�R`oHi��C&�Y��[,�Ĉ��,+�ƛڥJ��ʛl惉���LfǴ�$X�3�t��M:�é���M�+��v�7׈]����!��l��4Ӯ�-�Z%ك](Ń���GӋ�Z�o�S"JCO	g޽J$�mJ��ґ�H�USA.����D��.�a5	)�߾�OˁI�w�"E�p͕���_K�p���t�"D33��E�}�`�H��J�|o+.���r�<�[t�s��4'�.F�D�a�i�?�z�}��8D��`f�M��?w$+�������υ�r?�b:��B��e�ԵS�&���t	�9�?`V����:~�4���Pq$�m�Z7��wOimaZI��ڤ��'؈����%�ǯ���D4g��2�@!���!���Дe�ł��6���v�i�e��'�D���
2yA�O�U�:�l�y�WЅ3x(��C�L�ր�	��F�l�^^�_��'�<9�:�潦6V�>�~לzA}����io��7xpS��Ș�$]n����h�Awv�+��Gh���a�1�\��+��{2�Qhr~S�]xt���U�����=�!܇���d�v��TS���m���)i�J�*7��
�_G�c��p�fR��ɱƇ�( �Y�-�%%��:����[у�Ŋ7N3�[�-o��&�b�it������S���E��kTQ����j~m���F߮����@+�,�_�Gcu�<�M%��������z��˫c��g��[��C��ؠb���=L�ٷBNvf��O"x\�EJ�(�,b�Q���q�P�\rb��C��`*��
�]#�Ȣ2N~�x_�GTt6xw-h��\jZ��V�U7,ʟ�g�ku�c�k-�31ʀm(�ER	0���)�w����0���]���+���28e�sq�^R'9�Z������^Z����|��:|D�uX6�������m�����I,��"1�됨>����=mh��S1 -���)�d��Vx��W�Gpx!�|7�Th[��$)f)K�#{�ϩDN�R�	�ڽ���\Fʭ�D"�h_���^�5�1�F��Ja��`2� �u�1i��rW��u	WS�1�E;��M��8�ƨߵw\m��GL֦�4���3p���Z|��+��o�ÓY�q\�	:���*����pB5�y]0䲠v5�<1�:h���+��E�}Ό��^i�B�jGz��y�$�JIؿ7Q� l��{��WC� ���O���%G��Β��v_���)n��
�-�?�v�tC?>���f��ī@�b���c�������Nw�@}ow�pA���̰�7o�Ԥr�}k@��Zȼ?�7����q���m�r�60E�$��`(ʤ/w>wa�'ź��x�õbM4@6�+��-��޹D��f%Z5�tg/��u���oxۅ&�;�k�z��`�_QA�$�6���[����ػ�x�lc����J���:�H�6b���s�v��7�8Y���V�n��қKc0H)2|>{C�4A�>��.Oa��Y��=���X�.�`:�C���
�0�?_��jn�r�1�G� ��tX~�9ã�8�v��[�ض+�@����W�?d��$|&$�5���q��|J?�G�j����$�
��ý�þ���k�5f��y`��d��j�97�cV?=P���2��g�L*V��_�H��+��/?�T���'!�@���0�++ä[o��(�,<��9�/��iC�yN�D��Ҳ�cG����C��NW	 �[��9�!&	��B��p�Bf"�K��8D���g��bm=-���
�g%1n�*����<�(w./��`ql�)J;�x볌Z�� Ձ�r����� ���g��ܤ9I����q�9?��%4k����E�>��+w�%*��g!�7 Ҝ�j���i�Cfq��[�A��wm��wѐ�*3Z��P@~���([8�O� >����#����.��)���]塍
�~# ���<�0'�"cB����u:		�G�ly�]3�[E|�-q�-�e��$��UB�V+h��%�!��ۤU��o�
�l����^t���n��r�3�s ƪe�Ԅ�e��42&���W�]�(Ћ0ř��.�9v�e���l"���h���*� ���Z��sHn�y�~d�4It�J�"�p����	�V%dG!�P��znxF��_�R6�AЫ5����)�/1F��JF�sO��d�k� G=k=l�'	͵̷I�z�# Jʽ�0IU�8�aZ㰸s�m��v&��� ��]���.���'��,�O#/�/����	�^�e��<Mt�ќ)E�o�};4�׎=�R�)@�ĲJQ�|��&�4s%��;�XDM�P^��48q���<���'�(�0H�5���-:��B�->��k#c_��9{�Bx5-��Ln�Q�0/9I����FS�g�����.��Eh� �KN�&!�����ǉ03#ͯ3�|��&����g_�RQ��n4�Y�Su��M�(��.�jK���ӥ�U�e�d9 ���-p� ��B�z�*H�5��iF`?�9�3V��T�4O77y�H��l�߯�'��{ݚ���W�0l�'-v���Ԡ�w��!k��;�
�7�����
\N���$!7�ݐ��WHO�ԙ�bp�o�o�����Ԯ\�uP2���sz��B��@�yF�\%��oz>7�䧱p�%�X[��������6�G�����e�G��^���̝cJ��`�L�CՃ�GXԏ�O�}�8�V<xm��){A�\�榀���Vv���´TZ�y	�j�Űx$P�����Ih�*I���75ћ����\*�JȀj����@�rQ�/1=�Ǐ���r���On�O+Pٕ�?s��O5o�	B��ȯ���Fdˬ ��d}���(��4�Ş�ܿ#+�tVka?@��s��i󬿑��������/U!�1l^��#o���A�#܊ٌa�y�(^ʞ��w�a>�͏8��O���_�ټܯ�>�ϋ��]xc���q����B������Ӯ��㖎�(+&�]��4�B��=����Ǜ^,��|3�a"�Z�\�4dZ^$p/(�a�N����YZąGI(�*Vki�YY��iٌ�_,t#(� �}���|�F/�i������,ú8�ux���CR��a�蟻��L��o�록�Z��N�D>�q��-["�1�S`ҙȤ�R�
\f�	*��+; �������["��2V�gT���_?�}3���Z�J�L�(o��1��`��qۢYS�g�
U��%�\}i3���c�\23j#F����1H��"X����M��~�'��xO}
�Q�LQ��J�G?���!-��m.�Nz�VM�Se�����+g`��OD! y+�pu�,��2nC�Y�[⸨k1g��PK6l�Y���-�a��15?=`BU�~%+�W�f����A_h�h�%.σ{�,�%U�T�{���?�KL`��M������ �B�[��C[��B�ұ���#�mɃ3Uw����m�};D?�GC6�xLO69 �M!��.���������2�H1:���S��� �5���V����@C���>�
�����b8��栚���3�e���ɧ(�]쵡��Qe�0��.ɀ���&�P'��LOÏ�ƒЄ��VY9���k�&��:J����P q�(d������U ��f�jzT���:��͸�e54H��f��?l��g*ZQ^Ӕe��-ۿ�����>�Y�دʴ�{؂��S:=6�b�蟻f���	�M>8�1h9 ���po��PF�X0���'�9F!�N&>#�Rs!0�7����_�����D��rG�2GP"��pǩQ���.9e��!n�j7&0��iGN!���Ӫ;z�����L�wj�S�nsd�x�K曮ϋ�~A+�/oO��h���,�:���%��~"���.���lY	�)�7��אc�	���a�O&�u�I�	��*�[y�~S��r��+���yK�L�½b@�*�g�E�ғ3{�����౰E�o]E�q�K?���D���	Y����G}R҂�a�~���dt�d8>�8�8D�E;�U�f��JO>���l\?�.��Y�P �H�>y@�����>+U�P��;�󄳳7��Y�'c��V����yu�Ģ­�ӈ�?�
�D��_�D� �&�3A��(�(m���7�^ʾ2P�Y��yf[X����p��
f�<��a?��i�Y�f�&�#���!#D�Q+���tg�*��
c�ˈ��`�$�Q��s
�DL[	�Y��H�Ci�;�Q�OTk����P�tG� �E@oe��X��w}g��	U�h� ����Zु���JB�c ��q%�z���m��"�ַcL�o�v޽ъUvܘ{���� �Z����Jȋ��)$�d�p��d���m�.^���N�/�MO�?H��xU
���N�x܄���J��V�kUّg�E!�@�Uf���qc�WD�,R�@4-0���Z�UB�ǈb��<g�㗀Eq�i�w�5��O_�v�q��*>�� qQ�=SvO#9<��m�C#�k�EE� �_SF��K=]�<~��]ljő��=]l�34���l+�U4��U���Oz��D�*��ۤ�������v�/�'�[�T���n�j:�b��(�%�uŰ|UkϾh!�< /����	m�ČN-.�+� ��_a
FI���)��ږT����������N< �,��Miy�*i�n������,��bb�0`���x��߀�߂QC����Z$D��q�`�������A�����S#}{��@6"��3�KIP����7s5׷9v��G�e���r4"��G��/$�-}� 3����@O��A~/H�R� JG��p�d!��]'�\�S7��LO@K�PK����AP�EZKC���������:&tt�����O��>��#ԧ��oy2vN'd���&��MM�`쏙h�hbR>�\J?�J@���'�ڞ�ޢ�]�Ρ(O�˩w��i�U�5�޳�jj)�+WJ�d�A{�7�(Qz:.�z&"�5s�^�ۦFy.[tZs��:�{:k�{v�q�9���3�d����m�ZG�ױ�����r�Zm�M�Y�Y7��v��7��� 6 ߊ4,�xs@+GY����f��W46�fҷl�����#�C"^�k �z*a���≱Q
9k��j�;aqK�{��o%i�=�&LC�Ui�L�]歺��~�N��}`S21NY[�=}Ĩ�:(94^P*�q��5�A)BGY�����Y�*��d��c���ekף&;��/�&÷T��ep��=)�c������'�ㅡ{��|�m��(+0�*�7T�W�ﻠ��z�w���_`|�Bp�QH�Z�:��^�Z��
�fE"��������x}��)�k����^�(i�_�Zi�r�\��i>Q�tr��u��x|��-�X�
E�&�WK��>�9
�x_몰�r+9Fŕ�B���"Q^ޥjhBĭY��o����M�5�qNX�Qŭ;�0�Njna~�V���:O��5��n("���*��GX�s�$J��#���Z�7��J��(�d���^t䗛��J����{�1
�"|�Wu#��jjQ���x��j4��G�y���zc�E��o�G�[���
gw�m�ni��D5|o-�29@Vi�!m^�;��XE����#���2�W�<�;�����j���M�.��
�?�]U���8���M}ک�QYoZ�l�Y��q�/�>!1J�l�9p-DO@����#�k�+��n��yN���`�i���x��9>?T&ѳV �cE]N�2o��K��@�('�ad�\��iZH$�6�*Pw&+�^,i����s$\j�R����|�X۩
�B�� I$�(��Ϣ�޿�p����7� ��ڳ��e�Q�:���w?�=ړ:3
���L=��Y��W�>H��E�T��UX��%67������=�9�[۶	&n0.�< 0�'�$��m_K����)r]�ү�6�cb'���|��P n����������J<4�v�@o!� |![���n�v�����V�ǯ#�q��T����7a�M���X�BM��r���'�?�����m9�%��N4~�*��Ϫ�!DF �H)�����xm��R>�6�X��w�oN�a��?�}Y�v���u%�@i/B=�L��	(LH��%���@��z�}�?�f�+�J�z ��n�։��IU����e��g�j�2h"����C�`�v�&��O�E�m'��Wb�ia���=�~�{��8Kƭ�R�Z[Ӳ%����UJ}���j���$|̶�o�A���y#��= �B��p���z!VZhX�VF���k|�w S�8-A�S�l�Z�������-��(���b�ǟj�Ô� �=��l��S,��K9���:���y�B��+)���[&�O+MB=YX�S�H�]\�3�P~�q)�bn42O����ɫ!;���M�]jW����'G*:�u�w
*��v�m�<5�o�]��]F��@><U���h�Ǳd�,:��(�<��?ʹK���c�0}5�u��"r��鍚���
��C �n��r��C�劬}�n��2 �q^�s!'Ԝ��(�k���.�h�K0�n �����#�`I��ډ �b��u{ �&PD����}<M�.�Bw�ZX�pGf@iO��tf��@��j_�F%�z�FbE��R�$2�P�'��s�L���h�XC:z�]&�(��0�oM��[N���
$
8�9v:��},v��>���]���&n���� �^x	�^UB`������5|ْ�i�`:�:N��^6�hmaT��k{�n
�/bT�"^b�)�Aj��'�	�!�y��o�z`��ӧ��3����y��0~
7B"C����k���l���ڭ��74*��&|����pA�+m��* ��e�H`9�R"���0�m�7os�,r���B����|ÿ��t�h*���!�΍od��P��?4ڧ[1�Ќ8��PE*�,��th�d+t)�K�)NC�f�{�Z���)�U��P�� �.���Z�;�;t�M�=U�G�X�7�14��S��a{�Wra�C}�h%��
^F+ <�_
2��`&�	%�,���*�v�����b-��5���O�N�4꩓���_�����{��Vee�cƖ (�HYJYg��&?9䛶�k��I�/�cZk����p{�w*~�J���f���Uxbfw��Ȍ�8x�K�ּǔ�/���=&��h�q���s�|o֟_g # T%��ڈ�?��F���f�w's��sl-iK�x̨4���-y�����~|s��Q����N*r/}xÊZ��/�."\�K0�Z �P%\������ٻF.�gT jq���g�o�{~Ʌ��³����#E�nB����̱�c�Þ��dm��?{wo�6 �B���%���#Wۉ��=o���ς}$�1�6$�/4nL�**�@���������09�i�$�m$ݤ�`�O�d2�����?A�-9���Lj���Es.��[���F,���/b�	��_Tf��EHy�~0v�a!�&�v�I1z�hK�u�'=�Q�\aZ�B e���|�����I��)?L9����R�+sR���5{�>���!w��G��.@��H�8��l��� ��¶�x��������S��z�Ede�=N8G�K1ܲ�����ٴ�
W<�� gUR��m����K�\)/�@�{�z���I)�=-�
!U�I�0��b� @�`�JՔrc1����,j|�U?O�����.v�/O �|a1�7�ρ-���P��n�E�&�OP�^�^$s涕�.��]�����(��a`�R�8i5L�x:�x����k��"wC �kg+�;T=�8t@�ܪ|ok"1o]Vj/�=kκ��>i
�ZN2�?Lÿ`�U��
`���˶��f�-f��d�r6�g��R�����]-wF��Aa�&𕁂��u�k��^�c�?̓�ݪ�-Ƽ\�6�
y��e�EԻ�.�lHZ�s�����_���ٮ�X�Pa�m�Q��*ѷ�CC1�k��R�f�'�{�U���DG�E����@�p��Ԓ�_WωwjC;��|��A��%иe۞{fB�䅐x �d�"�j$\��F��Vz���+���-�ߗ�R����2X_0�\�<�6V�k���kq�ńY�*�|�#M��B��,���,��\�an��=wX5U�f����ݙ�ر�(�j?��9�?�f�fj����ң�+2��yYQ�b��T��t�dL�R���s����0���r#vj� �&D	��E^�޻��p�VI]D�O+��N����ȃ����:��8�4؜8���=��ugEA�D��V�Y�]s�@�P�ѯB�i]h�J2�_�yr�Dǃ��}��ƭ�X����Ȇ�V4��qύe!k� ���������@� �Iu��lU�؛���ge�ڳCR��Ō�Af�$��/@�^�>�p�����S����J�YUflckz�o��Uń9�\V�lx�.�Z���hD�m�y���we7_��%n�����Hz73}�w��	��	 ��.X�P�<�4�:8��Z�9�ٟ]�c8p�q%�߂J�M�g��j1��g���W�1�ѹ�������<�{��q��m���1�����T��_�1-��ex��wN������K�Y/hMe[D�5z#�֔�F�M�\e�J��3�	��^!����?�����b�d�>"�F�2�*}k�"�KD,��������䒣#lNۀ��c,%�p��|4������x�e����ޕ�E>x:Nf�����R>�������A���R_f�#qʩ6�J��O�qD"�^��}9=� d�)zC��&X��b�&����]��� +�㜛g�>f�v6��=�ܜ�Ȃ���"��ǎ)�e
���ı���7�s��2G)�4���r�"���ie&��3��¡�!�G�� ���=�p��Ӌ��@ʂB*�>��$^η��p��&�^k?V'�v�P�f@O�2�c_�Hg�!0��rt<���ʘ7��<�i�h�@�'��S��ڵyȷvx8��q
?�zL�oi�p���n��N�5��TA	�e%����7z�����m����P����O�,V<�%z1oR��F�ĝBܳ���o�ـ�V~�6.�����YQ�����NSF�L��8h�e��*�f?Ԑn��Q��(@ˊ��o�5V^��j�Ya�w��ך����8��
f�t��T�Z����,��t�2��:v�rƣ��˸�ZM���C�S;A��.:��۷&S�ʺU��o�}����3�vU)�tc�z���l{��H�rv��rbn9q�4�V��}[x����˱���NQo�ݹ��[�n!���!� �Z�f)�.4F���&�C�-�mW6B;�%fuK�}��?W.���Z̊����B�`&J��#�Oa�ʎ�?�3c�[B�I��m*%�1 ��pTl�'��k�1�*Ω~���.o��U�!t��6��uh�Tx].��N�,�b��/̷T��[9�%�.';2�k!�B�GJ��{��LM����LFX�W�YaC��&/*s)���{�*>8�ԡ�J���*>�m�W�̢Fq��W�W ��d*E4c�2���P��A3��q����G��r�_��ꕁ��(e�>���o:(	!�اI~�Tݿ��M��
h�~p�q����S@U9��'� ?�(����T��D���A��$v�PP�F�ӆ%�;�M���*wΩ�_���S�G��F�5��@ݪ�qef1�H���6zb{1ng����ԨI��mJ�y{̻�����IC�[����v�ˉ^n�M[�/Ȍ�E6JJ��ۡ\p8����M8C�s-靝�b��N����t:�SA/"�6�������8z�.s�	�E����`,�q��9����r��y^Al��8ǳ�*'>J���7i`˘b��� 7+��i���x��5_/���T«(���q.J�^�nι1~���x��>O�@R�xFTOw����B�;�%ro�Ɋ��k��a���J�8GJ��7���R�Z�M;��{���Ʌ�lU�!Fr���9'̅�X�fUA5N7���iA����j{PTq�� /��vZ�3K�����r1��ۙ9\F�o��
!	i�jݲo5�̌�?%=y>�q}��=��H�B��0�}{�CG�G'N�w����&�|\v��A_߿��U���5�d�f1�H=D���G��o�
��d��|^�zҡu�m�D�]�5��ǹ'�+ɇ����dm8��pQ�$Pr6�%¿{�rS٦Cc�f�;1���(���p�A�ya<crZ7��e�_�s�P�%������)��/l�|�9B�2ڑ�1�N7��DE���7Wo0��t�*�*�i�#�*�%1��B
����W���F���:tC�@ϳ�2��Q�Q�MTA7t�����,����ȧDF�|���4��� r�pO��e�p����$�S�'n�^2�T��u�Lq*F�pX7�Y��+)���0�W��plժ|����r"�[���v����?je���%1��ؚL�&؊�vk�����	P+�!�#"{�-%K�G�L�׳*���"�E��tѬ#�`��,4�'�,%�g���=T�Ow�P#-Z�otր��4bH:����9r��<�����F�Ʋb�#�>�G�a͵Ov��./Ό���oE�4CiU�=ay�{��Mn�E�S:�s����r/=�*[�ᰊ6uL���;��Q�n��4c;@&���c�e1����z���(�Y��~��AJ�'�*6��r�he��g'E�OAIa���?��Θ]���(vW�3%G��_q@�j�/5ݼa�,��u؉ѨI@n�ɚ;Sm��0:͏˔�?	�3O*�����n��%�T9��:tBb�݉��1u[��_<��-B�^��#�67J�w짾�uu1��yvW
���s��m���R#��a������HH�je�	���b{\T���>1�P ��tϹo@+�=l��
[��?�@�q�t�o��q�"V
�}1�,��~d��)"�[��7�%�tB��̣��~���{�*�6щQZ5�=�Nk�Mh����[b�@Bg�������tA�u��#��;n����@��x(���!�n`�?Qku��>�l�`�����$pĊQ�l���P ��Jݐ�0��=� �g�o�ꍴ8D����{>�SV�yW�Xw�c��q
u�m^�r�����Kq>�'ev���M-6,��t�te3�ŸR��W������[qb��-L�_��>�h8� 
e�NU�I:b��B�f~�o������3ѥb��`=��E8G�[$�n�d� ˷4�^,�� ��a���>�Y��E�P[R�ps���8c,�4t��*j�"O�20r�M;s�V{bG� ��4�.Y��8̳�0-|�_��Q"�v]֐E��9�J��F�� ��tq�����kE@ƺ�R�Iov�-v�����{����2t�mf�@��QH[񾧀W�^y�N�~w���zu4����t��Ĺ�!��{�ܭ1Z	�]G�F�����U'~�Ϯs=ҵ�܈��99w��D�/O�Ό]���j^2�҃�NvM4a��?w�f��3�WՆ�Z�`��L�9��gs�0�'��%��M��,�G��:����7�"d����$K/�"�M�A�Y��ѐD��3oF�>:c�V��Wn�o���<E��0���o�f�-x�+M��,\��(�~d-��E� 8_q$w
}Zv�Zz��i����j\C����V��D&�"��e��������?L˫F��㇫�e�"N[cd�ŏ-�����-��a>?rd�-Ag�i�`��E>���}҇#�H⻪*���1۴<��0�^���Yl�+�Yuf��6*�׮���ÑS�38څ��h���
~0+����1�TZjC��<"a�� '��c�1hÐ��"\?��_�r�������!���%�jo�^^Z���npz���b��1|b^��|l㿒��?���ə�!�qE�}���*-_�11�N[��hC?7��
srӒT��mť���2��D,RG�$hY�]�A�2貿;�)X4%J��z����M�j��ЕeŃS�E�4�[�<�g�&T�ԕ��`�2�O'Dg��X��]A!KNe�ygM��e�7��8����o��u�!/<c|�A����4����^�t+"�MB�W�?��Ku���}���[4���?���J�능�+ݚ�Ȅ�&z"*���\I��s1�D�NZZ'g���{zZ��0R|�0�}�H6Ît��-q��6�w$��HV��hU+_=���s�Q�l�����a�O��r,'�ʴ`ֱ����}/�Z�?����o���7�_g�q�E�ث7/M"�-у	�N��*}��=	�>�(U5m�L\.�G7�Kj�Ld�x�@�+O~�RÁm8��L�1� 
W��p�^�T�xf\��ڍ��ب��V8o��'�,������)>�SMx;е�;�@�Vo$�I�
'�:���ϴ��4J�6ݴc��g��ܣX���F�\��ϵ�S��=(��w�ŏ��������?HpG%��斉�w}�B#2�� �{R��@�*Ŭzu�;�y��Z>6i��Bf�m����@������\E�"7�v����1�Ȱ�Ӳ�Kۜ ���!���w�J.-�Bۛ�~������u��ܕ6�5�`��p��?ש�t����=$Zd����4��ZTI�����O3��A4h%���(��%Qt~��n�J��ċ�#��R��ir-kX⫱�`j%�hZ%1�y��q�Zʃk$�;Hq�E79�80t۱#>cei�����R$k���i�� K�K��4�~�	@̤�	�OS1掵�D�S5^�I:�|eEh9:5���1�CXTu�B�� �)(n/?TI�Q>�c"W�e����ў~w3���cE� 5/``�3hտ!�3@)1uy�A��v��p߻Ӏ��o������S�Fm���Y6�O�����z�Ɖ����-7[�^���O��ٮ_�EI�z�7
��.��D��W�f�̶��7G�Ms��?A���C1vv�lD�K�B>i9�̛�Ƅ@�F�=7���׼�x:�M�D݅�|A�����n穟I�V�gF��[iT[J~!\�e��>;�����E�1���è�n��YU�h>V<���1��c���%*gzឩMS�}6"!�����v�'*��Ḁ��N>�r�U�vVl&m�r���	/�R�k��L���f��<ށr����A���7�)"d�۾t	�ƔR�g:R�8�ڭ�-�=!���ք�B�_��Ҁt�C҅�|���!q^��=zE���J���H_dzD,���/�n�������x�a<#�e�I�Q[��PQ�,ѾȽ�|��Lw����:��#Û1<�jc�)�@g|m�F�8;���Y�Z����W��ň� �lN�r:���{���5�ʅ�l4���HE����=�\�Iv�<�ΛRdmŹT��2�m��ذ(�Җ������ �앿5��85�?"35`���2���&ě�{ol�:�*�5�b��݈��ti�T�!Qț�= �=q���?($2�@�P�5�a�8����b�y�܊�y�%��^M6޸�L�	����z��bt���{�����K�f:��0E^��@���iU$C��^Rgp�q1��:F&xc`j��b���(�,�R���E�D�$(�V�ܴpt��d���E���b@DH�(��ej�rE�tT�힊��id�������p�֖l&`�Fty���D���=����0�����28���4�^P�IEW�!,ptW��ŵ�&�����{��^Ŧw V�t��1��ܰ�!���9A�Lf4��������âr7��c��Mu�RHս/��N�c���ð��!�:"��޶�&�ɍ_�
0�V;����=�u�K�������}�F�ya�{"=�G�ރ��%{-��ʹ~�%X-��n�]�(��S<Έ�֬kN�gP)m��o��v�к.+�"�'#�?�5C�i��>�]��f+Z.q��ӝH������2%],�4�����Ѯ���|����AF��7q���Rdj<�g���e��ZK[)o����Tq$	��4�$�����vQ�_��'��/ʒ�����m��i�� q��ui�Mi�V��>��i��|M��R+f���v�9�];y�S]�b�;�Y�&���'��L�a��o=��������q��Ӳd��fsO�sn��hu`1P�l�&)�J��a,�mz�� ��ٿ0k����vY��3����#��R�[D��Kd�c�2��><ce�hY4�'h�2����U�g��Z��_e֣�@�n�HbRYɊ�Y,�j(1���l��~�	�4)�o5��N�K�$�YTb� /۷Jm���p%��,v)�-|Ս(q��]_�2��h�"0[>&l)��Hs~a�*T���}5�~��`��ס�k��]I�z@N*Vøv����]ꕝ���rYE,T�cI4���C��>)�B(���g�;�]ȻI�Ww�
���7��E���I���y�q߉��tMϰVƥ���V%i	��JeI���Ӛ}� xx�A!����x�͎nD�+:�jk��K���*cF"ir�����Q�W����da`y�ėa��̬㜣x�e�Ic!�֣z��Y(R&:e�4���톛9Q����L��*褿���!�3����RS�>i�Ӛe~�X���8�-�� ����}�93+�Й��O$3t)�_��N�Uk���K#�["���dar�i��	ԯl@u��u~���-L�:.���s�/�j�%�р�[I.s="���1�*��-��9"o$X^�Jur�mGvQp93L�Je��/�(�8�|�B���Yj���1�L\pd[J�@���!b/���������*���w�d�u�R�2e3��z���1=���ې���xS��� �_`��ğ����E����=�������,'c����sa#�N���9K�I7��`s�N��#�X�.�Y����%s����W�7qz�w�h�cC��a)�i��azM��NĨ��# �$���
����p����6�.��]~�*�w�?no��Hθ��H(�A%�N*5^f���<����d�^��w|�#����}6^H�3a�m�
�KA�j�rB%mI��l�U�cT똚�x�n�3��{��y�'�bR��Y��|2Ji�V{ǥ�#F�C}����7J�$T�����s��ǀ�w')!S��uYT-�c>�1m\Ϝ�\X¿��BY�8����,�|7'*�~P���P��.�*���q��󺧢�@��%�z�&{p�Fϔ���P�3t}����`2�̦�.3�'��ПQ�����:).����K�];7�y��,GC�V��6�v_���}�=�:�n/�Ma�T"�
+e�9�����OI���׸m-�:L%"��O���Ww?[�J-��ӥ3J�M�ϼ�����+AҒ� c�ub3�H�!r�Z�3VN܄x��+��A.�w��b���x\GǼ���>թi}�Pԫ�j���pa6O¼L0_����-��������d꒽h��iE��D�ƈ"H4��1�����YK+�j�k��S<� .3��v OqM��&�{�b�G��+}
�f�t'���P�-��PG}%p.7y>� �<1����Q[�ap�iL& ��,z.,h��H���;�l)��aZ�R����1�?�\>K��DQ�?6*��8�[7M�e��S��7j;�j4��G�T�E`�wB�\�N���vQpӾ|�V�$�*]Y��Cr�4�QlVrn{˥�Fd����G���`�Ũ�89��8���@����yp^��:+GF�g&�y:zU�#�a�w����F���E=Q�kK�w��ԡ�x����%���,X���a����B�P}���l	.���U<Z~��*1�XR�$�a�����:�B���$���ܢ�:���Vwl^���K�L.��_�w��B���`]}�xR�Χ����;G�(����������k��i�7�am�\�9m���캄e��N7��}�)�R�R{�(��vd'�!�o4�!M7�J��Щ?F{e��hl��u����j�&%����R�^%S�DG��'b<��J�4���'�,X�'�xG���)���p��V��Jb�X�m�P��%��W��|]�9����xr(�6:,�EC��F�׌
��+Cӊ���f>�$�	
(�Bv��=錱㽠�1�a�aE����M��yJ%d|��`��S��`��4r=ΔeX�S^�J2�2�M��Z4��1[^�jٴۿ�#
�b��万����w	C4�6lB��B�&�u�����Ym�l��w��z���@f~���WG����&Y3�)���ۄ�J�����٘hs+�H׳��sܦ�����"���!�X&z��3�q�x=�S�m���_�;�ix$"
�pH����]���%�^�[�-4_��������M�!�4a��t4��K��
����3��Z�%+
�
ظ�\�`M�6���3G��Mɖ�sD�2���o
����ŐTn��,�Hr���yI[��,�Fli�+
w���8�1�J�;���ͶY����*ar��D��`x?+b>��~�&0���!,�g�
���R�9�w��~��7�y�!��Y*ubؕ��tc��ܹ-&��9j�;�&�%K/�� "j�ٙ.}� \r%�S�'�p��35`P6u����M�ЗW�A�Ȩ�d!�k�'E�Dgn/����ʠ�����3AD����Y�H.�{�
iٷX28�ݛ\�\�Ǭ��j�sy�j�)x=N��̾�B���p�Ͼ�=�^�O9��g)���������&�Lֵ��I�@�:��9�
e.�9�Y��Z�?���O��8r��$O5����2����*�#��
�#>�6�Bs[dD~ O9pA��ރa���9�}���{�a��� |q��Y���Z�")g=-���FK���~����M&,�M�2ij�6��_��A�M��~���
�³WI%q�����I�O�=�;Fۣ���I�E���i���{��:^��?p�Ł�	��߃�V�m��61��o�ˢȧ&�Rsr���g��1�D�Y� 5�=GƁ"L�"�*�'j�05��A�l�KИ�G�\�-����#�1�x��3���4yMݒp,K�b�Չg�.����e�禄)�8GI-�����d�z>�� ��TAK�!u���^��o�O"8Oǐ�Y�HcpzPRb^M�nn�"