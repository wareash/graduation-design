��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV�@�fP�'�8�p���G�<3��������/h����a���7�&��7(SK�Jm��?o�w��0�끘���+GJە�	؟�Փ/��IY�]���1Q�(�H�`|"��{�!R;!�PP�G����3���>l�vr`�i�|���iU1{>x�п5���헚h-����dm�� �C�W������7W9���m9{{��vI��r|�f�������W-ǉ��37�P���5���Jåا{�\�u�?߷�dn@6�zf��r������;�amb����Mt�w^J*l|�G>��@Ȣ[/]�Z��i��������.��m���#W�q���46�<��@�S̪�EIE�������n�᠉��g�1yp��.?2�K�W���N�B{<���XO.�w7Yڲ;�H��\&�]���.��x���]T/q1��o��p�-Eӱl��b�ZOz�"3�%�O ���{�/V��Z,���(��¢�DGs��7[�/j�"�bUÎҹ� 頖��A��~��E�|F��"�������>��R��b#3-$4���,��H�\��B�7oڒ�?Х�>�>��:�A5.��Q��C&{�~hF��dߌ�<@���=�,��j�E��3U��6XӎV�m�ZK���¯8�[���)xF���s�ln#лy���P�������6әh��Z�2;yo��>R�~\�i���8��g��$T(��*�z��H֤�"�פ��5�i���#��s���ċ����R��kb�O�?�A�'�"�`kV��Y�ֵ����|��xU�����E���]	�\|uz���H��r�9�a/��E])�e *�ʓ��e�H&����C�zƦ�B�6K@�(��@�ֻh��6 	���b�Y��R���?p��1{�8��3A��0���&[��"F_h�ͺ��cy�$&H�7ȫ큲F4�>��b�J��b��^�f���6 ��P�z���C9ޚL.<k[ �*]��0���$[#U�����zƤX_����Ā�l��&��(�y3��k������;�'o�m!�P�hP;���~�}\[[����; �w,�rO�n�n_�r��u��^�S��1���z\gZ:W���G��`2�f�S"B�d�'h���.��^I�[�U��w�K5:��Y�,ݚ5�MQ���0%��(8x�@�co�������K����k��S��߰ڠ��	'�������ɺ���/��P��wB�^�j�����(pܧ��m�^iL����L�A��<�"t�^	��U�&���ܴ��-��t�d��a����+8�]`s�䞠��.p�܄�8	��������GHupjf��29��^ڮ��B �����3�����F�C�{�e�Q�cF�_6�X�$��+[���e1U��-��As����l"�$��_���C|�����Ei�ɐ�<�X�������K\�f>�;�yl��a*�.���M�mz��v�!��)��"E|V�U�>R�|���hӰ�nk���lԕ4w�BZ��;H|��Qw��5-I0��jő��.=�WjYs G�����x̵&%�,I7�Y-�h:�Ϊ�6���y�v���AJ�Eu��Wtz�q��+ �H_#�5 � p6]G ��z�a���~~���҈?�N��A�C\��}']��(tYF�
 �jW��<��!�'�Z�^
�^���#�� �eĖ%Y���0��ȼ�r~����"j�X�2�!Fև��hQ�b�����N��$FB�����M"gn�"� �����@��ʕ���X��|G���zFHN�S�ǰ���]�*ɚ� ��y���t����^.�ŧ6Kf{���n̥���8����G�D�'���,-�!�^?�?�׷�Ź�fZ4I�$j25ʹ�b&_t��If^�|�Mi���Y��z��@�5U�x�^�s~�	�E�JOC� �1Qf!| T,�*6��Y�Hg���T Sۋ�/�`�^���~Ry��;��KƎ�rx���f܏Q�aa`��s>����8�,}�3����G���	��v0�[B��"��1/ix6���X,�F��IT���:�˫|'H���7YK"�8���4M@�����)Ϙ��]��_�$���$}����y�]*C���� x(ݗ�nmSA%��ϺW��h	7�PVꊤ��,4hb[�sAV#��~!�e��G�V� ��o���}��jձe��@����'��L��D DUg�Q��jƴ<�ط���	��%�J:�[�`�؉�-NP���P�tt�ʷ8�gY}�&��h^�����v^}�U��Eں��ᅀ��g�y@m9�����,�����`�/�ޣ���%
zfb�Xy��Z�GE����4a���=�/�����vm���hC"�*�O/���tpm�7�Y?TM�/]u���=U&���M4Q�3P�JG#G�?㌤�3C��^�Q,¯��eL�4�e��ZU�g�F�_f�t�@s��7����R���U��nGT�m1�
�����x'�ITx��Ir�Xo�z>	�ǰ�b�5%Sܱ&79���x>>���#�	q�!er�J��F�3|���VP3`�3ĲdlezQ5(<e�ь���:�<zJ
P7| �1_{�����s�*��i{��eK]2�9��{���a��f��l�o��3�0�п�"��/E��s���_<|.�V����ΗL�h����4�#���%w�r*�;���i��Ÿ�`�N4V�o���7��h�]�W�҇K�(26���D-{vM�Jʤ*��5�L>��p��Q����.�)2�^i_.��������sGU������x�@l%�?��zI{��q�����M�-�Ex������Pdr��l�o�\�����'MA��B"���M@��6�&�Fan��A7��U�)(�.x����J�~��ϧ����%Dl���Ă_٦����!���#8R�T���v�`���-��^��\� �{�4cGXĠ�ƭy�$��kB��SD壞+��"R6v�L�-^�s�N�]�^��d39��o�����N�+�[�<���j��:,��U��_�����	��iQ'��d��xS�I���F8�0�O��p�}�&�[a�ȥ%i��>lۈ{l�/��r4	i�ZI�ix�@وDu��wO�_s!���7%���Kd�W�B�a��sS�ڞG2��l�����q]����c�N7?��;-ý�L�)��)��o	�wu�@|�Sn�S��a-���Å����1;�B
ݜ���Q��)k+2�ٯ���2�U�a�Ζ3�dZׅ�OeQof� �FBe,���m�`f�4���q�)E~�83L��e�rxo�:�. ��s�M�3��C�
0u��Ҿ��J�x��-f`>Y���O���0���,����A{|!
�y�><�˳���M�R�>
FU���[�}S���!�f	�;�5�>�f�ڲ�Q
��yWUwh.�����׆���T�ں���H�N��
��38-[][J����ǟ���Fg�K{R�����9���MT��CŘG�>c����멸1ޗ�='���M�i�O7���rd�ַ�h�\�b�C��3K�i�xh����f"�Nf�{5uQ�D~���/'L����O��Q����f��0�������
Vc�n�GG�Op8k�n�e0��b|��ǚ�U�-%��N�i^�D�R�<�_Qݙ�*D�p��������/����t@�>z���<��a�ZՕК�;��Q�4�(1�'�����}�7�6(��v&?�<V܃|�)|@ȨpC@�5{�Q�;d,�y��2�D�M�	�p�F}Fp�w�ʰu;�Y��ژy��≭y9��W�Վlk]��0�"A0рlr>��!V��s̗��U��_ѱ|�)6��հ��НX�"��S�|�\�:�9F�tg�w5�\2-��Q��IP|�\�lc{��JŬ؟mR/��r�XR3�Q���?��n���d^�B90P�*�-��lL:j�>���]�w�	o�Jo���b�^���z,& ��f��~�:}7J�h�s���� Cx���P��E�^�OQ��;�x1h=����� ]���q̼p�)�ƹV,<W䒀�Z�J9m���]�
B��[���r��S��Dv��FI�[G�zgX�ia�9�6���s��^_=�C��wv��,�#u{`'	�+>�J�J���inލ�]&GB�69���!82A��Ԛ�]$w��,�}]B~���eI�7�vJ���}��[azġ�b {Ō��K=�L�� 	�������of��{IK!&R���`wՐ��E:��?�!�Ď�j��7�����k��0����������㨌y����D����Nn��,#X�vd���p� ��y<�@�t���t�ܞ�["H����i�N
�ez�z9T�}N8�P�阱z�D�Pظ�;�����]��h��Z�y��N��~�	S͊����ܭb�;���&�ib�#r�Ӕ����Cn?���^{8A%,=̌˟�]"�>�l"ڎO<҃�a���=JP�]fL�4��֞�(�l����рٔߍ��UfVr�� /����QCn�3s���d3�Q\:qG-�n���7��1�hE��b�|�ɲ|����"$���?//~�CsZ崍���<� ��>ly�d� ӑ���X.��O��t,�K*���L���=������"�@��2ZDkqBv�4['�_4g���6�㪭��� F�C�Xy(��,Ô�W�V=_�i��u�D�͟4E����tr��5�>�<S������+MtK}X���qP��ԍe� �#g)gbJ�IP�=ce��v[^{�O(��+N�sW�	O�F��-���:����h����_;��궚�ĵ����WCA����2�Kt�/�{#��G[�I(�@�5K!n]��i��ٮ�IMF-\!��I�ƭ�^��	�R7ǄV�P�/�8�
�"p���񱂕��.)F�Q��H��,�:�n��u�"s��0����Ȣ�(� �n
���Y02j0�G�Z�x���s0ԍ��P����!p�ѿT r�iʶ4�X�x����"c��dj�H՗F$���c��54��_C�J��K�㦅{Vg<E���ܰ[�s���q�_�F��EW^�,7fq:
�\��n��Z�w	��ٍ���A�1L�rn%~�a�%�֘5� t)?��-��4��9ፄ^�+��*?-4�_���i��/�_���Ԅb%�A�LBP�r0�-�gsuĞΧ��x'�v�בX�����"�G��[��G�O�j������L�8$j�azS�$eòo���Ά7��X��ɦ�c�2N٦O�;<�7�xj�OA��������N�RF��,���ˊ��KN_C(<�C�-���QG�A}£Ɣ�b�Kh0������b!*R-)�6�?2���S7���P:D�Ѽ�cל!DU9,����=p�9�.�f[.���W��<<����b>��dzUK���/��O3����6���Ϩ��y7ܷIW�x�&w���c�hM�?\ Q� 8�s��k�`�za��:�Xpu�m�F��*���BM
g�JO����ֿ	��^1B������z�C	[��N���٬-I�E��n��Z�P�����e���\	���;��dt���hj*��K�~��ѭ7�/z������P���,�T�9|E��� �I�`�Pq2��/�eþd���&A0��q���D���_�#3_�j�HT���qf���wX߼T�����yc�b	>���u�|���%u�T?��Y��핹�����m���Fxrd���`)ʗ�@%|b��6';�A�{��{H��a���7��<%h���¶�{���n��6hh��ƽD�}D�`mQR�Á"����/^G��%c)�F� ;�s�Zi�8�N����H>n$�����,	�CУ<�L�uW��͕8�N�ų�9�����N��l��� E���q@���(�	�/t�/�z�*q��py��J_'��B8�R6�[?�����̬v@�t��a8��m�s]����M۬.���"���̭}�"țg
ɬAea���6 ��S��۹�#OȻ�����E.4"w��%Gk��wF�H���Q	��⏼]c/|��/� �"A���A��<�������:���h��X�s.��4��|g���L�0���8&�#$bjD@�<mu�_���ܣ�6�Ll�[�^�+�xU话Q%~���O�U��(o��bl�:c
[v�l��D~<l��ŏf!Yԋ-0y"��쇭
'g%���dD�&2`�J�iY�fZ�ك�|����WZ�a��A͹m��J��HAf�Ʃ�B%#�b�2-dʤ�R�G �YX�,��npt�,XY�QҾ��25*��CPN��w"�;�_9O� k�p�S�W$I�tY#��Ke��}签�t+</v��/y�z��R��#�������p�������m+Ҫ0�@��M�I�הƀ/��$<����׍e%��'�L�L�Fѓ���0 �����%�{�!�y�����k�U��l5�n�J!�8��I%��.f�ܥ�N�Mʱf��[��V@�9��@�q{O�ABM�W.kG�0p���(�%�3�v\�8+������R%X���y�.2�	6���s%cp�C���e-C���xhbX�o~���&Y���`6�0�~=/:��o�?]b?Y��EOB��A8���u8Lx�������x@���;�l�o�>m.hP����
+C�،�Ml��K��0o�"3�~�mu8)��Z'NQ0d%S:�dU���ő"�[(�vs0����T�4I�	]8����[��|/mdDp��a-��D�`np�$�3������7B�db` �v����Λ��1�UP����(&�KB��p�t��֋7,�EG^�f����\y2��`��.�ej��D���m�>�䈛G˦��큐i����h ��������F��� Ї�H��,FW�.��o�����c~��n����UWq8łɶR��y�a[q4�إz���#�:�J1�
�]vN�y]ؓ�w%�`R�}	�*Cz�Rw�>�,�ǧq�1Sr���l��p�%g�KS�$��S� �'�E�jx�m��i����P��۸%�)Q��� �&��ƃ��B�5G��h1�H���z7�z��ŔQ�bB˟ꭐ4傩�^�٧�i�x%�.����Y��v��ٜ���:+
�ժ������]F���)�\`��F� �}�A���P<b�`
u�(���o���p����OC��-2:�����?S�dxv����I&y�늳�O��7c�'�^s�wP<�j�ڱX�QJ�LD�Jx,A�/��G���*��+�"�6
N/=�G�䠰�Āe���H1��@�A����|�J0f\����J,_���0[{�W0VOM��D�tH%�1�D5�v��جq{�p���ܥ0��K� }�3���!��8o��g���Z�9�'LE�$�,T��ĩm!��͏�6mtR�����պ�;oKST�㥶Y�+���Bi"@�7�r�#��):yۆ/�0�^9���(��u��ٯЖ�d�sl�٫�,����z٧0T7μۛ��	r��S7E�����+��u��)���_�I�mcI2���@ʃT�x����m��n��WQ��?��4秜 W��y��l���r ٖ�+>��&w��j�:Kx��|js��Mi'��i�+k"���O*�c~!���6z��&�(�/E�O�4~��2�U_ ԕi��H���y���J��X�R_���ԁ���I8�YF�x��7g�,
�t:A��Tȍ~�lr�zE1��.?EID�:c^�a(	��H�6���b' �/ns���vZ9��w���'bح"SD�3�ĵ�쒗ih�_�M��H}O�,�W��8rA�!��¨����]?6!>N^L����S� �{�o?�>:2/j������%�}5X6����-�c��8��8Ke��:�D�f�(�vf l�H@J~N�1�]� ^%B��h��UQ���w�!:,#���]P&N�A�ؕ�r+�����1��dʉ�H]��[/c�c=s�:u�[s4��$tݞ J��<�oOI���,T-=���Yk����� }WM�^�'���[qDQ�5�ŸЃ�T���J~��-�'|���
��֢���=�"j���o
�h;dS��ݮ��P�R���G,��������IS%%5=a/��<�K Uո@js�	��[I��t���qOS�SΝ���A���!q���q:����u��X��@�p�@�B��Ջ4��{肮ka}U�F`�Z�mG��T�b��F�k�~A �]ӊlK��X9UR���l��w�?6<]�����f�{�am/|�����pt�R)�� ���}��1;��1ۄ*2'ǣ���Kة����i�j�h����O�s���H�T�c,�a��ᦹ�����,-^�s������"�?ӗ#���=�s4�H��Ó@��fyk\z��#7�Y��/.g��OF��91$Mn�b���&�E�m��
��m�`�R5S�4�N4�%#/>�cy��)3�k�ij/�pױ n�Z
c���T����h$�s4J�@y��j��V0ھ�pPf�>w=~4��U�N�뒮b�\ �>�s�No)h鑰��N���'*�	�4�5vrY!t2UA$'��%��E)����æ��F ז��hx:�ݻt�j��UD��_�?y��3�<�B�B�+��`�b���a;8���lt;��S�c�C%����Ҍ�m�	#E e�p�/�ʧ4�Ѵ��6m��{:���}=Ki�ak���͂V׶��Y`�L�8�N.^t�Y	��u'R�z��w�����xk�|��bL%\�s-��5S�z+%@_��5*���6�z2����㳟	ED6��	�����gy���"����'3�� �"��2	�<������vdm]$�����/}��>AGٿR���fH�}B*���P�(v���֌�S�w�	�"����Y�m9%��w����e�{9H�]�G2������ze`�G�g�R����N��?�^����K������
|��t�2���U�/��������ΪΉ���(�m�~�3�� ����fK�Bۙ��K*��&��xUU�Af�j�Ɨ�/�9��3��������Ψ�=��IW�u���0W�`�^U�UO��O�������Ux�]OX��
�q��J���N�����m��5Trh�x�^/4�~��C��,`I[̋wW�8�K�o�|�	�
@�a��7��PWcսq-�K��	�>數��>mg�Wx�1+�^��ԕ�%�Q����wC���P�f���Ȑ��8��#�W�mǻ�a�y���*�2s/�p&�{��3����6�������ך:oT����,��)�w���rSfc̢���.SͿK����j�^��O��<�f���~i��USC�x��t��k*�B�7���<��I��}R!]���S�q0�87 �ѲOtn�u�x�I�\����^z ��5v�<�:��՘�UJ�����+Ja �w�Z,���ܧmzV�I��k�zD����9*��a���h䴲GC��e�y�-e��!�ӛ�y���h�ƞ�C�AZ���5R���:�FXI� 7ƛ�_���5�������ۺζ/Sx�:T�R�Ҭ:{Q/o�_4��YF��K�@,�LM55�%� �W�d��zE�g�gs}L�v-pD	p����~a�WZ���(`�5x*�6�╁���G���W�z_�$?�A��i�.kZ9��<�̏�?/Z�׹�T���6����k
���`� J�[����^����0��'��D�qJH0��h�It��#M�, �����'�����9LM�|b}��n��ȁ&���&	 -��_tx\� �歵��8�����/�W$��w#f��@��4�WS�ƴ��K��N�wT��������Ȍ��gI;o�{<YQ ��-��x��-㥑�&WnG.`l��+�½Ή]c5��ϕêS�  H�*#��9��s������%D��5@kҡS�:�:Y��I�a�5m���O���r��~/[8���1��m��ԅ;h
��"U��"�Q��9]F��0�B���!�f�CIR����V��p��}1��������A�I��t#5 ��r��R)i��e�=A�հ�g��e㼱����U����F�w����C�:��[�Gr�/os�יp�!s�
���i�j����rI#�@�=1�R�y[i��X^b
��B�/���i+��Z�ZQ)��U E�,�����	h&�ǝ�� �ҫ�=(~��k�+�Q�v��UΣ�+I�;4�-I��:l/U�4>�s�%�o��C��.�m ���Wc��߻�&>��n:+��I���F�O�
����;�A���AE��y��ä���y��C�K��F��0�D�;1>�:YG��J�t|:�>$Ƨ���;�!�5�*��p�`�А��""i�8\K�V�,6��ӯ�c>&�
.�Ҙ�Z�e&�x<�	��Jw���������[�Q�S(�͠����Z�������'�����]���1�Xǣ� E���<���R^���1/k�IR��N
ʞm�m7~���+#�Y��Mb��ۀf�(�8��J����8y���5���O��E�բ-po�qV��h$*��Y�y2!#�>�4�]#Z�a-rL�y���Y�ZT_�� �+�v�V���	�te{G��k3���%���[N�F_'�����$\j�e>WM���6r.\�w�� �'�%*_�y�и%�E�M TWð�\�bNI[z�E�Ji�Dn��|s3p�(���<��:(�@d�U�q�&���qa�B���m��h|:��DC�0��;��mևȔ�<+P3[�n*��f��� l��I�>4�I��bQ���򾃖��s�qD H�����~�P���`�1��y�G�0� �7���	i6�+�IE��ϴ$�N8N�6��{0Npe-��uW�>�}�x���s�&��?�����뎺�A�Ϣ�y��;c:)�Q�6
�i�H��z����i��<�J1�?�Md���Q	���e��r��/N�d�907��K��k׿�i�(9o�i6�_���f"�R�r!�T>���Rτ�$��ܦ%�����w���%~��$��];z�KU�Z$n��&Vy�d��y��i�+�ow�6I����/r��mx��?e*�/lІebR�*��ӡ���i���U��Ue��	��Vϔm��6��b6��ڪ�|�}�d3>]y#�,�R-J{�R��1�%9���BݙU�1��Y0D_�T
����F���݇��̤�~�bח(�/i=P�Ơ��r�\���TH��?c��d�O���K1F�pWZ'�����?���mn��	Zr��z�ГN$hεy[�����1��f����FF8,�ʟi!�>s��fBi�Ƹ���8��acu*\�42�tW\b H���w���1u�@�����
Lӟd��N��pH^ ��Y�!�Q�֫{4m&�Zdop.�LBA ���I��)���4�^�nYA㩌�i=c�t�fq��hsO@�5,����M
Bu3<Nܔ˷���)`�0�wOR��#��sZ���خ%���K���k�Vl�{!Ug���Ϝ�3
l�͆�[�L��bs������^�s���
u����gﭻϼ�՗}�2���L�U�4��k���kb��]ө?h���_����� �����~L���5� ��hZS����ڟQf�w�J�H��l����}o��0�j~���7N�6�e�ڔ6S�@�O�φӹ> �Y2#۬���K|Ц>�@[F�]Gi*6^]V��(9�h��=+O"1�J�Z�Uh�޳1aU�i�S;m-j���N�4d[JB)� ����N|:��|��Ja:�������k��?qo�i�)z���`F�Y�ɪ�2�Yw-��m/��ֆ!�y��`��z�LG�#��ԈF)��2��I#�c����=]TM��ՙ��͋b�:LI~��H�BOb��;���	fI����)
O a��[@�(�ğ�"����Fs���5���t�\��ae�%��佂O	�����hw��[��6	��8�O$D���s�j�챇�N�F������z$;K���ʃ����,�/?mOM�|L��e���징��wD�993[)�#VF+�?�#0eyb�kZ��=fAf�k�}��Gx�a�5ao"�iW%�yX��<eP?4�f�<P��*Ѡ?֦tY�jh�D�6J2�pӰ�R��Y�s��82�4�u/�Ҍ�{���������b!���À��Ǔ&I4�b�P���Vz����[|��y�~��\�8�q��������.C+	�c܃��4��ְ#\|�|��F@p��hĦ��<1����������'�В���e�>�܁�F»ؤq�7�<���6䴔r_����=��8zׂ /�Ȳ���H�śb`BU+y�n.�����웏�����6��G�4�q�:�ʎ×������Y��Jz�� �W䪟ш�BEڌ��Q�U��jA�j,����vt��Q�����㤣l��	?�O(k	�^�@~W�8��gs��8a��A�r��O�@��u�����T,��ᶙ%�{�]Iô<m���,Q��P��;�p~��૜��ȑ��6Hⷯ����T{_��jo��;}U���BX��i�߬"����ȇ�4�l��mbY�����G�x�W� 2���~��أ�`Џw�_��������E��f�^~m����Tڪ��W[ ���=��8��B����Dg��Bb?�?$��\ESY!C.�v���)���$���s�'���7	��D��'�ȹ̾�W����*I���͋.��k���V'�:�<��ﺤ\��v��hf��������୲��aI\��&�u�>���X��������N�b�׎6)3���B�B|� Ċ �	o�ǰ.#��[����O'���DƌA�O���A\-�[�O�R+�Im%��h�2Փ;�n�2n=��k��2YF�nM3�b, '3	>Cz���8W�AI��(46�~K��b����ʯ�t���^��{I��ugZ\�^�fMU�黶_�ɄE�(^1q鯜E��w�̃:�ه��`I���Л�D_�:�#{�gW�9�R����i��>�]�<�9�R䑧ӹrƕ>��'��t�=N�kI���AjU�W;�ǽ*�a�ZÌ� �|%d�\u�K��i����xOb9��]�}k����h��5���ץ�<Ǝ{V��0	��5,�}#���fi����New3��qOv2�zx��w�Ŭ�����}��?d��5�j���!�B�EAG�M�Э],��P���k1�}�kX�/;����B4����*$�]BO�%0�;`I�,��[{Y�w�c���[J���+�V�k��u�m��X�֓
�-�o^�<�Ś�؂Ԧ�9Ps�D�+� upm��D^b��S04�(��^��%��n�AYS�V:���bۥ��5�4��/vu^��QY�x�qdlI�]�� �y���_��\���i��22��3��f��K"��4�?�`*�9(�Jd+�H���ӫƦ�sF�:E�v%�$�M�����g#?��%}Xj��� ��-><��6��W�⩫�n��U����E5$�(���Z4�}�1��e��3�� �bS�m�L�"*�Lˏ�PN9!�g�q�Ѓ��n]��ӺI�w[2����WI�Z��:�8�?�}����cn��;͗���T�$�Y�EJA�~�F��w� �Bhf{��*ù�H	�1WĲ�)�����Ɠ�-*72!�����_ݺ<����3^�s�9��wFw9=97׵�ӳ�-����YHRR_�@TK"�^.��x�]jł�I��;M�E��է��OP5r��o���d��C��^��s{O�T�M:1�n�����0b�X��UT�,0����޻�
"u�����y�l͑:V�b�������J�bCtu�y�UoR*��QN���f�R�\ඥ줃98�@�R�5cGCOrF�������S� �C:�!�ã|se�d�c�֍V�
��i�P1C�$ XFU�1y|�O�����՜�(� �vH�����D��S��1�<e�n	� 0E��V̿�7P]e����Ơ�`�iB�-�O��/JO�?�u)c�b�n��l8C�c.�gV-�?ui_�~�p��tv�nSTl�9$��=��]��3E>��;��ПCq�h/�����e,T�i�=�tP����]�\H��4`i�K'�&U0-��klEfrdZ���l��",
L��IWD���i"h��á�v��w�lA�T���;�K2U�����l���Mºʣ���3�V��m�E����l��4)}��g���C̸[��k�`��~�sa<Y������@W�K,��C�X�RX�-/S�BGG'��&.os�RU���|���16(&���}����C�H���zk�Y���6)��+�
�EI���$���+A�8*�U�6����&ƼMO8�3ިU������&�eť̋��yH`�βM!����8��b"k	�taN7cM�P#q��!��D�w�i�Q�x\�iT�;2(�U󻜚¦$��b�N���c#}�ҏ��-ĺ!
��-^��١y��,�O��4qU
����ڹL���E"�)�T)t���F�6�t����SE�lD�|�7Y�m���n߱ϥ�q�"�&ʾ�mz�$�-���c���\��K�j�R�w��=�"�"%�m:H]C��~�X�-{��r��Jf-8�mX�arLpy��>ƣ�~M�b�xh�/�\�{��ȡs��A4���~*��fR:rZx�v:0W�������2 @��7cJ�nY��{���;O�Y"�UX��	��Ŵ$���p��l�1�kƚ{�}��0)����{�Df
���ξ#?�5'҂B�T26��l�D�asG^Z��1 �x1"�(���ج��[Z��%+�t�.�B�bǝAzw��yPm�V��>����e,���nm��S���Ս���OPj:[���zS��UmE�I��2��[��m!\ 6o�e���"�a%d���."s�ذ����ә5H�V���F�5�Q�W�9�La����ZH�� �u�d���>f�����l��t��TDB��o��@��D/�ժ�3�z�Nz�%6��vF��+N)f�5f�y�:��W|Ԃbc�k�04����v�_�S���*����	4�>����.|�KH�����X�v���]؎+#>�:�dx�5��V��i	��?�C~�Y��1P-B�PE7,�U{��2u�`��s'��k���zC���y�./��G9��'v�AlA���j;�Q�Ƨ���~k�O�s�S�@�`��)�eJ$��?�������j������Xہ�5�w��t���Y���|!@�wCBυG�	���࿽�4l����{�4P�Ш�	��S̵{��o�N��p(4�0�F�I3�1�ۜ��d`p5��%��w0 F���[^�ϱ��9��=�*-}V�ˈ�k@o����]���ne՘6�� �-��ե�6�e��b{-FF�BSn��_H��ڎ0�2�C�;�8�/�i��tw�l���W��VF�;J
���3���h�PfdJ��"�Ud��R���mAqW5C�A��bC���xW��P��8{�&�c��������t��L��E���N�Rg��2�3]����Ps����.͔��@�Z˒� ���q�������]�:��
F��0�* �����D�m���'��+��t���E�3`\����j]*���0�aX�+���i��fج��E�|�t]1�l#c�>��� s W*�Z,Wy��-zg�Ыf�I��F�"T�,m�]��ypz��9��8,�n�crB�%d9]�u�o�cX�u!#�tB_��ؖ��-	�'�$�(����O�X�����&�eyv�c�9�P�q"m޺h� >����oh=����0�Fj�P���|x� F
v����n%Ҥ�h;�!�<Ӽ7�|�]u���v���H�i�֗�RWX;S�=h�U��v톐DԅNj�	d&!H�=R�QW�fd�ڶ��f�+�h�EJ��/ ��(,U�x=�&�I��Ѓ���!�����>�����I�V&�`�`��p��T#?/q5�]�E�<��f�<�D.s�c��'��+O�;즒��;� +����&���U��@~`O��� %[�٫��Z�yB�~.sB�V�tĈBM,��3�5�V>sï�8a�*�R�&>�#�À�l0����k�=�(����~����\�_y�DtLqH�?X�IL���d�cr54�O7��A 8=+�cX�QE��\����	r�2)Ua��3��ꃿCb�����͟]NtDj���~ƮЯ�i%�!r�u �y����э��Z<U}@N$A�m�����Ao� PWJ�^�9$�E��0숥'��ax�.��D��K�ד8�T|6˂�3+X)|��n��zu��P5:�wr��(ߎB��h�' K֒k���^S̝uo���%A #@�֡?BƟ�D� ���Y�m̨�H^�R9v6S.�p����y�ʧ���FY;�$��L���X" ��CD���p ��Щh�g�^�b��"D�'������֛O�����·�C%��=sY���b7�a�	^��j�'*��V&�a>�b���P�ԙ�Y�=W�<?������t=1w;8A���Fbz�kא.�~�����V�5�����$�M�i�r�B6?�h�,2��]ȑ�X���B�y�݅B�)���Ei
��	� ��.����!���aݱ���ܨ�_������q$�G"�@��	���_VzV��jB��H��5`����x�%H�@9�q5�\�33���ަ�ͽF�R��F�$F�lyf��3L�ǡ���뤉H�M���1on}��0o^�!��ƛ_��cY�d���96?����_aJc:��Ƹ�EM�k�r���FCPsڣL	c����˧d=����G��z��`2��,�����V���)��9����AG�*Xu^97�{�~ڕ'
zAq�G�UQ��@�'c�Gb�i[w+��I�����)̬�h^��q�}��-��𳖞�^Ԏh��*�)/<Մ?�$:vq_�u)�B4X�)d�e��MTt�F�,����������C"^��z�y�{[��jN�<%�cO�M#�h# �ත�����xm���%�Q�PXu�Fby$Np��</�[��!v��oHw�L3E�R�o�z����D�６d[��O0�:���\ݳ��vۨ��[�5^	��+Y��B10�x�����~Z��(�74�m���ex��������+0T9�3������?A	LA�q�� �l$iBg� ��Q�n��W�o��_��f`gʫWG���M�B��� Q
Nr�'(Fe�
(�Jw�\���`�._5T����k43I E+x+Q���S\/xՊ��KvH��2 �Ô��0�{��l� �ب��˫�?����Qv�6��D2�ߐ	lf���b��S�ٞ��v#��s>+`d	s��u|���,�������VB2�����>�g�v;�c��0ڥP8���
@�{���  XL.�����üm~�@6��fz6��-%���&��BY��Ҁ���]�  ^X�W��9�c��I�z�`��z�V 9%번�m�I���|Y)�0�v�����j}3���@�O?A���M�������t��5�P�K��Q,�礢 cڲ��}k��p�D2��Y��"-l��
/�4!g�]�����bmc���wF����v~d=�8U^��5�*$u��z�I˚��M�W�����ݒ��7�����|��!��q��Ca?"W�:q���u��^��k��^��a܀4�O,('3\�اf\� ~j������<��K�XjVC�(Eu< W�#��̙fӵ�Ը�W����H�P~�]hb�+�݁�%zV�`F�����'L�xL�;5�t�P�b�v<�݉��2�ʼ��>�ߺd["<Ԉ�AXf �ۂ �܆��4��&}i���ꥥq�>�'Ÿ`%AN7P���p�W�~���T$$��Weh7��+jG��gP�:ʮ3)�{���S����"JN��*�E�ǘ9Bq����bRX:cK/ܥyʓ��p�K��<49�ȮOI�ğ0Qu��a�t���y^V/ι����
$t���w?�����f[,�7NP�M��u`60`�o
�+�Q��!�a���Yt�h%nʶbC1Y�o�@� $���Ew�n}hwY墟`E@0Ðt�z(�N�PX��l�].�ܴ
Ӄq>2��]K�P�͸g5h����㴡x��$m���L����|�ϭ�����h[0�jR����@�ѷ��S,B�4c0�)������;K/ץ0뒉Gf����	ѓ(ś'�.�:��/)�JdI�[SE�1n����!(8o���G�	�1���I���,
�ka
̀��d��)7����)���O_<#�ؚ���H�03�\��r�s@^]~xD��_�����*'!8�u7�ٝ<��ؽ��0��{�p��V�2���#��~��a��[`�!%b���))��Z*�g僲�`�e���5�s��p�A�o]F���S��q�1.)Ś�H����ѽ���!�WD:S��c\�����]{2hX� =Ɯ� 90(�P%�4����T=_��r�1b��?���UP��\ߕ���	� nI�]I��1a3��d����g�\nӘMP�c;Fy_F5K���=ےj��H�����+h=܍�����}]��M��ĥkc����+5�N�AT�a T�T��7ϼ�� f�{�ٹ䟳2�i)4_�����݄�Z�\>�eY^��~#��q�X�����BX�^w{x#��yŌ��t�������+!4 5�	���aC��)�(�TXBY�����Y�g��Y�F��Y�C.�J+����8bHF��(����?{���ѩ�tG?d�Q��O�S��S�g����5h��<R3����"6���p�H�o��i%W��T�K�+p��2oV�t>����^�i�/H{��AѤ�$��DOP>}��Q�����*��3�D�.��V&E�z9X��U�Ι��"5�t�-v��4�g���ٛaz�n�b��WVT���f1í��ICҝn�ۭ�B�����IQ������_mH\],"$8#�e&�����a�����L�-��"��VR� �����@~@�u��?J\��	��kJTX�`|-�a&GR�g���<��0ull1���)���h��ޭ i�V����:Q%�_|P	��ě�)v�c>���I�	��x�%�͞(`�������.�����r�sIIi�$`�$��9\>-�+������J�h��[���ŨD�s�.� N[n�`�w�k�$�,"�E[��]�Q�P��?N��2T$�\�켆��)��W��[�|>*?E�W��j�A+C2Y^��I3�
b�tu�]��Vf�f �P������#g��މU���l��j*Ŋ�CI�����T�%�s��&��rx��D?��(�ܻ�u!��G�Ҋ�X%kt6�COΩƢ\R��tU�,T���,t��w,:G�^���݃h��+u>"9d�0�*N��x-q��Kݫ@"W�}��&7��$�G�'�r-��_R��Ryx�/�`�P;���@�K� ��{%y+i|�!k/���0�����ae�_[+N�5�X��(#���h�o^U�Ҹ��.3$㍎�M��*��%6_t� �7���ֶ551
�yn�:W�H]kBY�󫳉�������L��9��X�g2bC�c�����A�����8)Bfw�3wv��}Z��`�*��M!�;���+�)#�c���`��/�X��]aا��f-�萁_W)�w.��f�n��3OɊ����3��'�E����T�>��^$����EycS�/8B��z
f}���B��5��mE�ة#E �<t�R���u�'Hk�~{s��d��6퍺�8�R��%
�yި���y�&m���7:�|@=JC�UECC�Z���%�s  ��W�ȸG.%������K�μ�N�	�a�]ms��v+�
�-ИL����l�v�i:A��<���B�xzh�P��_��[)���F4����:��^�͂�����P��6[{H��������{p넁�k�wa|�9qV�X�k\�`����<���I���%.W����{�����t�м�d[*8�D�G��|�w~��t8іU��0�t�Nd��hF��D�_�y^H�q�֊Nz��8&p&*.u���E�3�𒌡�������9����3� �ȝ ��IK�\�x�9�5��DF�U��u��f!�6��!�|�fɹ,��̓�[��a'���n�ShJ~�D~^�]�!ZƢ�M�sC�>�G�h^�0@u]W/,v�꘎H�m�6��h�^s`��y	v$h�5.d�p�û�?T�9+�l�����`�Ը-�!�?!��I"�1���T����M�Q����W�?�
��|B��&�E�4�Ƀ*u�cg,��|�u,���P����3 �T�'���yv]�9,��{�Y�ʝ�/��ZX7^��ر�P	K��P�]Il�:a������&��s�T��8�?�Ņ�V�Yj	)"n�Gl|kq�Ov���\n��7f��/�Wq/�l_�}WͶ����S�W��Sˋ9���~��{;�2�iڅP�7���
��+�q���6���t���J���K4-H�{��WP=]�;Mp1i%K�}ɔ^H����Uۏ��.&-u����'�b�ބ�����g�Y�wNl>��Sl��GRf���o5�Cؾ�����V=z2K����nFnj1�[|��h��譃U���+~��4U�bm�� �)A�$q��@8�I<�T �8�yM��̹s�N�	٠�����A��h��H%Up�1�qA�I������Q�3�]_�_dB��������L���(�2 �p���l{8���2>�ʟfs_p�/������1� �X�r�e��|Hݾh�I�����N����@���C�y5�h��ev��P��\�Hu�����R��������*̨0��?}�����Y3���$/���'�а�2�ڈ��>�B b�m�>ُo����PN�#ɒ��	ۉ@��[��c��IQ ��k��Tڢ9���޷?��ɥ:��Bs� ��Q���8dN�hCa�yJ���r(>�\u1�A�t������R�q�H�#3v9�͈j�����?�5gҁJ�8l|<�
:��dE�R�����24���(�`6����� \��!f~H0��d¨��p1h���lGu�1i鼡'fJ����As,�w֞>��Vl4����t��X��\�fddl	1��]T�h<i�h;L
Vu�;�Ibi.[��,��[�����K]x�͋���}�俕�d��<@�8��y�G�3P�-ø��m]9A&R��	���5�,�^}�W0pV�i�����-���Ȝ���sWýM�Q�É�߳�G��2PO׆޴�F5>&�h�h�ka��;��fWg��0?K#��f�ԋ�7uwt� G0-6 ��5��YD�s�{���O�< �ˉ~B��^#�_E\78�Ӿi/�g��+�g �5_,�]�Ym��� 7Bs�*T�j�����/V�BV����]�o
E�eT��(��v+�,R�T��H�S�\ZtC��U�~M �˾�~u�6(�Ԓ���m�t�W�q��)=eU=�;λ̌hV���3�捺�;���ί���ɣÅ%�
�ߑ�a��@+��^�6E�)���g�����:��ՠu5�d�|GO��	���Lt����ؤ	r���1���u5$��.>�|���r�~��!��9#�DI�A��Ϥk�,Y�'������N6N�-_�K�ʑAY�I�j~>NK�3���]�t|,^������=�5a�b�Z ���(޷W��h�{904���2o�x14@B �PB�����O������lŁ�	����
Dż;i��r��lgɂ����-�uB�%��_'+�BYs �	����N-w-��8�ջl8B���y�e�ȍMa�NIb�	8m#fA���Za~%��X-m�?����7�w�;��4 #Ƶs�J�`!AQ_�~@��x�~�R��)�����v˂�U�X�%D�aw�/eM%r{`�f�Ʒ��� w>�Jd�oΧtm|\^�*��ے���?�O${Y�!c������w���c���]\܉Xӕ2q��7'�����:���ᤑa@�D�{��<!*F�oO�Þ�ү9X���=�x���\�	 	�UW� �9�IK	}��z�ov�w�Ɠ"&0y�|���JH�1OxvھP2�x�@$��3|7���$�4I;���U�cXJy��,�W)o�7�>�5�|�l2eG�z[��jf�1�,��`��!�i!�"1)��i����9�����|ѓ�UL��t��h\�#'�aC]�/M����e����6=�fL�y�z�J�F�2�(���U��MT��l
Hh��VO�pi)����&���w!���������Gs��Ogz��cVm'�d�q��K�0_� )X�h/ݰZj����L���v�J;��i�&y@Izjl��ǨPX�%���DZ�;��!�u���
�{�e"<�L-Qx2������������zN�owq�&2=���s0�N?R� 3�����v3;\�L�Rz�2��L&cR�'OD$��b4�rW�_j��]���A?����}Q�	�9x�q��e�N"Mϖ 
��|9	f���v�T��>؃�{1l�����K�$��	<1(�(Ԉ�\�]ޔi'�ɴV*�_b�q�b������ޝ[�H��Y�=w���T�{��XK�:Mo�FA()��Tg�6"y��z��W�Q^����F�⭝�T�A��N���
���:��e���ֱ��	v⊅:��u�%J_pTԎ	��O�n�6�V8~�^^�?�}���ٶ����[��1'd�p}͙^Q��(�6+��FF0��⥈��}�!&rq�lT.�&:�q�RX��b�;���'�CKs�YZ(����נ^�����*�S�V����5x';ڂ��u�P����Nǖ��|ybMN���M�(,ʨ(�~}�H�����S��1V�a���R#��}p�~ �0��I�CqUU�.�τ�D���I������f:h��0��-Qk\�`"S�/:�3��1��7�_k���k����H}Z�O�¿�1mx�36��ѧT=M0	z��ϟ�@�Gy~�K��8I�K/������� |K"�s*'Ӈ�1�;+����J��1';�����;ү4�#Ȃr�{����M�����by�ف8������ۗ��a��Z�s��k˗��2��qD��9p�E�n�
*D��B�VYe2��f��s�"�x��9Wi�����Ԗ��B+�((,&��Y��U������A�@O�=pH��*-���t?v:�(&�B�K�/v�Λ� �[��`-�NL��@L��=��) &�5�9�u���.�z�?���!�=��ـ��/����)B|�o2g��s���[���~@�!N�N���Cj����:�!��z��i�8C�UD�0tJ囃=�S8b�gJ�&4Czj ݚ��7���j��#A��`X^u绵,�)��j�%$�p;�eO��_��<�F�t5~iq�;ǝ���<��Zk�:�G(�*�^amW��_�'#F₳�̰�(����jL�#gA ��(�܏nٍ����L�z�#)��O�_�FɁ���}I]�U��=�ލ#�JӀ��Av>9�`�.�llt+<�+�r�@�&�����=;�[��v+@��b�j���Wr�a��uGU��\�=1O�nQⰮ=
������_�.
c{�������S�&��b^��X�rTMl�"N�gs%⚲M�x:o���ϿM"�	ze����k7!���AJt�?�W�Cc�m=���A"���e����}w�2'��o�Mz��ѥ{���L�A<�WG�J^�vH���� |�����4��w\ɾ�mU��P�����7Wk�{|�v#|oE�"��s���w	���9���4�J�o�Ia�W��(w�!��uXHgE�h[�A-�: Ґ�ǭ�^����%|�I��Jh,�YWQ9�ī��.�>�g9��AX��"������bo���͎���i��싫��!	Jd �@bi��՞�l_XC�m��*���mD�1�I�`��V�f�MMT����C�(�T
��"�@3�31�É�����ie�L"(�ě����.�����p'Y�;�qk�EK�U�[�-�s�r�;��`2�rM��B^�)����2!Z�t�4�Ј���g1��E������V�w�|�
x�D�����㈦��n��I[����EH˿s�R�M,+ʜ7��������j��f�M<��|%\x��]�"(��Ջ�T|4�L�(���j���а̠���/S��7�qw<hW������a�OxSH����'���)�P��֨d�\:x��݇��a$;e6�D� O%���2o���i�Fm���e|���θ
����T� ķK��FZ�&!Z��V8�ɉ~�M�>_��V!�̏��oz ᐑW��[��� ,Y��������5�j*ich�=u��A\��`��C�SJ�ͯ���yIv�@�9�b[^~T27w��]i?U&�nM���7�
�K�Tr�B&�f_�\OjpP#5S���-�y�J��b�S,�Ը��UvL5��vV���i�'��3�͵,��@YN��P���a���G�}P�Ϲ��&+�^g��n8VL�gф��!�~撆������uj*/����������������04��f��zVx��^%7�Ӄf&Z��{����kky����N�R�P�̽\G x��C(��o�G�l�w�.|�C�w��*+�ߒ�Ă�O�J�}	8@��s�7�x�Jy?���Μ*h~b|+��dL��b�i�ml�gC!.`�&
Xu���d��
�����!�z+���hy8 ���_��xY��h�Q����Œ$�/T����
���G��yI�	7��g�,��p5g��B��=Q��,��K�b!�s%�Q{6�Uy=����rS0O)d��2I5�G�-Ta΢��ꌫę1*��83:�e�FF�mVEM���X�۝ݣG����ȩ:0�Ԓq��8���*U!��9sɝ�����0��-�:r�����+���e��r��njR�Q�^^[u"�7цΛ��]+�)!]F�>�i%�Hݍ�%��>��1�������XoQ���OQ��ީj�5�*X�O��ڿ]WCQ�!���5Y-�u�H�I�'l阁a^Tt�fO�J�
}��+	áN���)��y;�_�42�������a�z���-d�� 㯰�b��-�T�ݠ0�e��=cԺ�XAFl���Y� �ׄx.c��&@ٶ�K��W���`
��|�S�[�(���HA�Y7��AK�⠎�)�U�*U�>qe�M;�*�ê�1K�n�g0Bk��f����)���p�1�+�|����vVߠ2�����L�1�|M����8���s�{p�Lu!��(��^���߁��N��	�ȻM2�!C7��]�{��[�ӹ:d�އ�u �?��Y�Hi@Q��(/��'�f=�;����m~{t��J��K�ԊS�O�m�tԒ�hx�k�kϗ���6��5�B�ȗj:-�1�o�-}=��l I^�z7�l�ؤ�Ē�*u���u��������b���<��#v>����k��������� �鞂Wۨ�=֊�����Z��}�W�>NWaSZ*�B���Ց,��c2��b}~���
���y�2��>*,L��fRG��̹�s����8��r󏸶^u����L��4��e��E�h�k�Uk��A��S�~��F���BΟ�ֿpk/Q�4����ڒ.�&`�M:h�+�8
AX����]&$e�8�h�lw�V��	��kO��Y�Ŧ=���b��Z��aj�Y�ʤ>��{8��,Ѷ�7��&&�T�ХFI0�}�j2�i�.����i�GDA_���	QEV	E��c����|��.�A8�b���Q��Xm���5=rn=Ba��O��FR�ZӿE7!`�h+�0�Θ8�0 ��qg������!�H�ȇn&s�d
,�+x�QC>l92�������k#`g�s���x�q��[��ȴ�C�0d��G�}�+-�r1�]���"7��ّ�	�z鼜�z�s�ed�3���*I<h4����L����������)q^�
,b߷�?�HT��h���/*�W�Gr��#�}hk+��kQx�\t�
����2���t��U�'�]����MN��T[�&j��ko%6o�����O:z����sd�V0(Q|٥�u�3 �̹h�=rE�S�@Z2�2���̢�d`�JD7BI S�; x���F����C)�|X��Χ��� NX�mL�j�f�h�޼؝�?���y�&R&�MtaX�-�EY�A|Wg�N��s{~%����|�"N����.}�灃_	���[lӕ��jq�}�8��S�T538�r6̺/>�V���5�5��i���/i+���������Y0�ggYT��&և���9�J�L񈓯m=g�b:4�ԭ<���t����&�^l���C���ɔL�b�t������p�4�Q}�Ը�H�ǀӳ��,F��4�˶���u�& �7rQ�{��B��*f1w�&+mۼ(h�����K5N2��/W���0�O��p���*��K���?;��vv�i�6��Ń���b1��D�P��ݙ(��:?q���ymXuDl	��|�a�V���ZG�)@���wπ\= Š��\�,D{��!A=���E�Rд���?y6#E*���ÝJ	�F4(�sdR[z�z�����z����1܋^����z1���hA� Ν@���Xf��k�sl�P!�.����^�ob(mgP
m�)o%'=���D�Y;���,�0-MI��Y�*[u����ݡ����w�'����E�q�@?�%���!�F�eà�P(��y�	���V$�B(�����\i�Wh��䟑H�eܾ謱��v��hk�x�ퟒ?w���F,<�	N��H�e�I�(4�������H�����1��8���b��$��4�x��)�����-��Q!v׈�R��|[ӟ�r�g{����(�+ϊ����Z�{�l��E�\��yߠ�Y7�����C��Ċ����Wr|��ו�f�1���_Y3��d�p�x=�	���ci#�aI^�¾	�罎?�d��j��ZR��f�p@�ߜ��W�P��a
��b�E�ɸ<Ћ��*2o����9l�?���VY�W5ϨT.�S�+��'J�!��q�Ď����G����7�[=�2$����ܴ�:�^]�W�7��dv>k��`>V�"f$9��v{�WQ`�д���c[r��� �&^	�m���a�SѠ�zK#T�[n]��(���&��B=����i�xu��2��1����#����*�����N�p:m��`�����M{gWC����;ᜨ��9��[�O8��]���AgjVc1��� ��ό�M�2��0�[�tw����ܟ*k��G-��[��~��8��֖1#���2��l��!�� ;E}�.
���<�'0�d��n +�R_�2W��K9�q�}����oG�Ҳ��G�#6H�e:�!�E�N-���h�\Su���G�̈́�/��}}��4��T&�Ij�PN��9�k��(�=��S{_�D-��w���wS���Z`s��gՆ�
�$6ERo�����l�jI���g{u>Vk5ɭM��6�۴�gR��Ns�L㙦x��={�W�{�>H<�Q+���a�������"եq����y��o��;�����am���-O�=���f����U��k�&ǀQ�Q@��b4��(��ۯ�=ʵ���ە>J Bfq!:�)����Bɐ��l����[$bIٻM��#�9 l��5�7��Z�/�U����)��;�9�F�
���b��E竹m׎0��2�:g������%.0�)��&�Ū�M37�7�7����92��$���c�q&�:����{U_�B��sو��@�ϡe�t�	�lH:�K����L��-[�@Zh��ߥ$c����+&;i7���LYh����$�'�V�]3��I����f���s	o��36�H��;H:&ʱ<������?�W[�5E>eO�e5}���&t�*4m�j*-���i��C�r�0��g���!�n
W��'a}0c�f�d�'�zG ����/g4��g>��!����>pI��xp$�`��qO�9���'�G�v�X?0	�_;ʒ9y����94��o���D��J_���q��s$�1S%`C�����!2����М^vFV��R��IkKo�
�-�^Lp�q�,�w��1����C�⠣�f��%_�'	U�96#����5�~g_��*s^�ѯ��+.��D[��ԆO�w�\M�Ƀ��oY����UK�Z���2�)g� C�Ÿ}��"���ݼS�����I�e�׺0�r�5&��g���S��i�!�4��@�XGu@J}�����w���}�P2�z)��ָ�M#F#2�%y�'a�v�I7�)^	����B'LK�6@�G'B��B��'�D�����	;�6�7)+�Q�D��-���;Y��6�\;1��CK�%P((M��w[�b��XQi�؄195�{���%"�����Kd]��Z���0��^�&��I�2��c9�?}����'�_��>���x~.���qf�wc�
��_:����1Y����:ڢ��<iS����c��N� _;Ō�F38��X/ϭ��Dv�z�<���a_��%������;0���s�-^7M�Lz-��[���
��N��$1�?�M��q��4���1&�.Ih�8*�G�* �v�rX���.EA�Y��9%�A�-�S�^�g���S����f\�ď���.�#�q�C02�G��Zl��F����٣�m�1�n �=>A�'O�s~�*kO@Q^��<����x��u?2Zp�(h'^�wN0��v�M��c�+y��0�{z���R�9�rs?�����0�c�/l��5�*�(l�A��m-�0(�Dߴ�N�?�Vɰa@�����{i��p��R:��?:�e�P]�J�p�����i鸺�Q����!���'���D �l����fM��)]1�ѸjR_�H��diXi�\v!8b��+���4�e����ȱ+ v�sz6�[	<}�GP��Q��<�eO���"'~JS�Lfz�� ݑ�FrP$���=��Շ���z�e)�h���rJi�F�\��e,py��T@���?_����r,"2����ָ�='���v-MKt���,%ퟥl��Y'SX_9[$��z�^���W_=����R��v�S+��0�P�5`#���٫k�fFX�H19����Q<�|�H6�k��H	�-%e��g�<Rf['�����30$)%�/�߰d�\|^B�r����U���Ϥ��@�g�_�mj���xa�hI�>u̕��������AN�;�t @�.E�Lx���|RCv5��ܗ�����+�̟
S�o��a{o�o=�_��'4*{-?�d��.>�������&�/�P�Bz=�n%��=���:*�w~_??䟎QE[)s���!��G�x�h�1�H����};��z�=������Zi*�y2u;m�CF�?��U��wLT9p�z5�Yħ썮�	
��'Tʎ/}Z2aH����c�OZ��za�L����>��&V��ߙ�޶r?(�]����5icU�U��Ч�7�����I3���u�vL	Q���Xzsh��6�)���%[��I\�:VJD�Q�Z$�����@�Y�wj8����vk *��-n��J�Wmh�8U���L͇,�}VA\�F��
DO~j�����˃���[�0�mZ�AYL�9�Hx��(�;]�Edɐ���ވ�qr����8�a!���z9@(Ig0%�MD����o�����������®���D���2�Ga��!�'Sr��.	a��-$ͦ����T�v�╗V��Y��l�@�d�}{��*�8&�=���^e�$����G��P��¬UL�����o������������sz?j���@���mbz��7R�-S��P�4ְ��ă$���h&�Mls{��»\ƌN�M�Æ���θ>H�t=2�\GU�s�D��<���c�&�b�D���'G`�\����kn���R�����t���_�ֶM
9���퉁��i�Y��1aO介��0�]^*�⢉=��N��l�Z�%���%m����ʫ�'��e�h�M�N��-�d.��z�*�f�h$}m��lQ��3QNc��H����&G.t��G]�2�q��Ҥr����h�_�����Z:��=�K��ڽp�!�)o�pX����0�Fꆌ�;I�82�BoMpF��y��ݼ�[����1Z��{�M�D�	�0��ҳh����=�䀋�+z��MÒv�$��z��F��h�f�ɍ���B?27��2u�O� Y��)��]̂�h�f�m�0�!#��4����]Ƶo�����o�5#|Y���`D���ք<�ؐ4�f:�Na�7��l.$vd�l������7�E���L/���eY�\���8�a:JYT��ϱ��j^�U:WrL>�Fd���.[���I��sv_�Rޣ� qD�I�xa����	�U�V!F���z$|:Y���p��I��e�p�����R��SJ�\�C��X���)��#���0���%^i	bGO�eu&/�]g�f%��pt�=�V҈*A~��G	�I�v{=�.{5/ᰶ�ɭ�{�2ǔ`�C&,xE����v�u��oN�zXWxl�x�"_�+�	��ڧH��7d�ˑ��M�
�m2�t���p�o0��1�np��?3[��������?�D�4��sҘQ�>CY�ʍ�6����z簛�w���$����D�c!Ư	�ԣ��/�`�Y<���Zë�B9B��*��75�N�����<�ܓ�Oj��j0L#kE�����o���0�˟j����.z�W.� D0���lG��Y�Ds��bgr�8J��b�]5���㙹-r�i��48�w5t*]@	��� I_	�q�J��4iɝ<��ޒ�>=�R�2§�d�ܞ��P{���ɏ�����ts�!GOE<�6��k�L�qQn�(#�h_L�⺡�ٗ�R?OqS����*����c:��${d�aI|��X�0��WM�Sb��}��؂5�~�����4�/m�vge����"��haV�3W��κ�[��P��O������*ȭ׫�䀃����i��{'%_��?7j�ڵߏVB�*^F�G��A���~� ��΂d����pܘAHo��m0�j<�23{��8L����*f"�U�ݪ�a�Md >؎�=������m��]VN��(��[��� ��E�����Q��_� 4��Q=#գ1F�x����TG{F	�YD>�(Y��o�>�A�m��J�A��G��n�^���f����м;�v�My��B���Ϩ�#�q0�Ot[�M=U]�P��NoD���w�=�.`�x��^B?y;:dY�&.q߬�M�Iqw1f�м��m�w�9� oZ��h2�[�YѲ�d�Ҕ_7Jz��݇��x �57"���	���7{�]F۷p�哟�0Aঋ�@��?����o���e��O6��t�:
�:�E�C:�^No.�1�&���{�����*#���)���EzT��cW�}�K
,��h]�a	(�8��Z�^�g��d�t�1a+�M��mD~�bd�?A��
��<b�b�7S�W]����)W�m �]a�`L�R�ʓ��;�����_K�XIU��v±Y��ϒ�?>m�\ϑg"R���\R����+ilm��Rޢsf6w9�~;���z��,ɻ�@]�7�D��ա�B��c��\*԰�h���ln���ϑ�)0�ZY��'e+
H�i�8���;��Du�R��+�K;UI8+^�0�+Q�[�o��R��\��.x�
-B��4eF�.|�- H�tʑ��X�Y�$Pe\N�+��D�K�D�A�BUИ$F�1���	[��cqA�mb�: �*��a8�?��#:�/]S8G��g�>xh�Ej@���\i
#��}��A�.#��0�9���u������qT�$��hN���౴v��`�΅�}��Q�ܢ�)�r�D�$������8��s���}1%����^T�N<��j�ǥ+[.���3Y�37�~���'��S�n��ւ�g{����d�M�����i~�6���H�'K9(��(���1�x�t@
������ k�7=���jz��^yV�*�+._���ksD����y舫�;�Fy6",�H ��ō?����@i�z�ǋ����I�+ID1��oTm���m�[U�zO@�e�o3'���EC+:��#Es�[[Hܛ�=Pߟ����V��G�~+���5���E��V.M%�O).��nb�Y@�G��	{;�o��9�V��!�5_\ ��}`�Úr�������Ƴ��\x!�/x-��@��(�5�tĸ �oC��w=+=�Gb�h������Z?ZM���L�C�A/�;Psn��$tB<����<�`@C*X���ֳ��n���f>9cn<�@X�x��|��/���k���8���^9�G�qġx������$��o��io��
�V�d�ft�;��rK���������\3�;`�KJZ]�˙a�^�}A�����:c)'~����Hg�~�mErw!�*�2�pr5�����u�!!D��{j���t�K��Fk�</8H�eY11����c�'�~G���Ӽ�ze���ܴ2M���7;��,��$w�ȁ��چɘ!:��% _��ʀ)�����H��wf�e/ȰV	��N'���Ҿ͖a�5�q����C[ƑoO��RS'�`蹰��X[	E�yzZ�����ǔ�Y�/ϱR���P=XK����;����#��O��ΧS��A�~
��h(�zä���`��s��]�|��( ~6v��c��JY�y9Jc�]��!���6��O����_�b$.V����{�3�����`��^ڢ2CL�k.�}1���ۀ�弮�G��.P�{�k�'��rm��!<o��$/��ɍW�f��G�h��B|�Cg/�`J�o�Y����@�2+#&S��L�S�UC�)1� ?��&{}Q�S�<��LN{M��?r��;q���|]�)�,�t"�B�VE>߷�=� ũ�(���-��:}�VcrGS�8>��b�jN�����w�w84����<���
��/�c]f�BQ�����{>׹>^k7<�NM*d��3�M

ؓ�R���ݦ���×���k�Lk�'W�w)��7mh$!�(V�S>�A��,�N����i�\è@rBǄ5���#�M�M���s������b�*8;"�����Dlo\7`��r�y^�)F����\R��QT�H�Z�x?���|\����ѭ��wң��>3�x�X��w1>�j�
ŗo���9�Y!�K�9��k�|Ě�PG�DЯ]������(D)yx�B�}�o}M���ٙ@ e��B8Q[<�SƘ�i���| �%���r�V���U�*�~���W�BR
]�w�K��^��̅߁�:Z}�%�р�ylC q�_'h�>c��'%�/� ��]s`�C��2J��gw�����eR$]s�~�+,��ŭ�;�#)UW�b�Cg��#n������.Զ��S�	���mȨ���bN�Qe,(��)�pr���=�l_�lP@�����I+��c忑Ϟ���Aq���3�F��x���J� iU�o��+�~�S�c��M�F�(Tq�;Cm�3�k�_E�D`�яC�I>��B`)���n�DH^�	�-a7z ��S�e��-�g	�%�^$ ŉ�����G>��R]����jdl#ȯX�ݘ�,9w�BJOK�H��/��ó����k~����)nG�G�Nv�c-��Z��!e@B�Sn'�8�������t�i�aq��n��`�����[��.g���c�:ڰ�4܎��{���fk���@**���h}��A,�b7,.�n�_�l(����� v;��4��_�
��!����Gp�O���$�|gFBq!��V������8<T���"5^�����6Ru>R}~����~�C�k����o�T�/#�Q��\���h�;YvFl��ׇU�;N'��e�XѨ'+;
�w\"69��!��ξG�<}�^͘&ER��P����l�]�"���?�Mҷ��Y�i��E�Rx%A.$`��&ˋ|}�;���3=)�aQ�4 �g�2�<ѣ����h�7y�фD�>;������Zإ#�eg�oU,OBi���7��O��@�}�{�e5�H���4�#8�m��?�M �ĸ�s��y�����D�;�����ݛ�<�k)��㇢w2�Sq���c,c�i��0��{Ħ��O�?��*������i�� k��^����P��q�~k�5���)�-�dc[�2�\<=��Ag8Ƶ5*�܌����gOmLN+�� �k��n�nv�l��uwK�/PI�s��w��H��w��>䞚9*���ʞ�q��SL-�l��w��`��4�`������Ň�|)c�Q:Fx��dEoY�|X���e�?�xZ+��:1`*ϙ[�쥚�� v�W����Ȳ��s�mk��S�E�^3�f%_Hw�cu�{F�,w��f�~����iEi�!�/�}g���2�/�- �z ď�p����ٹ~�϶���Rf�M&�Tz��-yN��?��;:�~�Z��l�@O�t�0��K���>���a\�諹��L�a'h��s씜4��ۘ��\޳F0r�t/�Ӌ�c��w�P��ag�[�����- ��d���˸}��"慍eqM8�,7��j��T;B;~�똟��3�d�'�'���ԭ|�-��6[�������jZnb�6;O�$`����:�>�t�,��sY
��݋W����8�r��3u���,�}.������&�oFbC�h�CUa��f�TrR6����k��+�W�����n\^��f��8�!0d1��0����1�VFKc=����v٩K=}O����YM�r*�^����[!��=e�Ց��z9Q��hc�n��kz��n�rg-���Fو�P������;$�5+DHM���"�*R��s��g��B0�1̰E�k$"Z����8�����!#��i�* �HL@��g���h>Ð6H�����(���
%���DԌ\�<���Om��꺬�6��v�'��=�W|ph����y{�rj#ﳎ�Ҙ�(P���$�*�-��J���p<O颴}\ky��Y���X����N]�5vK���n7��+�r�R�&�$ә@-��1���*�Zj2V���4����ț~]7����	�3��q�+8K:F^�:tך���s��x�����Rн��ʢg�B�aC��A�< :�״2��7oЂ��!�B	��u3��,�����#�y�)�:�N�O��4Ne����di=o����.����*��A&,큛Qu��:�G��\��_pO�����XF�R�,����R�6���9����b����Q���+��4�b��٨�Q4��N?3�9L�+��cQ�����9��7c���m&�Mr��*1KZ?k4���6���B��2${�mFD��D���1G�������)}t��N\ޚ_�㷷cl�������-fw�����ˬ���!T0��F�[TNk0��>(}p����m;�-+H�t�_N0.ȀαVŻv"���4����/d���e�¥�3�����3��8Qej��\�O�R��n��?8��W;�&�G����;3��h�{�y��iԃ5�3�#V�X\Y�iUoU��ð��WP���0��*�q��`�٥:cGG Jg�W,����Ŭc5��fh�T��uÍ�L:G�T����F�9t�3'�G�:/)�>�f��FF��g���PF�
�Zw�c*i/6�R�9�E��F������y���yz؅�`t�ݭcM.b�����2w����:�t������O�:'8"�<�6�$�}�TԼ�����啛`]7�vJ��,s7ac ����Z�[1���~��T1r-��D{�[g�ډ�b�Uy��𲓇'37O�+E�����ͽ�3��\?v��ƀQ'r���N�`)|&@0>���a�/�ZޣO�����z�q*K�[����W!"Ã���U��9'Ge�'G͵ӹ�� !���p'ϐU�TvV:��:\!q;��Zz�u"<�ҠR�٧�u���u�� sOt��Q^����0�Ep�G]Yp9�'{&S�b�[r>"�^�����u�4V��=� �}�7KF��"�ϯ����^(�y��~Yܕd"���-�}d쎚��.S�A�b� !ABe)T��̹��F�o����r|	3�zhB��vbšOʜm�'�(����y%I�&YP�<�������O�������^���c��e��d.��t�$y������H��c��J5���3����yQg�d�-��Y/��ﶔ��`	��k�wr�?d��H��R*�*��D�����U�O�3ZiF�ĭ �OY���٭$�N���B�$�Pt�e���V�^�&`��xo�E5 ��eh�5�׸+Ȁ���wA�A�'���~,B��_�a�ZY��%$�'��A��0;�v$�Z���}�c�R�%]E�4���!�vS")�,	1)�=6_�.�}�a�8c�D�u���AD�A�:����� ��Ph��~az=�߆����!�RK�R�e�GN|���= �� vp:b��Ĥ�n�A�!Q��uħ|�O{�ԫ+螮�<9�+6��Y��^޳d��V��_�t���U1�a�g
1�z,'��&T��nl�Ё�mh�� [wI�E�U4���X-��:n�2�� ��2G����\>I`n����6�b����y�8���8k\A�y+&W����!��L	^�g�E�,�۔![��� ���O��@D�si�J5�w��C�����o����劵lgz� �Iw���B��^�AWJA1��.#-u*��~&.������[жYA�(;�ϑ]���j6�fSU�+sX��7�~�w�T���W;�=V��>5���=)��y+����ߗ8$��z�~`\T�&^�	&�׾�	#�L��SQ�F��Y1�����&��~/;v�ꏭ8p�[��=޽�����Szf����]կWv.�/RP#����"dm��fL_�,��H��M��ĽbI�{��饲�-Pt%��*;iM��"�Ld�!�W�[J��m�q��8�kam��{��<�<7�~5;4�2�{�Y���SI�;�Ek������1��CE�����0��T���ɻ�Ұ�M��l���Xψ-�����*f��@v#"�/��֤z�u���z�]l�g���h�d0��
�!�k�,I�k.Rp�u  �)��5��7� &�=U��J:S�zC�v��9���(����ݗ�S^���g��E@������f�����O\��a��q���ws?�V��ۗY����P����U�P&m�� �?tˇ��)���7���#�6s��%�;�\ǡ�B~��<��?�TtdS*��1�������
�b4o3��!�qX*SYS�uAY�Mg�(#�����?)I�p�zZ���C�"�Hvu�Lu޴����������5iBZ
�����:AFg'X��R�E�]��*V����J{�Bx�?��m2��Z���T����"���O�tM�u}���u3���&� ��쥗v��;���E?�ÚtCg5���JJ�Y�X�]r�FŌ���,�5�D��x�SA�����Qŝ��	6V�͗�G�U4���[A�6�8�z)�t�s�����Ef�'��v�b[����q��[W<���g��1@�"��o����pI?${�4X�Q����g-�T��M<п�;DE�}o��k�ȷlo0#�:����M�$k	"�2��D�rͪv>�˟!=�aq�T�b�����t��uk�#�_����\�H�����-̬��'��;
�e���:(ɒ�0���a���J�v�,	}�f��wݥo�?r��O�ʕ{��%�KNc��A�p��)�3_>_7���oȲG��z{��T"|Fx�Ҕ����XkS��#x�c�T>$0��)%v����vU�	�/��� ��S���H�e��!y�S&q�`�)���S\�����1BG�Ztrr��Q��T���ִ`w%�c�����
�҄M/Ih�Pg������ݚ�-b'XTlr�xk���;2�&���:HC3��ٖw�n9j��g2�L{O�M��t���T��#��Z�V��/ 8F�a���g�t�~"���[0y*�pkZ�
3YVL�{�uΈ�v'hc���|ـ�[b�B����=f1E��;�o4��:��!�G�!ųb���Q�|��^�2�����6?�������w�q��pd�zuj�ӌD�6�** �����=���,���K�@���%#@%E��%p�7pQ���:V��Q�:LE���'��� x�W����C!<���`��+�,ș�����.��_��9e:1H^��/��l�� 5I����A�n�,��媋�2HrS�yo�46�J���
�׌�F���V���`>B`�
HJ����ł��1w��K�8��!�e�]Co�'�{��&	��0���2]��*�;�#���Xl��6����z³�:�.���;�\1E̡�L��K'"����4��(>v�lM�[���U'�L0y�5�@G�̅'O⤖��� �C��焷}���f�z�Ĭ�Z��R��������p��]��'b�_�s���Mf|S��2P���з����X�u�4j��-���5�͊Ǚ�&�ͤ�E힄x�>
���!!�!�x3��:����q�^Ck�B5��$;-�ƙ$��5�Lx����̶�З�~��3���c-6�ƀ��-�F'�z��h�x����}5׳�L�GP�i_r\��w�D]�/�sC�g˚)�}�P�l��N?�^L��Fx]��1_��{L�<v�a�)"��V�)\(x��(��h���m�����H�Y���]E��ӊ6.��&L%�Gq
7��ǰ��i�P���8E^�R��Im��[E������o�Qc��q\�أ�i�=Dl�������ᮎ����@����L,�a�����~��i\�m�V�a�P79"Q6���GaC1~�j"��`���Ӎ (�t�S�zMU��kF���Ҩ�I�	{6u�爛s�t�kD�h�h�R2���M��vt����������=}���($:ˤG�n~�퀌�M�}��ݳ���&�4����J�Ъx�W�E�R�=��A����kE��;�u혛��C�p���jA#B�>�M���]�*���G;�'��̭�e�+���2���H�-���aa���SZ�x����+
�^��rg��ˎ�]�
t-)f-V�0z4��Yv�<Zm��U�9�����GW4؁�;�;}LZ��BAk r��me��d�6mM8k�y�n�`����ŮM�	\��RmG>F��6���Ig������O)Lhiǣ
l^�FM������hI�ٶD*{�r��5·�p�5V�\h� =,�/��a�s���(��m����r9N�)ɕ1�Fg�Π?�����K��~\F%�u��71 ��a��0�RK�j�Iٶ��N[��>k����.0�?D��g��h2�$K�]���w%�{J��k���$����$ΰ������&
\O�Ħ�@,Y��]�+�V���yrⶆh���k4a���YH���ţVGq��,��'�������L�����m�9}Ok�����n易���m�P�Q�U��DYy�,,�qZ�R��|�f�@�����J��,�o����/�/y�y�Y�	
��X�;E�ۤ��l�z%�׫\�����d9��e���
����5���{15�p��=Tӂ�Z�+���bq(~�S������& ��0fsE��Xi5��SN�ǃ�p�{�o	�^�Vo�I�l�7�G��@d�T^G���G��[���o���Z®�N�\�'b	U�����������w�8�,�q
U�D�^�[h|:0�� �.���e��1=H�Q���h�\)INX��i��o<�W����߿�O��Kd��W�zõ&�,��1;_+.�2���E�+�E�p�
N������YRVC���{��z7�8OKY!�i~�}���v���Gt1̓��)��Պ�2���x�'㻆�21���7�X��u�������L���р�^�8����┩�3O���瀨jS��ܤx�E�m�O�L����W��� ӥ�kL��5!؅m�����8��� ��vx�My�ֆ^d��� �|&���a>n[�ɥݥ���� 
�=J
��P3�h�{�4u�}�@������-��q�����ڽ5\-E�ż4=G�O]��-�F]/.�Ԑ�o߻�4�����--b_��m#���>�W$KZ1�`�9�a��d���n)��\7�h�N�k�ToR����%����]�G`��4(��i�����\W���e�=����G��-�������M�O���(����yH�dX��q����+��v�zk>��ŭ�2U���8q�\�n���@�q�oV=�;����rh��)��_�A�PC*�3x%���a`���<Y�
�K��o���2�iFI|9��_E�D	�㤲j�5o`�p��
"s�
�.|����.67j��{���}����e�%�� )Z N��� l����6X��=H��p�\��o����x�w|�
*�5t�^L2���4�օ����G��Ǚ6�'���d�Y�Csm>6	᚟�u�դ���O�\DO5�|k��^G�|��@9��D�䘳c�Cֈ������M�-�5�T
�k�z�.Ҕ ��a)KA���������� 2�/@�_+��BR�W�3��M��԰�"�ͩ�a��M���l�ӣea�����XV/�� 4P���0Q���
)κW�+OSe�*���v\>��!�����C,�PyC�y�l�i��R%�c��g5 ��oKO�XC����v��_��)�N)�ʍF�&ssV�JQURٮU{(\A�;��	'ɾ����4
�.�gn�W'��o����B��F?������6|�^5ެ�O����9����!��,`����kώOv!��h�4��{Kzx��$�X���nf�z~^J<w���)"��4�/�~�]�ˍH��j'A�eZ�t�0*k�n�7�ڿ5��4�n��?k-��n�t�Q��g8����"7��"Pč��{��9@���F��kf^���S>��֪7p�J�9����C-���޽�s���^l��ZJ3���p^��v��	�^O�Y�Uw��I�n:⌭-p�D�,�shf	VR�q�_	nʹ����y�揥�g�s���/�ƘFhJ�a���Ͽ|D/��5���h����l�e' 0M⪅����9�B:��-��&>�x�+6秀fԟu�T1��r�Ѩ����)�Ӕ��`TکԤBg�1ޮ����S�ӵ5G�i3Ը,�Z�/-8��S^n�w�Y��>��K!F��7e�+y��z�BK�Ht[�@�"�=U
[M�66:���K�}��})Ϟ<�0q�r�]��[�V5��� tN@�kX�[�U�����f֤5	xE��*�Q��ȣ�V��?b�=D�y�T�����I��xX�N
BV�q��1���b,_C�-�^�N�v�Q�}�cMgn� ���6��63C4�@�6n�%:r'���[�v���^.��4�]@<V���`v�*0:��������pa�7���'�%q�B;>�2I�����E�&c`_2�ʸ��u\CM��T�z`�M�
J0�`��`�g�:����(���_�亞^$�'P:�hd�3ޭ���:��G���2l�/%DĻ_�� YdY�q��T,��T�c�mD$��Qt���]�����==�*��l�c'F"���Ը6�#������{+��&,�z5sX�XJH�T���Eqpс�{�j�+�HG��k]5�3d�'ޖ8��!�q��wٿ�F�P�y*2�Gd�+�[�X��T7#M�Z�Ւ��
#���L���ũ��/}�<K�a�Qd�T ΋��0̼9�:&sm+�ݚ��9���Τ�<إ��0����o�[���k�V?��a�~Ki�'.�S��33%����� �Z���$�X���A�f<��)�v�] M>+}�!s��Ig����Mf��S����Ye.���E�v鯀������'�ה�vG|HXKR��m#B��Ev.F��^�2Z5��vcY��h�6���׌W���+_��:Ϻ>��z��@��] ����z���@1#g�`��]�p
Ke���9�זw,$ ����5AS�4i�!�ߟ� ��m��x.`�
>�1�R�xu�8^�poù̳��;��l�| d������B9mʇ�n�;{4O� =p���hp���𪊬�E��G��hyL��cL�|���(�'li�S�ڨ����*�H�1T���a���;�X�Uy9�9����+�5��6��i�Y�r�7�!�ȩ��}f{/�^���M�P�ȑ&��WГ\��׭��-#�:/�ʬ���G��1i����D����1s ,i�b�
���i�{�K,0��Mk���z-���H_tu7,h�J4A�@��)��zy���?���Q�E��2AQ]"� n�=M��������Jж�ϫ3i�"΅�+�h��_!=��~l�Y����z���:���)�d����mDhuN�<Nt�	�;�PE��%+�dd
b>1�� �h���T":GG졸~�
R�X��S���Lò7���dT�
4D8[�+|NɆA]x63�)=k%~y��$Q�hi�^���fč,��B�q�o�Cs�ujN09��� g����IA�3A�~�sM{}�cc���myS���5��䋪+���g�t�Q�5OƠ��������V$*"�����HS�{�[��7A�Zǟ?j��q^��Ⱥ�mi���J�kd9ϙij��-Ң�gge����U.7�>bX���ݥ5f����&ߵ����=�S0eኛ�v��B�ث���U q,2��-]�@�pTT0#|1�+���f�=��GI?u�/��X��T�{a/�ă5[͒��"�;@��DL�J���$e�p��D�#Q$W��U��8ҩIrKx���DNO��ĿD[���Z˷_m���iI%q�_i"�Gb6}ꖡ�[>��A�QΒI5=_ۋ	��7d9�_[�8/���Mb5ƭ�2+����W��-8;.���i�O=�:���	�T��YB9q��-�)��݆r5���5�Ŋ�5x�1���q��Q� �4����O��Y88�(��<�~��Ky�e��[1T��v7��e�_l�7��c��0�C�i[�����W`�})��eC����`���G�'�ɹ�Τ�iXe�"[��}Se0L�Ĳ��Ro|Sf�{:��G.�娓Fݕ���tM�˷��q븐�߯�pR��С�X;�&;��-�aí̊0�4T+F��� ���xg�<����bw��Ҹ�(TN0���}od��n���J�bV�f�3�k�*�[{�_	�Lj�ig�@�|{�rsn=�w�]D��z�v9k�D�fNcz���$��wx�d>���I���}iT��@��˪�[7��L�����o�����Q��=�=I��3ߊVfa�C0?U�M�� �7ȫ�b��6ԋtG0�x
�L����>�����
��'}�hV�fН�2_7{��\'P��e�������bBҠ1]b.�C��(,F�)�l����t=��>T�����ɯ��#jub�Y�g�@X�������g{�L��?#p������ּ^�=N!A@Mo>��ka��#4�Կž����1���׎Z�b����A[�wy������IH��;B�B��E��;�ꢡ��G�ď��t8��1;P�m'��`��9�J��A&0I'�*�N�[L���[�)u)�]w0F����ㄙk+t"�����Q��8��	�� �{�������m�E��n�·s#q��(����N��Q����G��P���q5�m�/�
����ˣ���\]7.r��n0�RC{�'�h�p��^�{�+��~{R^;t�R����gR���D��a�D^\~�~�Ng��"���<��'G�*�α~1M�A;��-���U�m<K�| 8@UH�3s�_�@"3�^�!�]so�k�]����}�z̯ʺ�xuHwe�h'f������0�&H�Cr)�\�� �'��0�t$AR��(�VK���ť���7 �A�	�8�W�`�M̼��� �TX˚iNQ �hq��v������6U�߽��3�X\��ߥ~�]�p�u�Ȼ�a�_�����<7j�ɖ�t��
ޣc~HuieC.<�06Cj�T����q��N�
t5�'��P1��A��m�)�O����bo�ç$����R���ni^}-����e�8X��f��8\�ڳ�?��̢Xx	M�q�{�noڊY2��,1�uNr��\�j��C�B���V��Gjl���ϟ��م.#&�y��vp|�;�m`��N;>�u���)��D��!��<���_�goo&�"��Ú���e���8ċhp
ط]�q�ҟqѾ��^���9F���\��GOp�1Fo�r9� �k��H}�����I6�>�9W&���q�	��|WF��)��$} �TS�B�u�ܚ����Fj�r�G7WgV	y�"�Ut^{|��nX~.�YC��V0$m���*Sn��|��b)��ӝ�m�X]�L����!-��7�>���	����[��D�na~�E i'.V��mO���Ll$����8���mj������}���0Ja��{yjA\§�%�n.��혎�vXq����h���"�bI�YZ�|!)�2�&dЍ�K�k7��!w��Ǫ�{��М�P��p��9��žͭ���w�2�|��{��)+�=d2�W"��N�� �DyH��^J�u����
r���*���DO��OHgi����%'h$�u�����-�*hAY�]]T���l��jNɦ�d�5}v��-]�\�+�6{���;�;U5?��QS����p���,У�-�T�k�K+�ě�W��-�7W�A�'9�'��oW=�������qG��b_f�6����:1�t?�d�DY��iC����N`c��Y���a�hfjD�� �Z�n�e�-ʛB\�����1Hqd���!j�bFEA�O�8K��7��T���d�7�`�����1+�X4��f͇5�4��n¼�gG�`R�!rdުFfa��������vb���s��bTO���
� jYQ�5��$�[*�������]��>m��^�A��
�L�)@��[�^0W�����5����[m�Q�u�ӧ�ûjP�|ߎ��@�/���"��6*rW��� d�_�(�ޭ�%�(_��)^
b!Uc�Y��(g�Ԋ�JH�1��p���(�63�M����&S@�����s�t���!�f��̉�L�L-��w�]j@C�4ڐ�g��p�n�9��K�J�Z4l���� �du�xt!�Ԋ �u��l��+��&$�!���2���nJIfeJ�� [{Qb��O�����H�{"f�i��Oy�L
{ 4c՞���f����S�^YՑJN�@U��t�����ke��B8*.[�j��l�e�O�g.�Sk�A����i��W��D�0�=�66-v_e�V(S��m
�ϥž.4�y:��[)��������J�I����H'��,Eѻ7̉�r�#g��Y��$���;/��f9�
��������ƌ���sE�I6A[vڈ�ph�8�Yy��~pDÓ�#����v&���(�d���[�?��6쫯g�#	sd�!�y@�$��,���*r� -����[0��$g�Nd��#�#`�۰�s� �h�$C}}ӝ���,٣}p3�N��E���<�n��I����=.b4{}� �N�Z��jv��~0���87�[��AA�S�li��n_KJzgg����A�:8I�֯�E�r�ދ�^���2,_C�$�D�g�dFNlڄ=����Fse�͡�_��bw��6)�Ts*:����w�I�y��\�ר�b���"Gf'm<�|�Ƚ#��_���=��X{t��F���Τ_�Vgx�����X�35�DkZg�fX��6iK��n��E�� ��w�)�������;㳳7Mk7Eiz[$Hb�r�>��k`\
���d�KT����Ydҿ�ڼ�#t�W�W ���Z���<#����3�cQ5
���i�Π��ռ(T�ۺ����\��
t���Ëx��w%?�[����K�+s�.�a��.��X9#�x%�5?Kf��s&q0Ch.���y`"s�,,�f8���(X��ov��IK��p羹����D\�F��W =�װ��c;��l2�Kxy׭{*, ��� �5���(vZ�����<z��ZC��N��:�E0K�|ic�1�N��伆]�q�
�$��TT��B�f�?G�6N^��+��6��#�W�')=�be�mL�����١�x��)Nt�F~e��/�Hъ�<�Y��A����%KB�w��b��N���{�*|��`V������4�pYt��T�̘���TRT�=�\�Xɥ�d�D��z��ߐ�3�#4
x�۠{|w��D�ݤU`�DG��xlJ���~�`���1���(��� J�$)���>�`���z��k�_�n8�1���Z~�����X5ȴ�.��VB���|T��q|��e��40�'�^dlc�j$�����9�[M�V��3yu�W U�����Ū����2t�[�Q�?~ｭz'ѩ�OM��1kH���|z��F.U7�9���ʷ�2:kP�l=�az֪��K�! �jS��tb�}��Q�2�
���Z傃=E��7�=�hT	�Ry��0�" 9�[��a��Q�[y�!���{�~�̺�Ll�h�hYʶ���6��\ytqͮ����4?����]�P���<���۟��Ŗ��M7i��j���op����PX�="}��l깈�2�2�|N�Db4,�3w� �}���R���'�'�(�Q<1�;��q�N��c��Qf���y5.���td�g���dɃ|�e�����j���Z��<g�x������yb�.E~��������%�2(�D��.!?����lA�Hm�[3�K�����S����Uw�':�]Jɴ�m��r��LiE��)s�
���5�CBz;e�}��3�L� �j�bY�5	�E�L��މ>���.��p����-%Š���ð�VA�M��N�S�Lz��{'SK�_�:��F����dC��1g�Ɋ�O���S�Y��ޢ[�U��g�]s��EQ�T�ˆuu}��{�/��t��u�a���L�ؠ�����"�J�)/��;T�s=w��?n�o�5���۶���qG��k &�����}�@�%#>;��!�kA\4ӟ`���W�g��G�^ff[����,Uu��G�{���Bxs�O%
�rs2�2�8�B�'��D�m���c���t�ϋܗ�H���[�鿐��h����Ò�{�5^ Y���c�� {&�[\���l��d���+��ߖ��Y��?���K�Nn�>�����Y�l���X?lvAJ%0�vl����y��rO�����.,�nkkͼ���Ge��)Z���J݄{���p����5�hbw��S�a~��-�<�K��}��a��z�
�k���_�T| HA��E�����Ԛ2a�F���7�E)��l�V,>	@� �x�­�Tߘ�2��h�*��a�V!e��O��_v7��Z=�6Z�{ �Y�����57������؎�♘��M��
��W��>����(K#"$|�@_kh\��@�񂸀Uzv?�G}*6@���4���&�2A�\���V������	�KO
2�&��9����잧���N���JFr��F%i�o�?l�����/j�΃Wt�
2R�U���Ú��j�PA�w�$��D�d������F�|�SDd3F*~:< �]�+ d��P{#����9�>=��R 6��\���,'>�E��w�)���}��4����N�������d��G2Z��c'�C�MI�=xO��}�猩4@�%<�/��$S-��̌80�Y���eu@��ƪs�-�E%�iL��e+:h�s"��k?����oH�fT�^���l��M���gĉ�SCu��%�~[�}Z/�#����0�u�w�Uc��v��Ɂ[���3}��� U΄"\�(1>�Q��������U�nJ�I��
��}Ӟ$�Yw²9	|6 �b��w+���̴�D3o�:wD�j^��5���が�o��%�z�ŬW6��� 9���lrr�~���!T�7�MR��	 ���?�T.BHEU�,�7���f�U1���6�Qu+��v�Tk� �Hްw�����G� ���F��.��t��j�~y�\Teu�Q�qx�O�45�}�����ӻ���u�j��5�:��m��l�5qD��ի��:;s.ަ�ޮ�dN�.��Ft|)�a�=�}�B`4c���ɾD�/ �m<��R����75�$�}Y+j>���H)JB�2X�>Rgf������.���RE�KͭVKD�R��/z�f���K26�E������Q�K�t).)igU���{^j�?/�Io��IU
�\X�N=@W�:�>�X���ȊG(��Ð��q��Ndϊ|q|E	�
>�M�����Y�`R�/d�tȧ�S��s��r�5]f�P�=�f.Yz�q�������6\�ZI������bj�����-��	`����j���Ǌ,㟈:��� h�Sk��������j�"�e8G*�Lz�/���\C?
�r9�Gk�P":�_�ż >xn�h��h�#��_�n��i�k��$̈�BC�7�����-	�H���"�����>�h1�@u�;�r� �-c<��je��T�"��fǛ
^͕n�MO�F�nB���T詋�ܞB�h�B���j��ۂ	��%���΂�f�j|%|3�`�G�GV%7�Ɲ�����f?�e�*��e�ֲi{����K�b��P�D�U�)��ơm8�t�����Fv=�Z�Mlb8���� ��1��	� ~o�A�5́7�u�� ,ӗx?�'�%Ga%	RBv�?�!� .�:K�����2��)erY,�~LDE��H�c��@�^��X��׿�c� ��(��;L{��@� 2��_˅
E:}�'V���b��
m��m[� +o䛵)[6��(���V.�{`�x��z�YM�'�@z������h>b� 
�wcqĪ���y�&dĻm��x�[�7ƒ����5� q��2vl�#���,���\5N+h����r\��0����>�\B��@� �R BQV�	��^�h&�9
V��%l|3�.v��z����)�X3�?�miS��F1�0[��@����a���kH���̰���䖘��z��&U�%�0�����p|BĜ��F�%��2d:4O#m�dZ>��I���(�C_D��V��F�h�_>��Y$���7ed I5�R��`�w;�1�A>�/c
�.%Rϔ8+>�r)���¾��ª8)���>8�<\or 턙�%�uH���'=�*�`��C���m�T�q:�,��2��.�5���{��_XҴU��b��W��r{q�9|�)w
w�*bҥY�;Y[��-�j����:Qp��>��T��ю����Mr�z����J:x֢��[����u���45K轮�D�_�7+
	Cu1�yi�׃i�b���/�W�n�6���䥵O��a�>��0s�{è$j	pɻ�_pfDGFg��s��K��tSN_����@ �V-�w�+�ݚi)�7F�nx�\0^;a��DVj�?�Mp��")Ko��x�t�Bj�5�f]�����6�X�*��(1ҦM��嶔�Q�/�@F_�%�Kbvd�z����?��_�"�*%�Y�g�%���B���Q�ø=w�"�C�c����Ry�s�n�rl�i,�>��fh8��B��=(*��p��0�Bg�t����j��4�q�H
������kW���s͝�t6�Z	���G��=#!��\�19,�r�!z��0%�.m�v�!fs-l�H\�D���k�4�E�P�����ݺr�@�ُ$�C�n*��I{�*v��	��N�٠R�W��QƊ>�v����Qj�]P�5�ۏ�l?B�jV���� �5����}ŸV]|_�2�W�ar��w�L�"�G`'W� F.����e�1+ŗ���#r��h?iЉ��lJ�)>�āN� r�k�⿘bH��M��[�uPZg��,����m�N0Լɭ賎��~���a��{�K�1<@�G �ӋB���� �F��T�HI\�^�SQ��bryW�����'U�;e抸�E�p1�1�K}] ���bq�N�2�e@�@J�o$w^p��r�m0���p��%���2��L�E��=GܗsB#����:7g��_��M�c���,-C�,������)c&yw�j5�K�Q�H���a#�ছ�ؘ�����'�D�O��
e�r����������EG�$�i'>d�E�k�o8T����%�c@�4���S��=��������j�/�6y�SL���X>#mn��r�Zw��$t��E@ =���QD��?[��$��3}�5���*�)�j�"�L_w��WZM�B'�����s��j鬺תҢ�H��k4����r�	?��7[N٫Ƥ���aq�?�9!)c�Y��K=c�m�Y�<�����j���� �yzI0jJ).�����.F'�r�H��Z�[��CC�x働��܄������`�׆^���m�uw�q""��,��(%�Z�Q̤�y>.��b��]��˧@����B l�åC�(P`��曔�g�+xVy�(�34�#�,8�M@Ie�BR�pf�鵬�#��_i
�B��*�k�g��v�~Y�2����:�5f���ũ��b����ē�-
��Tx����}�g��N�Fc�h���&3 /[��Ζ���?��P�*����eڟ뜜(f+�0���B�g'��=E�c!~L=s�h� �mŖ�ki�;�i%�]�O������p���,/��,e��Y��[�r{3{˧³�:U(G���$��HR�Ov��YzW����w�^����(9���b$ʥ�e$���cJx?]��~��y,��}�b�HEt��p9�yE��\o���f���9�39y����2�دFbǖ����n��3~ >�h|�u�>�w�p�|��"_��Q�L����ȍnV��zE�qc�@�*ԗ�	K��I;y�98��X
���жڶ��t�kUU��\�o�1��@����[��OW�}�e@̓�l�D�
�ҹ����.��m��Oi��8��7z	��V%'x"�Z�1gR��]˚Uct@�e��jxA��5�8��oK�>Q`����2?T�M
Tl�kw�A��n�dfT�
�*<x۔�<��oxP�Z�| ~�#3�6}O�(�6��z��uJ�*��)!#�Ki'
31�����=�����7��co���v%J<�oE�ŏ�.s2���D*�p�*_.�Qڈ{��TŪ�� �]>���L�˺/�����Qt���سu�3���Q�j6!� ED��z���>�<���=��WpT	����-K��f~��"��+8�p���c�0uHWb'v���M�C=]����M4���L�u�g~����w-�x�T��vݙdά�4�Я���@���ը��@�7ǸB-m�)>G%j�	^��#A�H�x�ȣ}7�}�����pr}������53���������i)�ֺD�SB]*8:_��t �{"m��"�Ȩ.�p�@e� ��Rc�*�}a��cL����L#qy0�j���Km����5��h~"q��!^9V���2���O)��S��i:ΟO��L�,jLv�)�ט�dB*V�O3M��-%�Ia�nc�d#m`3�*�St>����#+a�"�b��/���yO�%����d�u��T!!���9EƆ��.��ʤ�K\��Ub��%��ԏ�����q�+K��!��
��}����e�
5�m"�Xu#�y�7�2�(cc���tZ7��g�����|�h� �/�T&�.o�]uo���8�̭ߊ󗮋��)�C��\GN����]��CLAЉ�=̦2h"(93ʄy�%&�dF�=�Q_spB�ȼ������;�����d���d7�42U�Xʌ�����`�&�:�0�b���n(��|;�_r��v�]��)�#m�&�P�U�>��O��	\E�^#�޶eE����HK�*�7H���y�~�
�a�+C���v�G��C���U}`��z!��3���Jn,�ܨڊ%6��IR�[�ts�J��������˺�(�:�7���#���<Ebn'-�o��t�Z�f�']����0�^Ke:�����\9}L�׏�`p�[`������ե"�k�l�&���
�K$ut�5�� �� �5�!�TԆǴ"�"ß��CS���9"�Vy߿i6>E�s׀�Ӻ���<��L<�� ��.�Q�4��
��օs]�����mjy�tthۧF?RdV*��J���҉"՟ӗ@p('��F��,q2�K�C��MS5`V�nNMyll��3`!rkO\
a���!�r�A�c;��o�E V{�
6�)�{� �z��+��hL��%��͚�D2#���q|�k���i$!�g�P�����eq7:��rr�ӄ����C�gn���c�����>�(y�� �%�kb5m�í�%�LXò�[4���� &3��Yk؊�~����s�&��<cc	
��?DzTLxi��ZbI�0{wh�W5�N��hE@Kt�(��d������A�jJ��5�;�h.L�(a�@wD%)���b�B�[Ȋ�^��s7�92����:��r�ޒ����ҳ��e֡_9��߽f��3u&v�.+��[��o��O,���qG_E�t2]��Pk��7�-���Ӻ&� v�z6W��������q�X���v�#���~M�d�k\/����摅4-�򘽚ߎ!9��g���W���3qbmd�����魒Y��
��+ǯ�Of%36��ƀ��3�?�]j)��e�j� �ڧb�ߨ�6�פ
k��{Z��c(3�MV��f阡����0_{p^=ye?��E7Qaխ����7n߰����vGF>��Ր>� 7�ő'(�����H��>uǑ7�s&�0$��K�T��&�k�W~s<��$���n	c���M#�h#-�u���` �Յ�_r����|�פq�/�,�If-o�/��$W��%�s��Hδ�4L��A�
�U��k���k*����Hs�P^�S�n1�bo�@T����4���Z����tK�Ū�>E8"��jF�+o�9e�ӧ���&"z)\�%#Z�d�.Z����׿�X�&|u�~r�L��#R;'X�Z��<1�&�;+լ���Z��]��p7��G������m�QL�*c�6l����^�^�i<��2�$�v��zwH��$5��'�O.׊Ĉ$����>/Y7�u��/�_k�5o��?Kg�Kjk+�"�[������=d��pPN2{ǩ�if�\��aR WF@%�[-���Sq,�j��$ݔX�������J)��ܹ�!���K���6J���"�9X�ڴ�(�a���Ə���s�1�S�iQ"?��<��Y���V��{���ahG_ݮ�Z�c���>J��/;
9�g㮾���D�{3������'���s���A�8T���k���)+D~�ݦ>���������GY�v�/rqs���-9���U�bg���$1Ȧ���裂1���xb�v)os� �>Bs���/]n��5�I��y��efv��IG�`Y(7��K�I�m: U���WX2��sp(\Ee���ю��r�S���"C��o[�w��?_�̞>���r�g�2���v����1�g��zܵ T�f�#מdk��6�ͺ��n��FM4h���OJP2}��
P=/ �����w�O@:.jUw^'�zbr�ݢVVk��}<�C3B��ƫ�H��$>���0����v�"V�
�A��7¨��q��z�.Y���m�W�	��I����튧�|�_�=��]��CE�����)Z��*������%����L�(����dT-��}�Sj(`��/</��F�(u����S�˖<,��Z��$_o�W��"1i|�$�p*�I�F����u[�Z��'��J����ٱ�ik��VH׾[H"f���������V��KG�Q���G���H_\���kI�y��3*���-}��*�قR�lb0>�C�K��%�>9�在���g��g��#Pg7�L�N����]���8;�;�9}#�n��_�����2���P1����}M���m��J5a�M��B�[v\�h&2�l�%����	"�y�7ݥ4���.�^��BP3w�ݭ�d��u�óv*���lbL���@�p%��� ,�� 7���`��Y�V>@���^���Z;t��(KUo��@rFa�mK���˕��=��I��9q#t���V��3�D�^��~�'\���w�>(��F��;�+n�̳��҆M��� [O�RUl2
�9�U)Tm;aQ��v�t*�^9�.��mb0X�^ч�+��L�蓹ۻ5�5,\���E;>�Z����-���4���5u�+�M��i��^���������T�1'�S�x����㘗��atuuh���Sa��f%�_���h�QWW�y����ӯȿ�);� ����Tl+�z���f�^��GޢZV��osf&$�i�
Ck|��ǖp���ܽW�$�6�H��K�c�/�ޫ�������*ۉi���0�QuL�k��n ��<�
�g�,T-t���K�U�\#\�xx�x�'����1w^�(��G})����`Kt�w%0�%��hE���PKj*�dx�S����,Rp�0�R֗Ii	���6bs��n���#�N]��?%�-_����5k2J�bT����c��jfY�^���;��_'(�7Pݸ�ǲk�u������^��S�&�mBܣ.J}��C?b��1������9䁞��I�P�}�<�H��w(��tB�r6j"�I��:�����KW�T�ZBf��e�@jYQ�J�l(\)Jy�iZ9��C�oJ�ǲ㒖�巋l�h��X����񁏦݃��o�B���w���9H���˄����v^�aj�/,�Ƽ|ЀX�R���� <�TJ�?�=F�5�`��<�Qy�d�V�.�J����7|�w���y�2�\�z����$�N��B�,�O~����ɕ%�E�t�Ϛ
�;:	քF�R�g�'|]�7�r��N@�,$�������M�~L�(�7�ٛ��S3��Ƞt��H�j�	y�Z�������駇����c�s���h�c5�j�3j�Щa�h��a�
����.�wrV�H�֕6@e�v�uA��f�=�oc|#T���d���o� �yvΔf��
ͳ�Rv��sH:ł�{RW�q��z�dF.�!UqU�5���)���m����7K ��Q�孼����M�o�D�<�L�]���-�E�u!E��ћ��Q&������&�_�_��X��/"E�f��,��M��8��V.���V�Jt�b=1�^3�>��Ϯ�j,��!�� '��t�i���ZU���d�g� S�2R*Q��Ѓm����BO�#>m�t54F��c�&4A)", ��q�?x)H������Ő�o��|ΰl�!,���������v,�"+�0������� �at^p�<�a�Z�i��6BuNΐ}'��˂����v�Ky�_/��;���p"�Ј	�L� �)7(�e0�<����z�ƕ���y����ߞQ���:1���}^8����}4�PF���^�7�$.�����v�jX{i�ɳk���� 
箊��\$#�A��q�H�1�G63�
;�f����˙���F�@�d"�g��ƻB�!zh%�����)e�����}# �-f�u��z�>�K��4�P�$\�t��ܯ�=~q�"`	�S�v(������c��W�3���ot'�u�F�Ʒ`4�i~������-=�;�]�� �Fn������Q�I	�!���ML`� �+F��r�'����U���M�4�ߓ�d)��Eī�����65�]�-M�c�ja�[�U�zU�	����l��<S��d첉�v��uܟE,H���gv��cW|�N�<��cT���P.x����9zHt�>n��U;ձ��mb��-mE%��Z��3m�������*F$�p�v��|���Ʉ�p�Z��X����z�W11R���R��wZ~���$�E{��0����I�6�R.����@e��Un��Y^���h��$1VF0�-O��Ƨ��?�������(w��������[M��zh��O۵��a���JP������g�� 8�PƌvcwL�@Ei�y��R��JQq���>�h ��O�>���#s|g��)\~g�;}�����-[O�5���S�Q�&��2/)! ��Y݆żY�����.Q�QT��0��K{��W����6���P�̅d@�9s��^P�l1\��Tח�k"�@oP9?��/��7	l(Iz����8(ҧ����S��ՃL���!�~F��L�A����/->uM �#����)��vE5+��d+���wD�j$ �z]���X��X�#�eFH��rr�u\H?��6()[�ft���� �̝c��5����I��"��.�8��%�F�[7G�>�D�zSBpJ�����S�g��Q/����-'��.���6htm���k�
��9>�6Z:�f ��"��a-�EH6�_��r�_��E>)X@�X	59/oY7#l�;27�q��cF6z=4�����>\�{�W�����Ȁ7"?�ғLX�R�@T|B��w�M�D�f*�>e��8��s�熠�U��v	R'��+-/YI�EO6�'��qa����0���Nj%]�o��?���t6[Y�9E��ռ8�]�l^h��a����s2����JP?Cts���EE}Q·.JDs��
|l׍�ݗ�p;���/nsD�i�����#]����({׬N�Vd>Hțm1�14_���2�.�<������1�L&��5ܯ騒(-]
���(�o*W���`���y��],��Si��wj+r��R3��p< ��%@��.�u`tՏ�k��&�2-���W��ug�����t�硠��ɯ�,�-���L؊XlƖH˩f0�ɲǇ��ޕY	>zg�Ü��j��<�ҙ]G&s/�>��&aE�U��9D�u���>$d�4�R�ƹl-��#�xA��$�v�Z�� 4QC1rFg��.6c 쭹��.��a՜KG!�Vlެ��B�
�Ǔ�L7�gX������}4.cj������!,Q3�L��猤���y����zy;C��E{7?�|S�F���u�b���p[?=�u�u˂��P,��j����'�1$l�X>g .��X �<E�+=��Ufè��`Й�o�X.��s+��l�[i�.ظ ���ƣG�����	ǃRRDAN��m�g��,�� �rZ R\e�܏���]MI*�Q��_	�g��������I6lڇ���[W�sq�L��_=�g^\':\J�5;�PK�uX�2΀��>�&�����1����@u	��&�5=.e��uJ&������6�!�SZ ���Pdt�l�p���&�c�'n���IT�U�LoPt�f7�}vJ�j@M7(���t����U���پj�%u����5r:�>�y�5�&���/�	=���(���h;��"8�ACP^#���
�V����O]<�N�n���E{IcN�%�rܘ�9�d�~0S��Qǚ����E�T?��"�w���z��<��=������$c����������=C���#q]��-��Pȕlb�=����Ԃ�\��%�ɝ�5�舶��_���6R)����{��.��2p�>p+���G�!�*:M�*~GC�$�(�0�	� �T��]{��a����ąh\Iôf�8/�7h���"�U��F�D��z;��D�7<n��S�L�G�(�q n�맰���~���U���(ez9'D"M_5�Y^X���U�̢�׶��.�]��֭�es�iՃȩ�E�����b9�֯
�!n�JRK]��҅� >�0�vv~.�`9#*bg���	��CՌ+&u��Z�q��xU څ�Y�3���%r��j���� 10J�@a�My��2��N�ٜ�2��@*ct�M$~Z�����JV��lf�Pݦ��A�pot����I�*/�����yY�����������$u��Sk^ʤ1�;�V�"-cx�4�,$�1�0C�+U�ƚ�rf-=t�H`KZH���Z�7��/�C��ˌ!�c��n����_�@�4$x�/�YY/L��˨�>VPV�Ǭ+��xs��ʴ�2�B�z��4�=zw��8@ݝJ4vbzOuύ�q4���)�D����ma(�#"��,Il*	�:S��\��Z���r䜖*W�/9�o�.|����^p��ȵ�,O���(�����.e_:RU�	���c�s�hރ�z�-�1k�}?mw�7�۩����Ȟ�a�
5�Ƹ{�����
S��'c����jLp����+�LS"���z�hvM&r���Ȗ��W�=�n��n��\ѶK;���_�a��K@�]��"�|��'��h�.صq���s�:\�����4V.v���yy��g�����nԐ�Z��D�*����@C �) �#�f�"�)��r��>�Yo�r\��I�6�d�B�w$=w�d�`�qi�t���NQJ��ڧ�o3r��2�c�}\W�mڥ0�+J�Oɩ�?Th��ۿ@����4�SI�C&�����,(�`D`��S�̗P�E����-�qͫ���|�O_���z̓A�'Uɢ�d��c�E(��Y}E��t�![4J �L�O��ZVZ�#`��{�²C�þ0A�e�toԲ1a���&O�&�wl]������L��Z�[7� @����z��~埳gih����Aƽ��e`�WkgZY�!9�X�Y�����VP8�D��~�f�%=y՝�GN�I���.�>��Y�e�����ϗ�����V��+��H�;�?�K���N�~ŭ{,ю�k�~P;�v��TI.m=�$��.��&�����Z���̓�֞�D���Z\��)�*,��Ä��>�k�7��+�o~Ȍ��L4�m���ec[�[�cr��DM+
`52�����f����I���s�
I	��U�ih��c�ʴ�Q������1��j�R��ξB�^)w��e�ANbP�Y�F�0-� ϻH+�+�HA�=]�n���M�#AV
x����V���`�EaHu���|�}2�e��-U������}�����@A?���Y[43@J����b�Y�h_�H�,�eN��X��/s�ٹ�>��7C�{o:_v:Z��GU�Z�,�(/�W���ǲ@�2U}5�l���=��zi[��Ld��J���Ӵ�l�J�uB�����W@�e����r��f�mx_�]Bԕ;�}�Y��*���K�1�n
����K>-\�ܧG�=s�V�(�~�<{{������qԶ%�*Ln���.m�@�\S(���P^P��}n���-�Q\d\̺aXo�]�>��u���WԦ�s���'�m���栚���氮���W'MU���CթW|mq��׋�Bi.�TS�����Z4��[.D$���$�y��)^� d|@"��">s��.�;��r��\V~7Y(��Ϣ��5>����[��������YF��݉��)ˢ���{E%�ЦN&�S,v�C�
I6M��@�~�E���o��8�i�j��N�-�͝6��
"��s�jc�E��+���O���{b�0��X8TIQ��Y� �����"��`Jp�����daX}/���O�HKgV�F��8��ں�>�ߙ?3͈���w��Q���Ӵ�<��V����u����(�0ӻ��>���sMoh����������u�;� <6�� �»q��N1�m��O���p�� ��&4��W�������N"�t�x���4a#�t4�������5�U!���t��4R��Ȣ�����i���O�r��v�q�Vv�R��-V�=`n&��'�!�M�C���ۻi�<�>>vk^����6�C���]�-O��ȤӹO�a4/]�sx��HP�۝�c���q2 �����$�
��;/o�c��w�@+��h���"z�X����2��.g	:MK
�p*��]Rm�#�<�]���@��l�>�\B���횞9{��ـ;��h\�]9�'r����!֡����?����N%�j#����2��b\�C��u�R���O�D+��jXn�w�.��ߊ�V_���D~�,ޗ,����7���ƯL�%CP��s�����ߘ���@q�3��:��@ܡ��l��pC����r�BDf���	��Ӊ0��dUg�1�a�.O	?Um*����6B��࢙�ؿX["e�6ީ.Z���8�����xO��+P�7\Uî�m��#�D��(S�Ո���M���r0<���iRԪ�]�&�ƗEi65�8uâ�ّS��-��L��xg)�
)��Q].^&�΁�Z7(��u�88�͝���/x�k=��y�s"���>&8R;M��7(������_v�f̖M&
E2�	li��Y�Į�"`���^һ�(����rv��m|��S�F��z���x�DQ?wx1 �P�ֆT!��Ҕb�k��A�x�I�v|��ε�\Ɖ5����c��0Y�7e�`yvq�#��>�V����@hS]��0�5$@3+xa��3��H\�X�����&��.:z!N|~�Tj�Q^cmDq{��^�In��Gbcn�t�"\��R=Gd9��ҹG����+5�-Ӄ&��n��%��&�Q�٠P/Zg �G9��U�5E"7��9��!��M!%�Ӣ{���S@4�bW�7�`=rѱG��#��=�wԇy�:�N���A(5=p7�g�?5��C���8����.�*sY3�[�e�o�٦�Ne8�뜼��ȼt��kb���V��5@fR�1x]
L"!#��:�����<��Nu�@%�4mR�?�S%;�D�@։dmz�4=��
ȇ��R]�L����Qb��B��F0��W<4�G�S�f���i��B�5VP�b^� �A�Q\�6�WC�Qe�VGT����-�t���ųn�Z�T�%�k��!��b1�;"1򅌮g��X��Bڟrť#����i�G��I�N�H*܍2T���f%����C�M��w�7�7UXg���ix��+���yAk���+`⁸���W��-*��y(xC��i��ܵ,aq��zM��ue� �U�ؒ/`k�ۑ��/?�d�5�����
#-uq��`	���<��	����V�U
zI�zF[��y�s�b�.��r�=�Dk��ƅ� ԍu�qd.��R��*�v^VA19���� ��5A��X��G`��!�O�,CS�'��l�3��&UJ}g��`��<���� ��%��]�տ{d���ү)�D�����5UI �6O�mؕ}�c�Rx�r���_��t85>>��D�t���r�9r��
��v=f�#Ѝ��Ŭk��=��ꎜ	��
��� 9^�҄�� V�. ܘ�X5�jn{�pO �Ԥ0��G����� ���!�b��e���5�I�V s]�~c�ZѴ�Ծ<}�_ð1�`͝����$5i��tC �CO�'�F� �^r^�����/�~�
�0y��?��=u��~a�e�k��M��cc0����.	
�D�������_R��ml���	o�3�A�`����T'��e�b��`�X�cb�����T)	��'y/��j�^Ν�O�N\:����F�.�$t���0=�~�O�t�# (��
`�����*�̡k���cG�����6���?�	b�� �1F;�/ q,#��%_�F��L���G?|�`3�p�V��CZ�Y�.W��Y% ��l�JTՅ]�d"6 B����Hh�<W�O��o��Ln�M��?�s�W!Rs������x+G�э4ӧ��ߦ|�a8��u�K�ԛi(뉻r:�+]���\��[�c�
j7o4�n�<l̘���x����xr�3iv�������J�����詊R��y�r;���p3���L�P=Ajǖ�g������eW��5�=w�,���SV�)���j��0�Y�m-`��"]�.�՗Y��Z�F�*��$3�/��S�Q�K>"S����Wc[�������������\��Je�Z)����8.��_�Z�_A���ǋ(�c���Y�)H�KW��{�OZM���|��OY�5��8:��bUL5��&��"GR[�是+����L��2��}�XH�Em�Ҵi#��?`j�o��p�u�o׎��儲q�X�D)��R$��.�zǮ�"�^�P/*?^qÂ��X��*��cؘw�/�1Ɍxd��%����f�ͦ�����͉��9(e�����I�R�����I�Q�('d�D� 8��*��?g.�z�P�J�*9hУ�I\z���:�t�Y�zqjB�@A#:�K�;P�K3.>n��Z>~Gյ��3���~�輡\��	
by��0�/��ᚧNF�1�	0����Zk�:��$k�"�2}�����$
/@�1���z
(�T9\'n�r
�kx�.�u�f>$��k���~�U�J:|���c��[?r�O���w[���d_v���%�����ۈ�7y'�������R��%�ظ�������&-{a��nr�Rʱ)���W�k������a��	k���s����������1}��f�$~�]���9?�	O��˼� �s:�CN �fs|�֮֞1g��1۔>8��=�I0�3�xלSTI�(r��qKB�?}{�*����dJŁ��/�SU��<��$�x�<�x��RT���!J��c�N��{�ބ����;4ҡ�d��ё^��7�ؘ�5��?�|?�v���g�u�OxcO����|J�h���"�nn��m  eFcc�?�S����F�� |-3PM��d��d"���nV�Fw�y����!Y��>c�gs�̢��}$��l�.0wz�aD[�8�7=:V�CƉ�� ?�$�h��;蚢s�|�(��=$���"��:�����U�����r����<�?�Dp}�¹�\Ն�A�,Q�F.�ổz��Q�s@3��2���R�s�O�eZZ��>��b��(���fp���Y5K%�[����h�#+R�u��Hذ�u�`��7�A
�}���;�s�Ռ\����"B*<�/l��1he�*�P��.H�`�����$�N���e$-ԋlmֲ״��d*�Ի���R<�r�KG��N�ƻ}+�䳙��c+���E�U"�~:�q|�{)ΘE����I�ԐW���#��.�P�����yO��xKR�$�b_mV�UT��"WڢTj|��w۷ct�G��k�Ƣ�ۡԁTSx�T��e�F.:�ҝ["���O�e���\�V�C/�M��K�*oT��r��O�jQG?W;���J����d�W�)�'���J=`�k��� ,75��x���=�9kf��K�s�kO~�.��NW��@\��F�J�X��B�^9��Ɉ��S>�V�i�l�z)�w� ���H��x��l=�+��L�9iZ����R�	lt�7���|;7uS�������~�c؝�ͮ*�7'վ샸;�����ڕ?,�F	�0���&���Cz\��l_���ש�U�	�N�p=j8N�J8$�DL���T`��sƻ�2�R#ڟ����)� �:m�U��S�6�dIy���D�����?�{ʯ9��lwz��%���@x���߈2|�8.�f�`�z����(�Trł�AI�ZTBN��iF���ڇ���������?���9u���q�1�A٬@�Z&XX��Mm�Fz��e'4���2��H
��#F��J��٠<1�[���*��MZq
�T**����]����:�|e�|7�@s:�\�&ՇfN6�}�H�PNh<��h�(�X�q���H�m�6y�jL/&��a�Z�T�bf��N���'}��sG=�đa/���;u�&�H%ԅᵹ(��a�H;S��0��m���Q9�WIt4�?P������Z% 
�}�ű+w��,��t����K�)�-:7�ߟ��W6�� P�ÝX��
���& ������N����o�!$e牫��̹��&����C�Ӊ9��j=�ꩻ$7�S���*,�����w�g�%��J��ߑ��|Fp�L�?�e�a�����m�.^\�A�2f�uA�21���b�lb�Q����	��P6����_����G�����~'�x&13��<�[�y�Zɭ�;�Κ*\� ��sP��׌TQ'�K��Rx��g`�O�'�j�,1еA5ep��Tcal�s%\�!��%��V�g���%g�T�c"q�#�"�6���i�ZC���CbB��16e�2�Ā-L�<�g������A�"?��_^����k�S=�x�𔴎� �;�ݩ,�B�V&2;L1���&|�\�Rt���g�"F�$��m�*�_�2�{��5v�U&��A�oY��5��n�����1������vkמ����S���(;�ي��W��8(�!Bo�s������טE�h��ڂ��۱�9��-�7!['\�r�Ԧ �$��:�t\���q�X�|����F\�4�ڀhO�lf��`�ۭ2���f�
BA��5�^�<_J���S�����$r�� �ɮ�� "�qa����0H�l�Q�\a�.�c�X�3��ԃ���g@N��U�i�m�o3��E��d���p8WF���[��R0{L|.�0[����>kb���cL��|���e���5��g����L�R-y<w��3�iy@iV�"Xm��0�y$}u��m���%���O� s�UG�`���)���g)/�3|9!����������L�H���\�rS������8d.$`wע�a@��ʺVKԷ��f�ϫ��k+�.��o3�����"y.��!}��w\���$p���
<&��Myzqs@~��b8�ݗ��T�W��?D��5�!'"�!W���m�a�]vG����O�NI~Ы�qp�PuF`'��S��7������R��!B�H�Jn�B�-W1��` tٌ����I}�Ŀ����W;��a�[�|ǲԋ��?� ���Y��b�м��F�ov�pRU�|W��o8[�o��Hk�xt
Y�����ņ`������2�+v�zC�|eF/�q�Ը�i4�;���UK%��O�e����iN��X �V�K}�֤1�?�T���%W��Y���%l&�o�� 
�i�!�׉+t|@xq(��A�Z� �t@���|�<�]�6��t1�����տ��[8*���r��{��65QߍP��W�&�$`1f4"��4S�V���6IG�J,���2���ʱAr�����'�-塓�98_Ѩ�7A01���f�<�k�(�]�l�H�w�]&�Up/g�U�����A�\�p�f�X�C�Ci�}��2O�J.������` �Ԩ��db|ץ��$�˯�X�}!�5�w$>~v�R�1[ڦ��`L�vT8%c���8d)�]C�P�"�b��_�F�E��%��O�d7:���r��l ��^yZ���D��l�ޤ}�����Ս���u��Sê-kh�&�K@x�l�m�-i�n�K$�_��4
W~��e�P����=�+H`�߂�麱<��Y^�p+��Q��>��~�)���h�Se���AF��l�y^����[j�fF���Ϯ7��Օ�,��h��6	��p�
@�>�N4��<�D������<�K|a��2'�Ik8Ӱ}OI�t���_vk���.^'��(\�W�o�`*�~���o͊�N"��F�^���pc [���k�{�bDG��H@L����]��ص�����T4��9.�Ӧ&�v]�*����7��"�Z��D(��&�NR	�I��>lQ��;�>�>��ͩiK�0������4Cz6�G̏��������J�*Eu���V�a?���h)������U��eC��?�� !h��ue�1A��,�nI9�N�����8~���̛k�j��a�nP�d�y�{_���dB��L���h��	����f��0-���`ҬS���i�f}P�vC�]�GJ���a�: �$O�0�.٘�1�"_�}�`�d��s�:�t��8��!o;�x�:�~�E�F���*�<��̲"��!U�ߣ)�Eo2?:�Q��_�ҸX�����,�������a�~K��?�6kX|�5�?�H-����2��~4�7�7���^p^�~�e
������K���f�"=6K+i�݊#��D)0Ym��U�5�L��
W:n��>o'�--~�,j]�@�R�w�2�<jSĎ���B)�;`��n��/��a�Q�/�_-��T�4�+��ǁ���/��jO�r+�> ���
�"ʙ�L߈���W[4W���Ͳ��P���%���'�wD�E�Ot�\�^���s�',b:�>m��D�폯���VB�8�|*�~޵w,�W�q�I�4&�a�Ic�H3-xQ�f�8�(`��Eh��Y��.����k{7@ma���^M���7�}�hm�,7�������:�9����y���/��Zr@����go��ٸBLPa�@�� x3�H�|�T�ɭo����YB���	
!?���T2��b`.��޳�ˉۈ��#����/����Ȍ��SN�D%�"��,b{e��8|��Q��`מ�|սІ�c?�v��� k؏�AۼM�����o��T�!��]���=�,�E�wl'�Ny��y'b,����_E���=�W8':,����)��m����D���پc���)w۽�}�Q2q��s�!k(c�lbu�����t4�=��������9��}�qag��K������ҋ�*���!�ԭLMK~ Gd�����n�X)'��w�H]�͜O�1f>�Wt�)f�x� ���������;Ţi��wqzN��`�&�B�m&����<Mfo��U|�o����`)��v>Z �S҈�\�h�nRׇB�+ˈg���㬒u�4���b=�ɐ�p^t7in� ��OȎ� ���V��H�J�I��W��pZy@-�w����(6j�|����9\Ǽ ��#�$�i^���%����	�F�a�����#�>���ƽ����z�C�G��[?�=�E{DJ�wfF]����VP��֌Bj���&��]�ۣ⾿��(��
qO��]Q�M0��/�'d��$U?L{��`İ�ȑ;Yޜ��$ֹ;P����1�VU��X��k�RBi�v��O� ���
��q�áua�^� M�\Τ�~�	�7Eq��Jn*.( �B�q��B��b[����j��_��Up��{L�4�M�ލ�}ΗM��Z��-�{<�I6B[7x��!�b!�%�2����{�})�w˅G�|ӧ��ܓ�+�@�I�L^�y��ވ�c�G�~��x[h%lf�}� �v?��)���L�+:Xm��8�Ƒ��"�ğ���(/�zh/�UG�qE,Tr�"W�]h�-�t�B���,xw�{��R�b*������xlCyqGZ������B�I��߯�Z���Dhx��#����˼����K}���E���v/�m�)35m+�Άӄ#+c^#�3'<!�H�c��_�97N�y*���H_���vBzk��
UP,�+H����S��{B:0�VV������z�i&,wBF��"�>o��X��b��S��H&���#���z����'�-�"�B^x���0��v�+��
�k��Mc�;�\�>u����c(���,m��\���O��aj�JM���l!���E9�}��:@ڲ�T%T���N�=�=c�X�G;f��V"�.Y��v(�F}J�\t6��b5P�&��.�t���(rcǨ��{��!\� ���>��OD��BD�h�	���f��.�=y�|�����D"QXJ�4��݊�T�
��fII釿]Dz�!��� ̮lp�*��U����?��x�˒���!��S���Lb7�	^)H��R5��"9>ϓ&�ى�cȢzr�6X�n2EΝ�Ԍ��D�X���9V̧b�!P�!���18�a�pd��v-�펅�W�ﳌ������/��G�������z�$U��1+��ev'���k��e�zxjv��"m?�H�Ô*�+���'�*.�usݽ�Qw�b��R9���'M�M$?���n"V�	�DLV��4���(���!�>T����3-9X�eI�(�UC�1��✛W�a �ʛ��f�'��L}j:-ٍs��׸�N-J�t#��T���*��:���	/���8�(\Q�8-ԃ#y��tP�>����m�^������i�����蹀��h��/��h7�,y��H����b��MG<TP��4��l�y�j������G
��W���sa1s��r��S]S��!q�έq,��*W8��,��[�&�Z�!�}�z���#��"�o6�%���&.�b�hl�z�셋2�H�V2'����ܖ�Z,W����P��j�����ά�s��R��f}U@�%�^��̱��»��<F� uhP�������O�����[-Pg=S�fԜ�e�	�Yii���N�����DD����<�vA9��Rl��K�������]-���������@9���q���{��<�����AP�!Idt$��n�V���$o�^�G��@N���C�\(pD��/ޢ�[�C�3g;z��=k{�sq��ޅ�CPw�+Z 3<&K�B!$?�6w�����M׺�)��6���
cB�CI�[���A�Gή4$��-m�7�f�E��-��S� ~8���O��_����:ܿӪ��v�f��'�	(�� <�u�$�\ '<L��TOd�V􅜶8Ygf�2_�?����|Bl�ΰ�<dӏI� !՚rB��,��7̯�# �����}y7��U�����F{���y�F�8�F�W�`�|���9���^�<y<����R�u>��J����@l�Rܽ&�Zu�� ��W̲ |1L���R�^\�ZE51��9�)����P�HN5��g=����*���%��o={[���]ܿ�}���쑻���l�*Z�Tϩ��� (�)����-� m�́�o:�^�nG-TY��ocǬ�|Ѩ�U����M��3��~�Bx�{볃���|�T� 6N��O7�K3���]q=��SdC� 	��*�cN)��I�*�K1�?j9�說;#�Ld�T�~����!B�� 	�^��Y_Wc�>�2)=���e�~� nG(q8Z
�P�Ѥ�D��<3<��4˼@�u$e�~S�~�Osw��R��c� ��W��勬1:��|xo�%�z��mN���9+�TfO�������~��Xx0޴���7���#0�y,lb�C���`�i�l���"�M�\���n�vp\Y��τZB��[s��ڒR����#>|b�î�5ZД$��&X�<n~��zx�F�0Ƞ�L�l�Sꌊr���i����'�u�
!E�3������n:LB��|�e�kU��5}RyuXv2L�V�ߕѳas���Ǫ%����NK�=���:��vp��ݿ�/?P�I�ɨ4�R�6�]��h�|*��YK���\���2�����.�\5�\��k�r;2
�uN3N][�ӷ�'�ء�a㴀���%x}H�2���	y�q�i�2d�$M�Y)���D�Ϧ!/�ʶ�,Ҷ�t6�o��,7��>�?&,i��[��F��E��?��K���F����mמ	P���ޓD�'�$�
��_�� V��Hȣ���D<�\�������AS�����;\k6
+jBJ�r��Ũ��-a�?���l�@ �����y�\~z�p!r��BByi�ܾ)�����i�y�<�/kF������N�J��х�b
��*�%i՗�.j[ҫ� (̜����U���Ԩ{a4�$�3
~:^�_.+*t�]h��@IΙ���?(@O$�BH` �Քq�QC����Ͱ�9��K�u���Sl3�/	��槬)���ãy�Rˈ���lӰ����Iz��E���\��$t�89u'u������Д��zz��x�7W qx��~���k��%�ڼ��}�р	��`�2�xPC !J��Z����g��Y,^�߸��)�G�DS�t�8��갵@�l*�]��65��ӓ�fb(ɿ���'���Y�E������3��Z2��{aZ�6��W�
����@�X�-0�;�+�h�+tgE`e1���z8y�Mt��cEv�&e��d�5��~?d5�Z=�`��C�8��pR돁���ч��WH��}?�c�K��1�/�£�x�����.��
�!�Г+�.LÅڀ���l��<�/� -(�ߤ�=m]��2������:˶�����L@7b�;��O3�t�L����V��ȏ%�ƚ�S����az�'�9��a���<3�0Y��ԟ4���<M@=���㯉�"�/m�.CJ�7�s�`a��PJ�W�O?W ����d�~APZr��TE�Xt=�R�-������s���������o�h���M���qɫ?��HR�,q�PH@CP�7@~����͘�gO�iuj��&>��dO�	��NE��	����r�� �;�	�����p����vq�9��.�ȽP�^"Z�0�%��ue���?Ms��u�FDC�|��'/�օ!*����dR&z�C�a^�H-h�h��b�����x;N׃L&K�*>� �G�FЅT�������ѳ�W`�ų�,?�洽�'��>���:��y�ry�{J��#M��Z����[�����b�j�1y&�8���/M��ɚ������*����/!�'W�˫����	|���G�	�j���ɐ�#�`��̀O3�S�No,�Z�1a^�m�{@GW�sUbR��G����-��䀮���>xpO2��m�Yz�I��*������G�{���Rý�Xn�� a�6K�&�}(�)�U4���W"i��'M�+T���\���7�掄�%�3}UkK�r�}T ��4A\#q����/ʡ�"xT5�؛kS�#1t�#Q#��� +	6��kdObא+vJX��N�җ�%B̮J�ν�"S�``%��F��!�^����*��
�%�akn+�d��P�5�@�~����"�$�q�'�N7��1�5҅��=e��-�G���}�փ��Q�ux�����0��Z��+�Q�ZS��|�w@#"s\=�Du;�k;�κ�C`
�kA��$D��;x#��u'汊D�8G-��K6t�zhyD���jH������x���+�xn���y�����QZ
��Y�IӣNF�F�(R4���RM�J�/�Yu���gTo��LY{��l�D4eT�~�U!��|�T;���*&Q5.J�'{Ա6��Gފ�?oUX���07no_���$�!9Fvĕ8�e?��Z����ǬO�dV�֙L��*�5j��]�L2���-:����F���z��V��W k�Ց5F����e�o�!�̖�}�� ;��|Յ�j�4������2'���i����D�B��:�\`�2;��O�?�X�me�lc��|ŹQs$�{�J��_P�.�I��?���I�<%`*Pu�*�;���O��r��<�)#_����ռ-���&B"eX/�(m)gt�����Ǜ�D� r>�<�[d �wtU.XE�J�إϦ4o6铼�S8]���a��p\��"��Q{(i�;	g����fl�����o�,;�����-㴲�X��p�s����y��T�Y�%�3�mh���P����,{��a�����b�";r,���S*d�q)�v�2�Q��l�p>���(��)8��*q��#br�	���ѳAvM 6Å�TsC�s�&��;5��jD8�?�@�`�Ir~ڢ��(	�A-��� ��蹇i&�V&6��A������4�iZ�P�*mk�ף2�k+Ó*ӟ'�ԯ���@��Cj�]���Q��S(H�΄İ�O2+���c<z<��e�_�#a�WDo}4rÛ( �2���L���A�Mm
���tr/(4uPa��c�$������3�3��4%��Cf�Yej�=Z@b���Z±��'k��Iē����_Lwo�E#���/�?N^��ijΪ��/[_+�=:�Ƶ�^�Hz�4��ȶrb���njWpFwY�U{����VyLS si�����f$n(ν	��,I��"�U`�H�ϵ�E��4�+RJ�4�����ʨ�i�]{��L�G��C؍A!0������UZT�b(�]�>��=��h�,g��M�(�s&�M3����M�[;��tYՑ[%]��Y薲�!4y�Pɼ���_^w�H�߮}�W~�ǸN$;�U��`l��>b�:��Z�'�`-f����n�'a�h���y��/�y�d>�֯!kD���)I�^�j!�p	��aw`�q�<�GS�ǺTށ��h�aj��D�/.7{k� 
9��Z�-9�H�4l���P���s����W�s�o�]V�&�H�X&�л�i�,���Aq4y�����n#���1��&�u�ඩ�k �T*��%[�I�v;��)�����i�j �9[�
�K:x�F��ӾVp�	�\�B�İ}gӠ�p���(�.�mu��I�*��,� �0���N'l�0Q���.z�V�,�� l=˺��؝��|8|���r�$A�����a��M]��;%�o�.?G�(N�n�!K�To��4ߙ���JHxnv>]u����&|T-+�v�#���^5vG�讕��B�RL�+7C�P<���HE54��2�`�P��jMQ�W����2�p3h��]�mª�!�rn�Y���W���3u����mv��K�h �']�Ű��`�P�h�Gۯ8��R.�L�_d�kv���e�&N���I��vM,>�9�0�A���ܱ)��C�'���c*t:��cN�$��',q� ֌���P��H,�K_��v�#~��P��9 AOm7��s�Ʌ�9Nm��ƒ�J�:�Ez�� :dq�ə���E �Z�g��M7�K���?� �W�-��B�t,���,�_��(-����4�w�f���4�c$�����b�e��G������I��F*�L��u��i(�^5�T���U��/��pO�O�V���%=I����������'᧒e��Wx�H��|��gH��M�jp^Z� ZRӊ�s��`�vK�X8��8N�^�`�YI_�N��l�;��o�e���䳜G !lut78��sv���ެ_k�-޼=�}�p`b��b�0ױ�Sl�ۡ�W���[���SD[u>���ʼj�׎���`$߇,��"��8)v���V]nnB�Pl�J*\i�H��(�3~�B���?�~�H&�F$�|J���T�W<��r�������t��q�}�S�&u$�)�c�g�^o�X_N��s�MWȰD���B$�!���ʇ�{Ux�X�h-��(;���%O�5dkt�_V�X$h���X�Km�=�~�,E��!�+�Z��x��<�U
B4�-�/6_h@-d%iWs� +����u�9��'��!|l��;2��u}��tc�F����~ތ���~*R���ۡ�+j��u�f��vZ�cj�ItP0?���p<b�H�EA�4�������X7�����D�5Fy�F&�Yhۅ���Y��	��2D~c+҆�p�06=ǃau�Z]�튝�������#�(��̶���R��ȾsUG�FIo�Xc~�L���>.��:<�t���;��Lm�r�L�oPЍ�)���3��s�X�{�no��:��ؔ�w��#~�T�������j��c�-㽴�g����a�F ��o�ɣ뿯V{�f�%F7�}�ܲ$�R���1��p� ��$�c�2���g��f�zH���+ݬ��nc>nhˮd����S�r�U��ʝ���_Ew5ơ��D�E���/�.�f �!�ڎ[P��}�Y<ҡv��p�b43Au`��iSZ�l6��?���}��?��NPކx�J�ǔ<��Ւo�&�Z5h#YG�f�
~�ҕ������_%+�˘���� ���3.ѩ��q Ȗ��n�ݾ� �x�����Vj̢���!K����?�m���ս�Np���y��h�.� J�ɤ>���5�Ê��z�
=��������V~0i~�U?��wD �M۴����u;ڕ�����Ŏ,{|Әx���R�A�B�������t� g(�\�/
����0�����t{Th�/�&3u�Em��y�z���a��g����������ieen�jL)Y���x��]3$Q���~�ej�NEv�ֈ��V�,ANx��X��������$xz�o%�7�*�x:�^iq�ঞ�C躘&�u��P�H��H�|�D�AC;Y^)k+:<�H>jt���"��%`WW����X�/�����P@���p�S��bX���@*�W���r׶1�4��.��^��Gͅ�/_r���u�+\�c��
qn���`1:����a�^	{臚H��M2�o�@��Q@�-:����kd��0��)k)ʍA��#��O>�_�����E���z�� U������F�&m�����0]��)$Xku5|�RY�*�̅�%ZO�������p�����i��L�P�A�����nJ�ӭ7�?�\�=��Y�����J0�n�Y����MA`'�{� �B �|$ͿGc��F0�?e.2�RI�i@���Q6Ё ��Lk&2�-4q w˫s�l��x&U�H�.&�:�-�8OmW�/Ƹ�7	W�^a�����k��7nK ��6��T<�7%�"�ip@����W��Ѳd*���i~(lhy����wQ&�-Z[��pi�8�o�G��I���?���B+�{TRAb	�ZV�����V��b�]��U�ܣS���*�=�nN/�/�y0���V���ϓ�+��i��Y����A �<�p������ 4޲��B>�B4G�#�k~�ǙP�fG�F�1�~H�t�:�ƾSch;��� �z�,�Z�)�pA�ܗ�������+�˩�'ۚK[.�j֞�Z�
�d�~�6t�gڧ3ϛ ]��^���yHb��LG0�׬�s/�ߏv�E8��處?m����hje��J#�nɭ��/5����w��a޻bKʌ3}M,����<��(�?&��Cv�Hs�ю`
+��]٫��3e�N��2�"���e��(�Q�S���.n��%�%X�w�8�B�w��(�I"�=���𥧩�_}de�>��s��d���Y�x����y��0�ڱsH�����+�b�(���{��)	M����(޼*���~m�[�`�d4.�;f��5��c��MM�4_-�\���)fJ�!����Cu�,�-x����-��ʊ�E���Z�?��V�����8 �ᰛ�`B;x��FJ�0�tGꀹ������E����31���0��ni[^&�Q�ؕg|a&�\����6b��ķ&a�w�	|A��ps^�M/|�I��p�9k-J�L��B#����a�s�~A����!�oI߾��*�ZoE�=�*Ah�ԙ�@j9�ʾГ+���3�$�R萗�~��L~��K2u���P>����{����v�n#��O���h%1�N�a����20�Ԅlg�b��ߖ�q����]
�`���b")���u���䇴-�3>�}>�4�$��X���3����ɼ&Y�!q���s���b�#~4�a#���C�YTtP(1l)/��{N$7wgF�������fL��O�=�$�)�D�=�� _����5����#�,�Y��0y�̟�S�l�A(�	#4��W�΋\����g����B<�ہ�X9�U3W�S-Nca_�;'����d=�bh��$����8�U�6�u�@�*�P��L�Dy1=-��K�Z��:,���mL���'Xyڱ6JvC���a�i2h'!���2#r�0��b؀�6I�D�މ��������bM�A�2!��D�ʂ}˔P���)�a;�A���۪�#�ޙ��֓�t��賆������ ��9����&�t ��܆F-���fE��>G�|����v�ll����=���d�3��ǻ���}�R�"�m���h&��L��h����y��Q�/�k�b�#�ϋrH��N��@V*�w�v���>�(�[�~�HDΡ��{X�f'�{y�Xל��~(���u� �:`?�8)8��,�.{�����K��|l�Q���[l\�|��QiW�Y\��S�v����J�E�w�١�T�g�(Ե�4R�F�V�bw���p,U/$����σ�N�&���:��n�s|�S��յ/��p��S�j�JH:��TK���L��j�I��q��2c�3ᖴ9�Z����8�F���y&| 
�gT�<�Tb�b�ʫđ@#lw4k"<�8Ou�)bZ��V͒��۾�>J���.~T�Λ7��Q[H���ԅ�D�TK�H
�m��O&s�7 k�<�k��8�M`�*���J�W�k��z����~���u$�@�nD-�-�/��M�N�j'/E6K@�����}�9��(X(�����;]��g��Z���IH{	��]D�Һ�G
Ԭ���+�"7��c�lj~�� ��� �g�����k5,��;ji��sx��	������*`��H�Zi�u���軀1�Xp���9)5Yh�b4e͐�1[^Д�y����Q�3���@>bR>�=�-�_%X�Spe�*>$�~�׶����n�GxW/c]�x�7������U����Gb�s��v�ږm���ꏩL��ͱ%�1����d��9�i�S�f�N�b��d���hb̠��b�s��h�J}��M@D�����g6'�~#Zw��lח���Bu��(�8��~����<7g�@fR��S�L�/1�\�[��+2�|��&)57^.
�$��y�Ec���$G�ηz�rY.kx	�\����>��FI�T��䗩H(S�H)F�1��y��G�LH��P6@j�-8X;�^<�i(��]���_��z�ȣ=���kR�7ws6�Z?���L3��;��[!��p���7?���2��`ê�YL���NO�S��H2G#��{�Y�"xAW -�i��ޚ��Q����Y��'1�Õ3�FRY�w`H���Q�"^E���&7�~{�&�;�8^��y�@N�}�r4HMnq���Szn˩;[��}zI0�C[}�+��Y���\̩ �U8*�r�1��RD�Bd}Ş?�ӎ������n��U�;����.<�YS�L���Z9K��x[��x�ga�%i)���4�A�&X�t"�i=�u���h���I�߄�fE��n�h`���5�%���R���>J^�*�f/&;n�@��"L�J@�D���Ur����Cdv�P�S���L�P�x\y@�ɼ�-�(,u��Æ$�{��
��y k��M�c(��_e`x#�|���Om~>�|T�#�z�`���>�d΅�"L���u>N,����\;xe%��D��=�qJ���!�jVz �� h;�D����v�̳͡>W�s���8r����"������hߍ,�ޔTB�ԅ�C���[�7���>��2>�*b˘�=�����P��`�ʽT�(�h�|WMG��P�d|:S��k_nI�s�Eo�cj��������p� �۳���#�5~���*�O�Mn��|Z�Q�OZae��:�l��a#��x�!�	�� ��7y
��s$�m����5��g�.�Z�!蠤h�+o*>�U��P�{}�f����{*\���
�����)\Nep'�d���A�*��-��b��5X�FHc�A�ٕ��N>q�"
e�B���������X��zt���C���J�Z�u��|.��ȡ�2�xh-^��ʃ�i��;�̧WQ��C9���a�����e�����z�l8k�E�a!�-��D�����1`mu�	m�������n�Ā	�%U9=яLx��`�K~ۦ��w�GG���|��hT���i�v�h�|0˿3�Y)�ŷ+ppGY�r���)�s]��8��-h�1�d&+��>TLAHŞgۤ�g�ҏ^7�1����F����_�=?�L�@����7�6�4B?��_	��|�B���s��dzV�.�u��"��񳤥q��ѹmߕ������CV*ȸ�;�B�e��;(눂BOF�T�����\K�*�owI)(�\�����3�?�{{u�N���(�*�P6ܺ�D��� �m�e͌��b;:�J��b�2�������N�{�WN���d4��-O���vb�հQu!:g��Ԁ�Jd��mE!1�GG�{s�o�2z�{j�H����.r��҅�d�� ��q�l����i�v�󳢝:�5��N�ë?�V�T�|]�G(��lob"@�"U�<�;�g5��&)B"-��mC����Ͻ�:wmqG��q`�Z��e�v�23�k{���Xb^'�%��;�M=*M�s��`Hh���aڪoBz����s��U�Ls��ik{�m6�*
>ƀ%�U�|�B J#��� �#�#�@AMLxܜ�ľ�X� �1T]]��9\��|����� ���`�Q�Yc��4IiR�K���I��\�a��p�:��箳�\'cѐ"؛�Ʒ��F>�̄��h[Z#\R>���遁���k�|�Ņ2�i��<ө���u7�����x���4���c���1��~Ϛ������o����`�^�}a����\E:�.�	Vr���������B��`n����'��jb��HBm��v�t[�O�f�YX��I_�����N;�m�����$�B�7��@��T�Y�E��P�c�AZ�}����&�X~���Hn��I��D,�{t�^��i� �"�+b (۳��aA��n-9m�����\���&:\e��~�
�4�H$�S�p��e��޲pe�]gS���
x8O�� (t�G۵^2�D���%l�U�ά!��V�跩��q��,6�[U�c�1���%i�@�K#��#�fRT멥�R���������!�Ы�)��];?�;q����<�ro�)K]D�kK�����*���hqwy\޸�jl��]�����k_]3��@Q�� e;2�֭������e��,%&&�1�.�����'���}�r���	�2��[��}lָ}%�8���t�W�p^鰷�zH��/�v�}�0G�	c�v�4���4�7�N��Մ��D���J2�G>��A�=���; ����ML�,:E�#}�8�c���~�����p?�~u���B9�У��d�U�.��Ygw&#[V������-7Tͥ.@����[�m���ۚʀ�5�fU��_΁�i��k�\�|N������_'�t2uVs��c���;XF|3"+fl����.w�We�r�a�T�"�Q�N��rd����b*������e�lo֌�Ux�/�!���f�	i��~��	�꦳������1���^�{�.�Fw�IG3�#��hW���c�to�-|��>��Ĳ�%�����Qr9O�g�������}߰nI�=���&��O��Ԭ����\`�8��Gs ��`;�BHEb���0�f�jtB���y[x��"�|��;R��m��������sJ���3|���I=�p�Gu�Y����}�x���4�GȈ,�	9���3�i�2�����)G�,-��8ٵ_s�:Vq�ӫ�o����cN����aO�Gc$@g�s���А��@���Tڄ'��4��&M/��Y����T^���(��+&��DwY���/��,���8<YK����R��=z��/����!����V��0D�Lit�R���5nE_]�4�KjW&��۷h����@�����?U��3�T&0�,q�Sb��P-X���P m��ڰ�u�����u�~��N=M��)���OU�"�5a��{.4T9�կ?�H=�HT)+e��@Ew�R�|4����p�}�w��T�m)��[��/�R�/_܈(:�= �i{ǌ��0*a�1Z���*ь}���p��r�~P�!�r&��r�ɍWτ민� nц��ƫYLw�k���1D��ܮ!�)d>��Z��Gꂠ˵�i����)�Y�� ����X԰R�u!	��=�����\v	К���복����֣�	��Z��Pw��b)��5���:ʤ0�V�I�'˗����5y���lЋf^�S9�>����%e�������â��Ȝ�D��09������6dj��fuj$ɸ���ԛV�H3�Ƚ��$0�C�m�T}�C�;�V�����m�j��i:VxS�u>�XC���Lx��}�m�4Y��&����y)���������~�!l	]�i�e~�א%���V���غ��s�`q�AZ�$
 )�����,�Twį�=�ސ]Ēg}�ѳ��W��0sz�bxx~:xr�Ӓ�����dű�d�E�[�[��I�uX$��\>g������T��J��/�ä��{�f�}�VyR��l�k�Ţ�tS69���'���y�	C
�d���S������f�RS�S3�a�%wZ�@<�}D�|��&�J!$3{U+�¹\��H������b]ǌ���j�V"N��b���L��������8fKu�+��~�pA�y�Bj{���o>�<�?)E�)��/���+N��c#0�!�M�n	�?D�~�(�x��GX#V��6|?:b�����*a.�Ə��F��w�R���2�Q;*M�mx�Ň5�P-�S�Q�c��F�M�%�?HVE�;jԄ���Pٚ�3kH��^�����ȉ�y�A�~
�03��ɛ�f�c�%���=v�%Kh��8��B():�i�(f��oWʼu#ˬ����I2#�Hx+�,c���+�dXю����c�F���r1��j��5���*�,a���vQn9e����Q~�$������T����@�(���$x�E�<0[���b]pgD���2ь��\=9mP}� ���Fi�����7�`ǹ���AR�`�� Y�.���%�y��,X�hP�@��ٶ>od}J�I`��r�;W?a��W%V���s��[����Xɾ�ĵ���e�<�Q��H9<��fǀ�S89z��t�[�v�����pX]�p|֒�s�ᙱ����eO�������|}t�'92�����;�J�F7�߅��r��n���`�Y*�JtŊ�ؐ��i�g�hu&#7_�����;��u\"��:���s�Xbd�����{��fu����ü,5�I�쫨SvV�yх��cbE���3�
�'�^1宀�_�ͩ]&����#��1t2�A8�f4\п�E��y@n��ב:��s��������I[ɽ�E�pj]�=�l�4���iwSzp�Ԁ��_�ugЩ@�œ�K���ú��r(_�x������e/G�呀��?-0��!��ؖ�	 �� ��������`���a�sx���3�2Q���L�_�$*YI�%~)?4A�8�E{�B�RZF˒��k$�"6?MۤzG0^�ފ�9��]��*\�	dK3�$.�Ȫ_@�.(�-8�Ҷ(+P�B��4����Clk�Gإ� 򎗻�~�ʦ��E�&�a�4�ȱ��D�M+�Ia򓖗�3���gr
��"����`{`�tT�^攭�6��JK0�Λ��d��*�rP���l�I��ķhr�3��F�!*�GH$J�wG�D�Bt �{��	�Gl�	�����?��p$Ӄqy�в�"���UF���@Fzv B����'�/�3�&Q���]�X�Qt���pJ�@d�����P@�ܦHrL߆r�e=�і�{�Da���������V�õa��PF�kB8�Q����opP`��@���E79�	T7���>[P�&�>�d4N\[�t�OQ��??}։6�,���'޳�w�b�&��N�;tPp��I#�*1��G�cWg��9*(��tL����0v�/ @�?����x���M`�X��m��c�5��홌y�u&��y	��e���c0�X��}I%q�'vg�Ls�#hfxn}�D��*H�$�ֲy��  ڂW�7�2`,���$ժ)�[���j���m!mhe�}�Ľ�V^��R#?��.W�s�< ���qgJr���ղ�EX��`E�U$h�꽿Rx��?)U�bD���˝��q��2\<�Ц'~Z#�Q�=����lP��>8�j�g`F��T����K"��"1|m��H��{�+pCˑ�Sz��
v.�ͭ ��%O>��s�E���%���z ����J�y��|��l���T�C�ji��ML�5��_�v��,P�!�V7%R+Di	��|��eѡ���N�_fcL��%��Xy���l��	щ�6�����#��a*('�%"��qA�l�����%�X��gsX;��N����M��=�&�=��/�c���ە�}��,���-Û������oZl�H���)��b��zNm��B��6f��Ҵ��6iܙ}� �R����l0VI%���~�����a-�����o��w����P	��~+sbǋ��������g:x?0Y��*�&��I����i���V�-�n[�K�8�y�]���Yk�"E���J�3�h�X�$�ԩ<S@�Wq���h�k�jAT7��*fg=9��п�D�H6��i�P�^��&^�1*�(�~��� ���
O���a�k+mY��,�
j�=4h
p��_0�-G�2:�"�Xi}g�#�&��$vi�8�C��s���� cGw���3�G/�{G\�FjW:N�ʓ�̝��YN��ct[�J�*ƤJ����y������-�+�YFF+w�b-t��vc]	Vš�v�o�+g{NʯK�%�Hfn���1�C��:���*�,tq-�Iڿ=ؤ���?J��Uz���nfq�=JިB�e� O�C��@oB�g��Q����F���=�ݲ��9t\�0c�n�N��)���DC{��lgO����&����5��U�Kb���9�����^����
�v�|�j���X�ֵ�{�x5-�Z���&Z>�@Ej������D<�%�I�[2M�	�7��Ǐ0��J��#0@���r�S��1�񊄀o>��ck�R ��o����A�����a��՘+~^�V�~yݾ�1���x��1�����2ڊ��
B���(��#��HvA}= hjN��PT,�	|Z��,i���o��� ����d>Us��!���()�_fS �U|X�h���F�W�upѠ� �׳�{Þ�O��f��)�[k8v5*�
�m\#1՟�3}�����U�m?&�!i4(w���n��L��U����2���J����mX��ܠ���e�"Z�
JS۫7~p$N�:���s�ςP=]�v7Czc�6u�8���$\w��w���������4b�*y{H$	�9t?�-��.�uZ�4�^w)��>�����<�فW)H�žnJ�Ā<�C�YC+�OL��D��	�I�0��YC�iW�:���J��rI���O$D�u�U��lցyr�{1e7j��U�gJ	�ۥ��	�?J�x.;Mq~c�vnt�"NQ[Y@��<�Wc�hR�W�ڶS-"ݠڎ�Ҟr�X���}�=~r|+�x����I��k�KP��������������x��Gw���M_V�,�qԌ��[ v���G�hT��8i�-F��o�Ȭa�m�pF �
�iX|HU���k�����<�S]{;J��g�t��'@,�Y���kT�OP�u�C������w1�����/�DW��K;�`�*�����JZ�dxL�n�Ԕ���ڝ�X߽��e7>'h��) G����=Kg%.�d�� ա"-ԭO�N8����`�k�E6+�~�EB�p�GqT~槛)�	��\AM�uQ`-[���{��m��YXkM�A�zްD��T�..g ���~]F
��P��KM�gV�x�����%Y��r��y�'���t��Ш�Y�#�3�n��U�������D&�����^\+���=�}�C���g��$�R�q��7Y��T����O��׷FiP� ],�$N�Н��T����rQF�S�x�i�A6���J�ɞJ_�%�'Y�h��[!6����Rc��V�e��H^)N�)%S��F�@8�r�펀8Ϣ�q/mRTo�`��un��L�vm�����W�D�B��%w���q�1$@�<2!*`&�-_=��R����a��tV�a�⮋ɇ�󚠨���j���M,�y?bE�$^yn�%j�p�Nv���iYOio&�nL��@{��d@��U��K��8WIX��ɭ��x�e�	����;��8G���{k_V[���0�(��b<y�O���A�W��`P�;RڻU׷�E��h����F�$��}O÷t�����L˙ ��9�����~t��^�����)<Rp`l�٧��k�����"���h��/_�T R����v|�����2[�A ���V��؟M{e'�̺�kO��y�o�)w�[n~���l�K+������N� i\�	�	��SxN�f���4�4$,�=3�,MWl	!��y-�E�\����ެ+Hd�۸�=_��WR�HǮ�k��YD�v_��Ǩ�a��&���J��S����X�tf�m��*tI��;�|��PY�:�T�pN���Gyuv�!Mlύ�ְ���r�\4���i%�X�8��,��F� o��\�ډPq����JSWF��S�_h�Z}^��X�r��;��¶��U�����!rUan[u� +�����d�������IЮ��/u ;����xΜ��E��)���5����CI�]�֊�dJ�q�Z/ns��{���Nru,�,}�Z�<O�һ�hi�˹�+W�iQb�վ����]�sZ��G\�=���\��26w͉1۝��>��x�$8$1~���M"W_{>+���Sנc�,/����H���i1�d��%"�IG/O3��dA���(��Jɘ4��׌�ߙt�G�'��Q�q9�R��-c��>��S|�	�ĒS\�������87����0���ނ�;;��3V�	�Z��?im��.���i<|��&�v���	��*8��+S���,������~Q�S#�P`�V������'��td��%�l4u-�i���u�u�J�v���!(H&�����z�8��J��
�	BO%d��������ܭ�U��O�<��A9E�
&Ȍ
h��V.!Ma9�߉��Cjf��~�5��h0h��W��c9xgBR���/o�u�U�D��^7���ޅ�639��< H>��Tȹ{�Ʀ`�_����>�ۥx�M"�+�p�ʩ���T����D��r���s��I��Lv��zz��*�2�J�U$n��<�ש��9,	��`Z���k;�X�?��Gd��-]�a����&�	}j�F�4���~T�V����U�ߡҥ�	�4�s}G��8j~��a�)<)UH��O%������&�QOUs�n�9o.��6΀2i����a���ƀ$�`����oPY�J�wI�=	�4&�{Ԍ�_E������0��_J��A���:l�n�#��ء�"��0��(Ĩ�B*Ԇ[��h�ԛ��	JP�k� �Ȓ�|��-�&;�����C_e��l���~��O`f��X}�,��+�����=~4aQ�4,ȳ��2S��>ܙd*�ׁv�~���K	�p���c��8)�q��s:��].�$lY��/F�Jm���G7p��NU;�z4��jg�����K�z��N�`W�)Ȑ�0�C��?}�SID�38}}O㿕��ꭎ�(hzA��\�LG}�f�2ΐ��~��%�������c�3���Yo��D��H�@0pg.n��©�o�=�����TweI2;z��L�Mi�,~��h�? 竵���/��U�>���X��}���`$4e�{)[ �Hz�����d��qV'�J�d��]�Ǝ�b������(���EY=KO�#b^�7�U, ��Ψj�*���Lo� 
6#u" +�6��H[RL0�|�&��r*1���W�� �����ڻɂ7,9���kW�-��!M�!௕7�ۥ'T�[zpl
\�2�1�,�zyl���:����8�A���F�Y�ӿ6�3�]�ej������$��6������K����z�>��AaP�]�vu�!�V�8G�W��G�m&�u����qc��/���^4��`���b�A��s�:pge#(7Tf�ŕYv��������������N�6�kh�]���I�,x	6�u�lf�!�#����?^�=Pe�R2/<��Yh:�NÈ��"��49�����F�S��9�.8K�s� Ǚ�%)������� q���/�_Ȋ��o��΅ig��i٥f��I\-�ڸw��ow;�լ0;FQ�� b�H��c,�n�3���r ��'ŧ* 1v��'�e�����6K�(k������O��AX;�!����خ��&�����ѶM�E��s3U�Yi�8��G����[���iCz�Q�,�����h8p��+̴_��z� t��*-�l���t6��Gi�l����(G_��T�G[p�M�mS���3[wխ�����wY�:�l����ꕾk��)@�ζ�]~���	��Y��͘����
�C����ʇ���p��׀�}�\T.��N�sr�;�9"W�8Q;��P2V
�����p�QeJsB�̺S���U��"Pğ��#-+Op�d+�J4C�T����ݘ������x"Gw���V� T�5c�t�s��j��P{����}��
Y]_
GX���ܶ�)1{��n��U�55)�zq��%��3�nM�盒1��9d׹�&� WP�F��_����?�D��.�M�(�~�g�����zI�b�a.�����.��Ø���C����l���N2(��*�Y��y�ľw�H2F�;�w����J������)��'�t��������f������3�r��x���09l~((>K*��ɐҤ�
QY������i��ڟK^�ƿ��^�|�� �'&�_�z(��SF^�����J�Q�m�ӂpPt�h0i|�G^�~���s��":�]��v���|�L�!��]LU��r�=ˎY˪��µF�a>�t"E��ƔR�ǌ��y��O��L��4x		+��%�	)���<�K2��?����B����ϫ��\����L��O�!	{{������K���T��<������%�����U`�ٿ)E�>)n��kG]l"�]W� ��%̣׵�7��\0�l���6����JSD�Z���!}�ػĸ1�Ux���<��N�� ��g�熋���3R��8Jmm�⻾l~� �qY`J��k0��AH|3a(�`WB4Q����9ÿ_L�ʙp޿����+���[�/\ŧ�3p
Q�t�q7[}i+�gT/�\�h
�l;�rj�!�	EXX����6,}͠דJ����g��g�V�Z���ڄ9��1�ޗS���ep��`���� ����3�G?�������O  0��~���Y�^cCk���%�P�'jc�#W�
�pm⇽C`���$�"x~�t����&UY����>��t�NV̮��\�_0��I���kEd9����jr$\}K�9����3�9�N�NG�;�0�k���\�S��޼2�
����]"e#�2S�)�=�B�󈜨�1A��h=-�C�A��cv�D�y�{�#��wQ��^>�q(�	{�~�썼/�$�6����
��S-��T��K��b�e����߹8�wY�Q�hъf��*ʮ�t�� �ٻ��9���b,���MGߡ��q �I�8��j5�DJU�r��J1��89a
�{�"�6 �{d�!R��)����
�|�!�$�&���]�h�C�إ�O�6�͑Ň3/�;3����]z6l�������D�>,Uv.^���8W�'&�9t�%>�y��@l�VAG��ݩ���A��|�	!��s.�"�tG���Ia^ nF���q���A:��Mx���ay���-�gK�|��~����סFc.�?Z�N2���q��H<�	��´ ���r�� ��ӏ|��Ľ�Mmt�
)�	:,
{yEh�	��Sϑ����"Ԑ�V�%X�o�d�,����W�!M�e.[yy	��/m��fw[�BW���TMQ�C3W�t'�����:9�J�2,���A���S��˷���T�Ч����V�,��t���s�D��[#���I��B��,�����T U�0̋������n}��[~g��zS��T�j�P�Ha�\�s�֘�9���E.�~�����+�>���<��
�wJ
9V�:.����RK�) 7�fr��7���%�r�7�{�9e"��#�L��&_j��L�j��2�n�`�;�Z��0-1����rKQ�1� �oF�#G$~�����R�kYTl���	���÷"b�%�PM�t�s݈�e��L���ˀ���;�؈ �M�ﶔ.���Hsܫ[�hM�:��*Fr�tlS���s�G,��1�VX�o�������5Vl[��֚���bF�8޳ߪ�7P�<g_��`����P?�;�pi�x��l�xM�hó�rd���n�6������~�i�Z,K���d��kS����Y4��Ɋ�דj4b�?r�U��P�}2w]�wi`�g�j�ҁҁc�&/VQ�%e�$Iva\a�6���3�	��e�ח׽G1n;"��
�6��K�s��؀�ʋ�S$���.v��!Nh�o�dܝl8�(���o��ld����wNWo�`(��GÎ[�S#�C�:0��&��]�Fۭ�Y3�/�p���P�;鎹i%�7I��wA����JM<)9���?���������T�$�j�G��hÑ��-A��RX�t`fc�_�Tg}:��$� w��Y��qֹo�,�h��ߊMɷ#�h��n/�
ƴG���͈fS�R�ɷi����ܣPB��)�d7T+�~���5���k��cq�T��ݱ¨+�k�S�=����<�(���ZhӜZ7�Y5X% �M1�"3�W�1O��uB�j��H*Cړ��Q�T:�qc2��O���������˼C�׉ʇ5}�L��K�L=w��-�IB������R){/jDé(�<�)4�����Щ����ơ5#n_#��� ��i	Ig ҙ˨Ƿk��I��BY�>*	h{��]|�f�y>�f�2|�O <�:0�z]�~#���n.�L��UQ��l� �J#Рt[A���0��40r|=uъҥg�ƍّ�µB��ڋ!DZwsj�
 ��;b&U�Q;�|�Ux��cl�H
��Z�B����ِ���p�s�XQ��D)Ē�F�L��~�a�6f�6���3�r%�+���P׏�%��N��$��0���G����4���>��^.�Ǯ�QH/9��G��_�?^�I�J�ſ�vT }��.-��ԇBN�e��ʚ���,)�ޮ`��?xT��o���uv4D����׾<-�)�$D���q�O*�.oa!P��M�X�705?���-���h�f5�vW#��F)���~�e� ����PT���Q\�G�t{<�h2s�r���M ����n��(�^��k��p)"�+h�5�G}�v�Kr�����3�����g
o\�W�U��g�
d�k4?����ۓ��HRJ% ��s^��`pۏh�+S��⼨NƊ��^�U��d���u3�1��=�{n�	M$�lj6��F�z�Mm����l��e&c�����CD����x\ҏ'��q���[�&h[!�0����P��Ÿr��?��-?�$�#�{)1%f�����)��~�ȿђ*]��P����׺<�-*O-���p�XB�Hy~�l�ͼ�Q�[�����PG��r�*�o�<K����>�
ABQq@�ꕈbV8<��%�e�����K�p�T���&P�H���A>�洅�P'����7k���\�&� ��t.�:�X�A�"g�Z�)M�/Hq�zc@��s���<_�r�d�
���"�i`W\��aK�� �[�z���#��ۅjcc`�h�����,P�HF�K�/�k��Fj�DV\�W��0�#��~��l�3�iHF)K|2�R�פ��J��i#4z�"�ӱ�l<Q��N�l��L*~����	�s]�YC�{?�h�4�O�<����;�:r<����(v���a@��N���|z�lц�㿝B8��)�s���D��W�}ދrOG��j����D%-142k���!i"4`?�j�����FeJ#�2+��9ʶ<������D�-�����F�Ҵ�;�d����m�2���ԏ3c-%%��&#�m� (8�mKl5�2��HL���q^�i
~��t���T��x��\�S������[Q!��@�Ԅ�Ks_�t����y�����҃f�ik����ew�4J�b"�f2�eV=n�*�Wߍ逃��(���d����)	�О:��r376(�b�cȼ��� ���F\��ưWFh�����g�$[�-B&~��	G=߱�P�ߴ_�q��EM��`H�#Zx`��bii�2����C�O=,? ���E7��&��@s�B��`��`9@t�1ԃ��:�an��pd.��J�k�����T�}�����ν����v۵_
+���_r�|s���QrQ
y���.XM��5���v����3�-�$m������F��7�L(j�dȱ0��t}���m� S��T{��"O�(u4:���l�͜k�,�
�bGt%h�'����p*�%�i�#R��[������!4`ɀ�z)vY���L�!lw��Uo�z��ryY��`$c�J�sCV���=��
2��9�3jy��n�Κ*?�'�tu�os���!+�e��E�U+Bxy�d�)�Tr���7ip@� �V��48���k� �J�Ҵǫ�گ(��_5~�� PTb|bO�@�U�\�����W6�j7
�y�Z��j.�Ki;[��=�rz߆�Z�qW��R
�Ē���k�]�R�v��Oǚ�A��z�'"#�����偾���Di[E�`5�Ld����å�RoW���#/R�}����r��K�Oy%
s``���a��-:�6U�:�<S��Or���4��%G�,T���szT\�j� �[��ElRZ7%��ٶhȾ@��w=Fݟ�*S���I4=��'�zC��V�oB�!��1�e�M���A�!�J���{Mj��ɧlV��	�W�;F�QT�e.�����עמ���e�k�^�(��[��p9ς~0U߿��^o�� n�\����%�(�{_��}:M�����C4B$��;>Y���v7�*���������t�ݍu�)��7.#��W�A�73�M3`m(�� �\
B�*�ܷ�"�L��Y=��Ax|�TT<�
Z+�S;凒+8��(ΈW���$�A�F��u���9Ν�%�r�{����n�mH�����L���/���g�`8��|� �6=�x'��5s���L��К@��yqi{�*C� rB����˦(o�Z#�����[I��g���F͘<��G����H��2�@�M ���[� x�4�¤�Ias{fe��x��B��z�^�6S.K�5u�9#�1���3{' $�])���܏�R�f+c�5��Te"f1�Y��1v��ʝ(1�`2p���qy�U]��J��u�U�~n���V��5�GMPk�/�ZAo��>C*�q���L�����T45������D��"w#a
�{�Q�u$����	e��ޥGL���/.��ǂ��1������޿��t�\4��!Ǣ�%Z�̧i��{�|Po�4�>��\_i��ͺ0�͌]Ӵ<-��B�-y��c��]-�[��̝=�&#�Q�	��i-�8�u�9�M��` .wg�a+��C���_�)I�^���o6�=	;�}�+�!Xs��bi]l�ۏ��{��꺐�W��Z�[/ �*g�*��6�����t%t�&vY���'� f���Y�|�7h�>�~�-e��UQK
��zp���V�E+�g ��P%51��E3�	�/���:�'̇&�'X�+�uނ�X=��9���e�S�
�o���D9<3�Mp�B��9���I>8<T�{ɚ�aA��;�(�0��в-��zC�+�S�<�r��a�=M��7�7�x 5/z��M�=�5"�n�J���^gD{�F!���4�01�#G6v��6�X��#�a�8���c,���=UUFl��d����/;ć=���Ts����^�a�w*oQ�gP�	$��q�+1�1<��(�e����2�	����� ��@����}VinLί��Z��OˍU����x˒)2s�7�'�`�v�ݟn�5�@*� �̝��;�Hp�3���f�F��y\γt!��&K=�-�=��>K;�O�D�)E{�b�_���<:�н0{���3�+��V���:y��]�D��0ߜ�P �+��3���Q��K|��E��p�FFه�3`��s
��̲jGJ�����g�w8LY�,��������?���g����"�& ��%�0�#��E:�8f�<��D�1���y��Ȼ��'!pUv�(ݐ��p��dJD&G�]O��~���=��~hJoK�'������˝I�C���W�-{���JD��!�'H�nI��ؖ�?&C+y�}	s��)�vk�$��
~�@�����c[�s��>�i��{����w>A,�PsNiEW���qe��T��.�E<=|�!�@��~z��e�@ w��܂Rc,ۖ�a� w�� �u���|���\��T~�XTs�\+��Q+U�:�r|�B�{������z�� %AD̶����w���4'�ú�qrT[N���?�#z�ɇ�I��BQ��2�}�C���v��%=q=�ߋ!s�ɖ�Aϗ"C<��ȣYm�{�g�H�[��C.��54��RGM����pikը@�%��r�����=��.P1=p�ZE3����;�ޯ�?i˻��l]�CNd�Q@G�XGݳ��#��i�|�s�YRͽ�ʫ�rcƒ��'�H�8��Q�<	���U=E��
���U�Ĕ��b�䞃�L���}�a�����iT���dm8�ᜯ5ga���4ނ�dg���l���p3��.���ދr��u� k��P�uI��K��7q�'�j\V^�M������� 8mC��&��>=����M��3�J��E��I� ��)c� ya[̺>�Tph��dM��S�7Ӹ���&P�*�z��u7F�t�֎Ś�h;�;��ח���BQJRC2�