��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|>�qT��>��f��AR����$� y;]�*\uȴ���ԉ)��`���C]+�g�tpgV���$�[@��Tx�\Y�͜��B
�ȹ��3���As���+y�]i�hHRi��s�J�O���[=�t�'���<�[��K%���j�߆?y��-(�-�p��Y8v.����Uĩb3�X��J�� uX*�J�s���S>�iÙ(6���[��ô���_��w��t���/��D�8w�Fg�S�va�.&�~(�	Ǝ�rQ���q��@n�i���.GڧL���a���)���'�b�r����ٌZi�6*5���\:���C�4EFrYC�|�9�����d���tج)�uT.!h�A�l�=Z�	T\pų���G��73��ZN���F�L�[���4ڃ��A���X|zx{�Ծ�%�E+>
ym�������LM�ط4�x�>p��~=#f��*j�E��S2�џx� �,-Q���"�й0�͚���"Q+��n&hY�<u�#)6g�JH���!ڋy`�n�x�n��%�wh
'+�� gajL&���e���
��=%K�]~��~��;��ّ*
?&]\ϓ��#h�S��,zs�+��4�Nd��N.^v�(���J��V���_=-���3M�������7�4����p4ڝ7u`F�@y�"�G�����N�Bj�����4�Jv��͂F6p��6�n���c|uV���!js"�D����w,sU�7� ��"<��P���4~O�s�w]&Y��콃�[���9�2&0�=}��8AK����&ӫ���z_X�r^��3o�_��F~d�0�fȽy1e^������&՝5u���7�tl���wQ�B�x -�n�D(Q+��W-���)7	̙$�
����"�d��6�wr���	+��K�H���ʑEd�WkL��D=���-�'���)�>m��[���o�|	�!�8\׻��䔤�< �9 r���s�eh>)�x'�EG��p"���qe���1C���$��������������Z�
���� �/��*�[q"|��٦�vL�Q�Al�PbB@g}�6I�1���w�p'����bx��.�򻷒t�˅�M
�o:F?�r�����26�e��{�T��"Lg0�%i�J�g��0�>���r�Fs�Y8�:�O#�&9��Ls�v�_ʥ������e�'��P���r���$O� 39Tg=�C��V�_�t����$g��Gp�nY��Co��o]s�ji���y�/
���=�]^���o`�mN#�ta�_�H��j^��`�Ν��~��ڑ+��~��n������l�]lf�S�RW�ܶ$��i�������SD�B���t����6�SOFs���:@�Gk��hTֳ�l��h�
$����ݘ9�y��j2b�uĀ��VP�v�o��Ԛ�˩��fe�\L��ݬL���4aGw	�G:�;��Q� Ĳ�om]+���؂�k��������M�O���},�&���mFc=���!�%s&�w2!Odkﱱh�1����~��P9��b8�(d�%�"߽u�ɖ561w���,�&��h�FL6{TO+��;O���
$�䜑J�wmi{� �z��s�ps�!pQ�&�����R-��J=,�\\I��@�X�g�Uש�U�f4%���.ˇ�~`<EA��P�e���tl��}��z�+�Td��������s�ae3��w]$wQ��O�.�J��	ӕ*�J��^�<]�6-����j����,��歎;
�R_�-	����T�� &GC�f1�9l=��g ��A�p�F)z��n_ ��z"|��N��!�Vγp����<1�G!I��u�MƯ3'؞�ܛ��P)`�JZ.��광�G:-тv�:FMls1���{��1�٢�x)Y'�JeB��~K���*�a��v��x�\�o+�Iv�}�k�r��^]��@J��U�?�`g�ͯcJ�a�.T7f�Ij֐_D�I�iL��"��}b��%TֆQT,��+F���hZS�Feq�WXҥė���Yi�t�F{���IoKg�5���M�u�A���;�E��.@�l_��1�Lc9N�w�h�A6��,��^�u>��ȡ��ռ�%��B�����0��u%����R_�o;��/���Pk�D'�SA�(z�!�߅K ���y截}#�Ej'O}����sc�x:8#&p�U�t�������} �5�F�g��݌��Z#L�(wo��k-f r��nH�W�{g�)�gΦq_�|:����-k�yC�	j�t����N�b�[wfDx��Q�C����w�L��H���Oȅ6S�[4q"}�cXg�í�ׅ�=�-Dsv6� Yj7?z��SR�����0<���:��) >�^I�,2�@�Z�_wFd��_�"v�>���Q�9��\��z� �>o0�>��r�":�OF��ֽ+$�)���UnKџ=*(��p��9Ua�����X�}N%7�MF|�i�"�M'@	��:(om��jd�+3�>��OSD�ޘZ��ޢ��\Qc���p/�z<5_�dHbD�)�3�- �I����o�'��sw3��/(��y�µ��P���U��4���]��Rs^�xR�{F��65Z�//�g�
v<B��%���2`��'��NA'�}R�O�=���\l�6��2�;��m�oK�)`���|P%�ҝ���"B��sR5���r���T2cx���6qV6��.�����9ܖ��Ch�0�)1P#B\
�.���|��[0`�{&h����P�v�����yf78��Pdp��]�_�=����#�vA��-���(�ё�������&�"��Ban������w	��v>��B�S�3P�V%hy܆���������8Z�w�c)Ҋ�&���^�=��ok��t�T��T7��r�Y8����.���yb��ky�+l7��y枨W,�0���p-�}JE���[R���H4ܿ�`M�3����،_1����|���.s%} `j+CXR��@U����4�۔P�X��#0�H�N̹�}G��������s��9��Q(h!�NT�!Ob#�_� aG0ie۵
Ӡ� �0��EOS�[�ہ�vP���1@���ɍ[RH�P@Z�>�����j�A�?���#�wk����W��qH$b���r��9�IPId�L�a��Ii��v�U��0�)$�;�:Ⱂ���b�Tp�yϦV:I�I#��B1#�Yî��j�P�~]�gftP{onj�VT����W�P���D�f�C�z�q)��b;i�_ @7ZՀd�0������-�+&�^k�	nP� �����	2Oi*�[5�m��?���<$%��������9N��5��q>_����׆�A�.vV�  "HqYv, "La��-:@�P��dڷ��*�F0�1�i��y�����kX$��8?0�[&j�8a�:�����Sk~��4��۠w�b˖�C�u1����	��XLA�s�Y�Dw��e��nj�Ç���kx[ԗwC�ʅ��i>��9�P�KW-�߻B|p�����>f�0R� E��9��X>�P����̠����+�jb§�b��r�4�v����O,S�cpP�����B�=�M
��/b�v�� 6|�1_Zy=�yZ&��6��0;]G��P�c�*��3Bt��'06^�1�sʑ��(�)�j}܇���Ҳv�M/=�!�.��b���t�^��4]�`�㥢���u������竘ie�91(~�G��SW����(� *�ORz����u�