��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_����m�e"kxu�Uٲ"#oB2�-g�j��h�p� M T�(�P�+M��&�[���+ǚ��.n{Q�̅Z����&�;3j6dED=�Cl���ȸ����8�^+����K�\u��8���f�u�$$��LF���ꆶ��xV���*'7}�� <���.rQ	�+ed\���M�����$0	���I�����B�<�.�x���1�\��ֵ,i0#X�;s�djuM"Y:����&�H80k�_@��B��r��z!9�GWlOC���C�ݓo������i*cVg��F��	c��6��h��^�_a�~j6��@�������[�0׉�2�+7�Զ4ۧC�a��e��u�v�a�R<���+T�W|Ės�U��Ľc}G.jWV�(*P�{�.$I��8��mZ6�C?$��!l*�0J��6!^���]��.	mT/5���lo#�o�(u`ܓ����zC�A���hڔh78��iC�����l�b�"H���Q+v����j�F��	�f���E\'�V�aI�}8�x�[����Ņ�p��������2�$�X��?v� �fK��M�cVb�`���P��J�(�m"�� +��{SU�V��m뫽�^m^ml�S�!p�(ZiG�V�ϳC�| �h(���.�G�L�X�p�Q�<�6��ٮ'���4�yQD����R��������]��ن�u�*~��P�Z���\j��(�u��N(�6Zp�kع������߮#�͛�B�a���6"�)�D����Pe���ol/�.��m7G�존K�Xr��1i~\�~�.玝��J�]�����>��=ވȯ�}�.�C*<�b<]g���q�����!m���b�WS���g��(.��U���^G-//�nJ&�Q)PB���A�˙��<c�r���d������&��Y]z����v���l-�S��K��E �,�?'o����K�݅���ɵK�K�]�5���`>7���CA)�b�7�OvP�g�_���/��L���A�[��ʒ�&l�]����6a*�n�R���8䦖L��i��t�O,�&L� �J�4�"��3r��1�������$��`H�w�0]�Z]�^�%��!߳\�x�`T�M�yE�Ѯ��C�WB���+�l|e$�=��mH0�v`�ŝ6�:y��q�S�h�d�\������ʨtCG�Cc���g:��kV�/���I'�~���"���$*/��p	 W�`���s�H��ߟB��r�4�ţw���,�r�-�e�8����'SE��*i=(�7H�:�~FЕ��
5��?���Ⱥ�	�>��e��Jl�-G��kPaXE��X��Q ��S�S�k�X���]���cE�&�!��R��@]�,�MF�#J�/y����6��^�d��x� _��	�x΂ț55�����a��3Q,�������������E�F^�FҸ�ewR���|0�V��{�Ż���#��>	j����B,�ߌ��#�S�Q5�=���+Y��>�"���%�!��>���}��Mg��j깸&�0��%α��V���
9�]q�e=���<lV兩s��˓�L|h~�U���vݴ<�y�Q�%����J�b��nX�L��J28��r��A�eF�_���u j������Ow�c�4�YbM�6h�Mnw���0@ݑj� (�R��}�#��:Cc��dg��?k+4���52�	�k��z�u�0#4'>�\K�GR�7�s ��@���Q�P��-��8�,��7\�����E�C�4!��G�!�W�u�҈Z��Q8i�i�[���Nd)������>|C��Oq�<���m�̄^XK#X��ɪ�k!�ʥ��q�-����R��A�����w�T=j?7��W���#,��pw�ݟ3}�O�@a����~ƕ݊
|�sƽ���D�^]���Zzq�H��R1}>%­��DT���3x騻h
��B����|�Lp_MR+�&s�c���"c�YK�u$�оl��쌗s�</�&|���h�u�\�F`jɱ��#�f^FM\};�p���6���R���wr������\��8@ ���i!:%���M�L&^ns���|F=��J��Zsi��XJ�c>�/c<��k�c��9��Kn��	�xl���a֦Ln�+����%�pݰ�<��o�7��$x%������Á�& ���K�g�z�0�f���`�h�����\Y�V�~쾿�~XJ)I���)�l��t�ƿ�[���R���,�5��(��arj�i�-˨��3�	�y��)��Mf˦��]���+�{�k=�A�S���J�u&9����E��<1���"�M�D����8yx<P3�җ�5�#����F������
����JA����O;J5QK+?X�8��zJJ@2�S�� W([�+��[��,e�[L��&D�ޜܽ%�F2S��xv�h [��Ud�s�0���p�"�7�bp�`2�fA�삤�A�i���BIaÚE�Y�]�@����@�� ��A+�M��]dZ���Y_���9e�y�,�˷;�_��ś�U1�����Y�*!'� �6�O-�gx铔�[�Q�������M����Ϭ0=y� &�w�9�;<qdW|�d���8:Q�� �"PP�. �$d3.�.G�i���3=3&���͸Kt���)}5w-+vv�ɂv��n%�������T%cr�s-��M{M��OD`��s@���5�T�iu�U�߫Օ��Z6���nٍ0Ӈ�ؠ�g���Ϟ��c�W�,�Q�;��͟���@0O�%��i�5Nz��t{