��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�"��F9s�`&���a�oq���F�g�O�]�<ݲ����eCL��D���{�5��8̝DFI��Zp\m|Q��
�}�6C���UnF:<�jΈ�2�����<����sf�k��,jڙ�����2��X��Ss�HL��	�������+g?���N�Ż�����|�v7�{M��VNB
��Rs�゙�Ld\��X�'��R :�J���^�����kMkx�Q���3!P}�e����d���f{��@����S��>���4{��ת�AO�Q{���cR��G��u����vſ�ˡ�;� �-���&Ϙ��\M����&(�)NSF�#�%>���p�
e,����l��4EL$�ݏ�Hmڑi��THIհ�F���}u����ݨ�|���@�P�-�ͽR��PE�QO�<�$9c��͡l	x+vKm��w?9O�C�)���&AOZ ��j�Y�H��Ӷ�O�\V�d��3���4��?PBOB�f��S1U5�Pt'4�?և�*��*<���"�VQb|�C�O
M���Ze���\��=Q,~��w6$��ֵYT$V^�FAšE>�'���ɞ������-�)����	V��]�\u�jR��T���Հ�ߛ��Q��Y����NΙ���q��(5n�;W�cO����(�V����u����*�t�7���E���X�6������C��>�r��!��e��$\��"ܦ�R�?��	�3�+6����]���MT��ĸ����0��x{@����(I�����|�ZΣ�~Z�e5ջ]'�"2gc!��Q��S�,��3����Y���N�J�'�m��WvV¸F����G�n��_���,��2����������!TZ��	�ބJ��/��Db3�,""=�r-(>�un�!b ���uyn� �+\�/�9=;Y"F�P�aH��aP[L��D@����n��Lͷ�]��^��= �6H���� �[#�lI�7΋us,���3�
�d��ɱ���S%��Ib"�K�#�a�FԈpB��Ό������h �X�N�1k��ڊv6G�T���N�[XC-LA��6����xR�����-8Б�AZ��24Ӱ���"�T��#C����!�P�rѕ'���ؠwY�K؊c�_�i�W
�Nz+ѭ�'�T��Q�i��!/U��ք��³Ƣy%��{�����o�m�|����������/6b�OGW��Z�l�v�(��̦8�B���9�L/�������cD�0Pe_`���47�ul$oʨ��lQv��Q��ۧK �r�	���8/d��pL=#I_ڬ����-�<U��p�N��+�'��u��
��O�A�Ͻq�z嬍���2�
'l��_��}��*Պi�U-g�A%���0u\�����v�Y\�����	{urs/��EI��i6 ���[}�0�.m3��k�;�N��^'�u�J� ܥ퀶��s�o�,���r�f��^d\��,o��OM��׫�;S�I��}�|�j����`��]�!�;�-&^�+}����j�p�>)��؞IO�~f0��m�ݣ�hC��I��i��'�'�"�Z&�8��o��V1�g�xW}A�aOwÉ����4^c��tHp�xW�������H��-2[F��m}�٬&��җ�v�*2U�4���"q�ФG�1_��u�`�R�V�e瓙���v(��[�����EݔQ5C�2���G�T�id����p[�*�����ϩ�XHƉ��n��U�i e]�E��@�'�/ٳ�*A�\ፁ��x\��ob(��r����_�ՠ���)ea��ϱF����G⽆ ���`E�j3���C�j^�jː��g=���������6�_k��/�!��J\ +��%I���D4H�1��V����W���M��~^��ӿ���r�C�4�*�A��2��f����#ܼ`����2�Jd;H|y�T�� tN�ԟ���d8J�)���l}D��s	�$�m�.�1� ����$�7�2O�4Qd��l�KAL$9�|��F�MW�n�@���#�
d\���@7m�PF+�b<眽|�z:)!j4�Ì+��������<�	m�L�d?�@Y;�K��>��D���U�&	A䷨6YT�~AWhh&�sa���&�b[p�C��EB
�!�`/���1��J��GH{�6�Q�\C��0��������E��5.��B�hxC
� �pΆ�Cl��Y���p�dH�>�2/du8[�lѣ����&��QX���,������%6��!�r*�s:,�����5�������'P��񵯥��`]g&-P]���%&/^bW�����n��q̃�|����GFmb��/g�r*Նqc�^��L��Gh������+��a�=��[Y4H��_+�@_�\�����/�I�a�B �IR�f�R��%����>�W'Il�U]�f��|P��;�Ꜻ�C"_@w�0L`�/X?�y��T*��X�~��6�]��?e(-{SӢ���u	�N[���߬���j�W����P�=E��5*W������h����)8-̟�}o,�sLx"���}\b��L����[��eg�<Bs(`����x���
t�� �#�^]`G�g�i���4��X�8qI�23sm8��b����I��3������i��_N���=m�����d�� ��qXۭ�B
�% ��<�:(xC�\��n3��1�(�=�EmM�N o��T>����53�~�����h~9����Ѐ��5���V֔N��� �o�+�K�=	�a���%>3�Dl�_j���s���Y[>�io�=�br"y]��$$U�*,µ��WFD*N�Pn,�Q!-A.�ٕ�u�P�D���z��Xl*�}��Ј(n���%H�Qy����������B����fxd�?@��1ۧ��W�I�r8�:Q�0�3�2ݿ���@@�a���l2������BBA3S�$�6E���{�{Ӛ5�^]�!�]�A�WЋ�N}#Cb��9�� ���i�D��:�
��QO
�Aa˝��(!�N������`�X#����P��V������9�r{�d�h�j���GYHn6��[�s_~�Sv��_�ЇU�G�J�ݕi�1�
�nB�Ǚ�Bf��������@�L�,,��}X7Մ=F(_\�k?�+�sx���h�ߴ��� gsk�n�=v7�X�Y�8�8{�?��`�����̯�jvZ2DFwpd$���{_j�|�6O�/�&��e��r�h�F	����(����%`�\{b��HG�K�!�7��6gl��L�桩co�G�2���^i̵�[�W%B ���\( c\.c�h��qIfmu���\@��aVY][é��-uQ�.�\��ڢ<�x'�#�{ơ����]yH3��U��j9�:���E@Q��7uNʎaR���Y;P�/H?�������r+�Hv����0j'�B{���5ޔQk�u��c�eױ�.��� �Ć���[8ȓ.'���jܐ?�,�7�o$�%xT�{��,�����1Y�޼�U��K�h^`�C��ZE��K�;���@آ�\�ITX����7t��}ǫ�+��-�G���u"��_W�)��bɚ�2I���%�C�1/7�+d[�F~���3������V-�����+�hB�^e����gW���	��.�l|X�e+�ށ>z��������������?��H��h�gp&Z��l�G�3�GXml`g���&^��i�R=�8r�F�cr��/u�\�&2����$.��Sȯ�Q��+����*k�(�e��T� )ǥ0�7@��n�W9����r�G�w^���=)Nj�m����s<B��L:^�H���7	t��>�S*ӂ�e�Y|�6$��ڢ�u�r�6b�b�k;�mEW��M��RȬ����,Z�̼�=�@�M�%801Z�0G�W� ʻ�4�QVϥ���Nn��U�0势��0�]�c�����2\�|���>[KHT�<iƞ�@��)@#��ځ�'��k�eb5+?�J����O�B��w����Ӟ�c@Ϧ �/�3��%r�_�U4(7�ugk(VA��&�B�q��8�g�<���Y�V$��-�CU��4�{}�x�֎��Er� >�a�?Ȳ|~�;L��+��Ǯ�h��%�wo}ጲ]F�h�LI*DL�?l��T�;_���kCl�x��qq�f� M����\�0bv�	�]�#������0ؕ�G���(�I@�<���%]�t�L�
���i1� !0tAj�Q��)��"P-�(�ZZ��ex�QK�vy��1�l17���>���b��Yf�I�݊�������+�'1}NsX�Z|t������G��a�nu�n���J�L+���jz���(�K�O�J�;�1D�(e˪���nm���-�6I)ҫ���'�6Ťr�j��H�a6��:'L��.Jv/���cW��������Et���G����n<(�fN���ٱKx�.��٪�%$Sr��?#V �`[L���hJY�S!��6w�'��hKyλ�~���N�jC���LB���y�X�Pq4��6������ѹ��,I��-�3�Į�\G�$PיK�1��5�tsʽ��@4�Vݲ(�(����G�@����{�0��1T�3�o��fU\�vB�"�;;SL�̆2C���g��Z�xZؾ��Q#}N�M[���1H1�kOv<t�m�K����C����S���i8�у&���8*�;��7-�����j񆂯]_���F�?#͍�'!�#�A�C������֫ݣp�嘢��K�`{��>K#Ԧ/� ��Q-c����W��P�De�T+�j���fR2�J$�K��8M�yݸu�\+QmPx�g1���]�]���8;���Ɍ�}3�oxPۂ0���J-��SgN���ڹ�4����od�k0 N!;Q����x���'�/jj�(�7���I�gF�1�]uv��9�o�� 8LF똯��OP��gM�~h�ť�vV�� ���;�*����/�mG�K}��Z%�2��,.l
H )����"ƿ�n';�戝�t[	�9P�p��9 �����E�Bg$�3�D�zt=�O��[HE[���Ѻ*z�%t��QD�Go_�b���6�\����U�Eb ��0鴍���GNV�#�?�������6>���yj��+j]Z]i�N��xjۥ^�����HU4ɢ�͵9uDM���h�
.$A���1 15����"zS#Ά�e_b�a'%m��q�;��������Ȯ�;�x��*�:R�/��7��̻����O���t�{*m
5�>N�OP�}+�����ˊ�g��m-'�}�����)�ti�en��P�;a�|�k�>>�:f�)��Q���% ���?�tI�k��'z̀E�Sy���ʌ�ş)�eɼn���`]X��"��5�:K@*�����P�E��'� �g��?F}za[�L�$(�気O"EJ�^;�P���.)��`�}YE����>-W-��ϝ{��ED��# ��u�%�͡s6ܲ�ʟ��T1Ć�F)���`�<���f+ӡ"�D�:.(���~$E��j.&�Ȭ����&�F!ja���EI���vRM���5(߬���0�Gtl������8�H�#u%*р���z��!0��I�I����M���/͔j��TD��^��_.~�+x�����%���y��u�[t��M�sKU	��U��u�b�V�[�r,x�k���Lk�tr�#b�ɿ�G��cO�)ҁ�،��6�#@:��rMI��u#[�#�mwU�k|Z�S���������J�$4��ё�����q��ꨵ�<��|���Ryջ>�1�߮�X�{J1F�_�c�U�Et���!���>��j"�u&�cxv�9��U�6�9!1�t�Zu��F�w�/�1�}`��Ƴ$����\�{׫r,E�xZ��֫�5 �u��w�c��W�^�����c�S2�P��bG�XkK������`���@U���%TK��3�#K�汣�e�s��
�-�;O 0���UR"k��h1L�֟Z�D�D��4��ŷM��p�@��~3�:N�Gf�β�h!�"��	v��OHR�M4i@�%[J��q�fH8�Z�Ջ�9���`
K���&�B�	���e���>�6�+2������C��J���D�Uh�'����]���2���9�+�� ^�x�^E��J��+�#�����Q`GçL�2L��wY��Zi�!�L`�����������^��	�o�q�ޢ��Z���rD2�h��#�P�cp4"e��\�+��W�@DP|�kn8�fA����ש9p�ʌ��|���G��(Q��27c����o���^.D�\(^$�|�@b��w�6ػ���g<z�W���q|q��I�C����me��1�<�����V�E�i)������|��'�eI���UjZ;<�0�m���O�N�d�7� 0(>�����G8`o��yb5���M�1b+��3]���r�\bR��:N\/����E1��5���DZ/��(k�BS0��Զ�'������x4/[���`��qw�xnx}�R0��~��{���VN�u�����ѡ1��:�,��f�	v;$��3d7��t}�2Li*��TI%�l1�w������=w���#��Z;;,X�RC3�+=q����Q�«z��
��P<m=��4 B���}z���I����@ة��Pᢙ:��ÐvAG��'�܃�G^!X�J�i�}��~�N�0pD���j�i���4�d���8N�Q0�3���"�f��0��^$���A��9u�%��.U�N $c_o�8�\��@�
�o����!:���ZI��h��+OIIž^�|fy X�˃�ޠ	4��~��a���1#<��{��n	Tn� �]�!AC[�I��W�)��Y�_���kѴ\�o�xC&����Y����0;�F�4��Ş[C��J���$ X��es���n��a~Y�:�<�ʣ�w�:as�4�x�29E�������Lb</ݗǼc��5[H���Wm�lA�|O��Q)n���z��,�*����)�Y���|�6!&.�yۇ}�As5֒�3��������qс�^���!��T"�)��1�N��
R����#;9��˦���=h�9�LN8mIi��8�IQH6_�2��,�	`�P[^��M=�I�tgu5&L�ְ�3}^i��/��s���r���|�:p�%�<���HU��A���(M�"���c��~��o�K�(���U���L���L�+k��h�P�-���F��	Ө�0Q��$}�5��}�c�\*ށ��0N�_`��	��{v�58��OR{4[{-;� �>�y��}o0j!��^&�L0�p���vׁ�(��� R-i3���ph����c����������
HQ�(M�5x��d����tn��o����J�����ρ�рԀ�o�<���K��ț>�i
D�dz�y��EىT���'�3�NT�J���as9����,X�zl�!�7�1��(��aZϖq���>f�)HF����xڷ�Z)�csמ��m�6��M���UR�����v��0����ɩ�Q��w���l|\E�Ť�,�a�Bz�l⯑��N�Q��+��l�70'�,� �{<�_"�V�!��8�(�&vK�}��nuqqxix��0\߄+5\"�yT6�$�'��`�K��x��/��[-�������
����R�8>��	9�lݡ������X1������j�%�� ��`tߦ�8������% ��乔�玏o��Q���G�FƅV|����4��GDCa�g�M~�ru���e_s �+U�݋�N�Vt'/�ŷ����J��Jw3H�~�]�á�P��T�	��e�C�Ŭ�9�q�7I��좛���b�$�k��{��,����S��E��������4���'EyjO�����W��O/.���F�$:/cH��߅��6�čR�U��������,�+F�o���QT��p?o��'���5�6j��,��j�0�mޱ�]`
%��W���d�H�&@�E^pwE�tA��^ >Fl�pqB�
�+F����H����O�	}��M�/���ڙ�{SpuEO5>c���4\��d ΍"`�\�vݛg�ݘf�ŦMYȹ�EB�ҋ�D�1��jD������b5���/�E��.�o���>��G�1��"���W�8�s,�=��G��$VYPbc(A��m4�! �vU����^�/�I� hο�в�^.P���Ÿ@L�i�l�LQ�o�����M�+QxE�q�j�6l�1j�N�V��{����pX�+�s�C��B|��H�(>2~j	ߤ���RXx�c��)*��W�z�"�~1����橱����	$AF,(z_cσ�N��zG[��#,=��\���g8r�5mL��#]�8`L�k�Zw���Q��u�3���p�\6sn�z���>u+�O����x|$��uy�&�b/&��ϼXuZ��!����6�(���������	+X]!H���_�hen���k��+T��YIi!#	��r����a���5�����L�s�.�6�&Wp��>�@6ԫ��"��gT<Yץ�h�8?O~���yͅTf��Fh�v����9��΁k��������-W�K۪U���m��7�ݍ�	���v�T9�{њ�`0,�7����8C���3=+�cށ��0T�ZR-�q���x����.�a��d��/L3:Q`&�l�H5P@��A.u�ix��0~��`���LW�J��o�"����=�Ɉ�)�yB�0mE,��PY�D-�ή���ZM# /���V�q�Ij��TL\ɵ��]�����2��Fc�$��O��&Ȱ/߃K#��ēŵ�KJ�b-,ˊK96�CB�ӏF����$H�Tv��6��fK��+DN �\�vD�НM�\�-p�FF�]z��(����7�f<�r
���9c̲8�7�q�F��<�V��5���YafmjOr�L�;�<�r����L[m��D�z��m�}v(����m&��R���i���(M�z��w����w��<��C��YO�2�8GԳި?��J�˕�?��vMY�zH�6�&F�Ɩ��=��M��heԋ��PT�G��IL��2������ґݢ�W�`EOqb�n�!�tم����f$l t�+|��Ûﱮ'9��xu��MI�MĤY�Gcd͔r6z�^s����7+�sF8�e�O,�Q�	�M���/RF��k)h�ҵ�'?���+�x4Ӿ8Z1��������5I*�����i�M"�^q�	�
m^ *ZTT9��|[4���	�����|��%7����rqt[�gϻ��v@��l����_!gz2D4?�.��ȴk�����w|���^|Qv�T_���Y�鏼�G��j���\����:��&�M�����A4�O�}��e��k�*mO�>�ʔKv��2���M1ۮ����_+�n	6!5��"��#��}��b��:q�F�Έp��b���Cpn�*-f���V�*��O �_����;!��X{������lݕ���;8K!<Ƃ���Y�ñ����EY4P�����s�B�����!*�do�9�@
���*P��Y��P4�)���7L>(�T���Ȍ�1� �h��CO���.�����h]����|8���������\o�#��vF3��õ1G@�]�%��Z���8�������/+���Qy�Oۦ^�~F�"&���A�{ð$��K��;b��uUg�"�1��t\�?��2~No0�g�З;1쬌1/r��;Hզ�w'=��V9��|y^zWQC�ZE����B�V�]v��XE�d�HY�~���i�7&�-�xmi-�RR�P�p�����Re��������������f�'�r��ǉ�Ȩb?��%��h�m��EB,�C'�ߦN��@`2GF�㙜T_'�q���+���rBTI��q��({�,1!�	���C"NK�f�	m�����.i��̭�W�A� �AO�g���f�
��b��9&WNGKO�^aϰϣ�M��~ �Hv���ɠvS_O���J	�+�R�U�������P�����,�rS�'���w��� æ�Utݸ������#�d_˞�N� ;G.�	�
����Lb����[_��1�Ұ?:7L�e��7�d�*Мi�wxɌ���Y+Ȍ�̩'ʝ��\3�3.^Ӏ<G�9nK���a8{������_鴭>�}�� �a�nJ�:��NCo��n}����G�G�v�Ja��!�}O	DF��� �ܪ�����4 �n�hj<ťM(L�����xj*�<�܊���9�؁vH�d�ўZ�<}+�$9����Ƒ�IE�n��.|a�����=����޾������!k�X�ۨ��˔�����d��4m�h��Uu����\�6/Q
y"���L>[�@5oF��dwd�N}����.�Y�}��Ƕ(������]��b�_��#k~��o��'x�1";>�0!袙	ͭ�
 8�����_�v���	�6us���� 0��j}�?NN�S�LB��
�Ng��N
����3e�&��#���p�Ŗ�ua�>�)�U�V>�2�ًW��b����c�yή��9Y����W��=Z�6�`X�_��>1 �����`���NE઩�l��@��q#U&t�k�"�O��a�'�߸v���-�/M��!E�;��C�pH���¶h�ڣ�L*7�ے�D��f�>኎ӒÍ)���{�-a�acr_q;��<��J 5L��P<l�cnQXH�:ON��lfc���l#g�t�4���{�V(�ST���@/K�?�a��ܔ+l�O�m�_h� �#����6��N�w�|<�G����]s6Je�'h.H����V�g�__d��N�*0��f������)���*	dN^C�e�Ϯz��-���yu?o��R���=�6��kC1��X]6[$ U���$\���w�wcn�������O�z@ĎV�#��9��h8O����y��7�}(�mˈW��+�
2���=$l��`�j�Y��(K�P� �0�Ft�}�j\��7�R��Me�ю>ӯ(�.+��r�g-�o�2N�}�k�iV؝��H�hM.�q0����W�o��a8�h�*�)�y�)�nǼ�J�H����1;"����go�w�x�^p�A�Gc+�DK��e���\|�1ې�5�&��.b}GE�z?�s��RӰ�Vw�WX�W�!y�����K�t�0�S���Eڄi�F�u�n��1�����V4:ޜ�V3G���>n�*;�M������"����MQ�a��ѽ#���J-3��"�5������8p�r�+��a�R_v&�[蠽4�I���X��or9�`���~��{�(;�$9��Q��� ��Z�$8v=����7��̧�X	b�t>%cj7�&�G���{J(X(���Ua6;}�,o,;�Y�\�YM���p8�/�)��02�1��K�,�\��R�b��f����!as���w��4��n����#�@��z�������u��>�8u2hw��{>M�.�>��8�ވ%���s���ٸT;>�?�u?��ǉB�F��QK�H�a*�f�"�8�N�,�R�n[�YA�R�g5�������A��2�V��*�]g����l��a�����B��x̰�.�K�kq����ߎ���r!����ݗ��d[�y�l�%�%:P���ʈz�(��p;y�[��l�3[�������'���U�ӧ�m�����_�B�q�]�]e����'�'?$7##O|b~�f��â7�:��5�ԛ��:�:�&�{*HYM�%~�F~�<����
��H�۵���ZR/I����y�_i(��Y�ֻV���^D�	g�?`�b���M�4Eڳ7�����-����EBr(�Ib}v� ��v��Ni*�,޼���VV�`w�H^����`l����F�N��3#��Z���+�l�;"Y��P��T����Q��а�ck#�aku��ƕ�A��C��~����B5�,qI�qľ�H��)��X�h�t�q�� ��t�US�rBt�K>�ǩ�<�7"��΋�~
[�u9>o�#g��0Ȋ=Y%��!��d���l����0�iɬ��B���Y5#�y3ɑ�����:!��]{FQ�Zک�����ɉ�%�FpF��cG�m��mM]ܸ�`�F���3���M;�w�<��b��!,"w<��@?�����@?�X3q�~�ϙ`,��mAQ��*�o�N�����Ԍm���#"jJ�˗���Q�EGO�Z����P�Sa���c�msll�g!V���Q�R�M�F��oy�.��)��ȏ�3�%��4��Ȳ�قs��4`k�7j���&�Y���ޒ����:���4�T[��0�G�Ï�����Ê�������&O6���ߓ)��F;�Cd�����kU<S�(�;�y�L�*X�k����c�Q������7��`�ߕ
ir$~�f??�W�`���g1�{`�+h}?�Hh	vf���>��@��؁-g��준��q��&�4ԭӋ+�M�����z��~<�'%V���$�S�C>o�?�9_�?��K i1��g����z�}Lʳ�r]"����Ejӥ;�tye]"�4Ubg�����h�U+�[;W�ק5�����{�x?8`��efi���Rw�g��ja��J�����Q<Լ������汫gh"+�j�]�lG5�$�c�\Vے�2^ۑ�KQ���IS�24�]���������@6u= �YB�F�'�*�/�|z:��jt+7%�I~l��R��jB��,.)S�b�/*3z��r��3`������qx�U���7�ZgS{áG.&�[
U����������xe]v�)���s��E�ԵeR 7�\A�;����X�����W1�a�G������4_;�-��i����m���o�7d�{�ƲuU�s4���d*�R5*-1��ğc6cL`8��r�����_z��>��1�ᨯ)V�6^cO�S��p���!QE��e�5���.�f?�*HI�B펷(�I�Wl�;{��������]E/`E:�� ����Yɤ�Ӵ��ߐt�T[�����O�Е�<�DM:��K������_c���x�M�|��7�j
��ٜ��?����>��֊����@P����َ�8���F���ο�Hh�~��?h�YHAu��^7(yn�R�Ω6��m,�@��5�$�� ���)��ApʏzH�'{*�t�Mu��X�Z���U��df�?:�)4��u��`@%�V���H(�;�hpޔ��ҫ9��^=���`���ǡ�8�th�FN�v�C2 ����aq7Q6&�<Hᦀ�F^=�N���9��O*6�S���s#��Nwk؈�>;�(n#e�0]�kʼG�ԌC��j���)k��e���Z!���;R�	P�ɧ�����U�'�Ә=�,�������AO=o�tf=���/ٝ�E=���9���ZI���0�Hu:y��cx�B�,c�C�h���ܴ9rAT9�j~@0�Q��B����V'�~O�_��M�պ�J��!WG�p��ekh���nq�[��R�+ն��!e�˯�nc�z�����͋��dx�e6�F~�Y]���=j�X��s�N�1�UFi)��[��Ϥ�/����/˴�e���^��*7�H�L�H��=��c�K��!�N�g���je{X�q�
�^T]�B��%��δ�M����P��� ��7C��"�pm	�*2E�b��x9�0-�Grj����I�������6�������
|=I��B�z9�8U�������hl���A��NR7{��(<'�"7�)O}\əev�����J"��+��w�<�e�x�q�Knw�jt<kF�i�T�4I���%��YA�$pU+��x[ח+��nZ^�b�"Е�q��A��b���"9a	Yb��[����[�ۑ �C� ���K��4mn�6[���.߽:�$�@/ޓ����"&�F���0Rr=ͮ%��m���u��S�K$!aV�&*z�)���>j��>����D��_m����7�n�P�����ٳ��$h��4�z����5-Μ%Ȍ$+�e�,���PZ�6�m�D��
u��H7!rąܾ%�N���#s6Φ�bX���zx���OR�ϫ'�
���|�U�z�s3赔Z����o�)DQ���l��ܨ�*b��%�P��/h�f�[7l"ω��@t%}�k~��!(Ё����^ZP�ۊےB�B-3;/�Л'��I�t����&�u��R��VC�	�O�(�@Tf�j��)�/$��b=5c�1��|m,|�<�~#�qE�B�3�
t��̧���	{�gʗv��Uo
��u���1榉o����G�<.g�k��h����Q:�&$���s�y��l&�'#������މ%�Pc6V��晾%UJ!a�� �1�ܥ�[�����[��w7�Ѐ�3Gn�~WC�*�ea��/��R�]_��F���<�2���[p�"���p��%6����R�xJ'��+ś��b�?�I몄�~��m�ŗ5NB,�փ&�4�lG����ѩ�� ��6�6Mpw��߯g�" �~��΋����Z��)��}��;��ѵ�t]l�A��*'{�n `�.�k�����RA_ĥi�$�x�AM��E��	�����R�Fc��;���L�<J��@�Z_T��Ѝ��ݱ�5_��������l��R�&���?��n�&53����|C�2���� �F�pB[ǐ�"6BZ�h��y���z��H;��3d����>&���y���ԡB	�4�e�LI�5��9$?gj�=ڢ����� �.�o�����q؇OQ��UN�*�z)�_-�	(�u�<������C���|A�P�fs�Tз�����__�#)g�*��F����[7�lg�0��3�bS �M�J�T�i�n+�0��)~��$ݣB�^I1�d+�^��!N�m��/���W�8+��\nO���g
V��4O�G�Ǖ�$��T��`�6z=��8���$�;D��0I�E�H4����h�x)�g`W��Q{�����F �*aE`O.@ !�Ũ{ ����e}h_Ŷ ��8ܾ�����n��k��>��P�Ѽ�3���|�m���;tFV38.�0hLt���_�������_{���c�Mnuo�4hj�/�ڡ p�p�(�y�G� y���3@�q�����`�4p����	����[�����M��5	9��禶����74�Z�ꈓ9�8��7#�x�h%�L�d�䥐@��\��)N˦��cc���!C�K"�j#�\iS��A�w�����x���O���O0�r���
>k���;
�l7�
l�0~H�Yhn�:c睋�0�!��I|5[��GR��f�^���vd��X���C��p�$Z8+��\���9:��h�I�ő� ��p�e��X��ZS8�&��K���������	]�`W�������|�ΨԶ��0���x�4�8����Y8�9q5OM)��R���.D=�{ڍ�{��%�l������&��0qc{�K����p1��ǃh%=��RR�!��|�/X�b�e?�K�.,p����|�j/�p��syS�3�<��ꕾL�+���6�vQ�&��h> ~�t�;��MM&��3���bQ��5��e���#� 砲������t5�T��\ks?2��H�� Q��oa����"+���q�7	>	���R,&��0W����^�<��%ó�΍��W�X `]��j5
� �_����>����Z�6Īc������Nq%{;
�p���<ġ$Cf�EkG�04��:��B�~f��Lc���:�	Y�dF0H�����5�k�&��I��P���Ƈ��1�<�/b����>]�q5��:�n���}n��H�� %�T�[�i���x�aZ��&�]�^�ڟ� ���S7�"dd=��ŞZ��A�KagN�Q�%���۵�һ���P�9�5KB�����#�����c���;��yH����/���)�s�0CIF�pI�$���w
G�E�:�3�.�����R��F���|�s0���;�6�����eS���Yqyp�X���%�ሸ}Ў��N ?��%ձr
��Q��g8�D q�����1��ܽ�1���bisr���L��3�soܯ�ȽL��W���ѧ�F���O���N1�W��u|�d����B3I��6�K�M6��fi��V����D����ڬߓn��#���"��
�GP�	�<]�h�r�U�+f����Ԗ+n��7��\
x2p_��L��]��[/��{��Ų�6F��m]�t�Ʌ�]4��M��0�Lwi#�_;�ϫ ��Eb�}�

�(�(�@���b1�D��ʧ�E�a	s�Wӝc�	:��n|�\Ov�\�+����N�L��-�zŪof?#Y{;���U��o�M�P=�G(�d�j/&�w�afs���"�x�M{3.=hNym�k���'����`����� � ޝ[����~�~յ�0��>ȳ_�)~�Ϝ��Uq�6�WS�~�ܙ�q���qD�i�n_�j��'MY�+�co��Y�.�����3�B쵝�}�FZ�ìpl�];�ƍ���:�aC�k�P�b�i��5��!͑�s7��,Γ����L �	������t���Z�g�Ipv6�V`7ce�s(��X��f��� V���r�	M>���٥��^���&�Bw�?T|ߓ����2M�}@n��_���)ڄ�T��'�)��\#�Ծ�*�ǹP�������s:f'�v�>����lk�T+����y7�-Ҿ�񵢓OU��mRE"�`�e�oyJ�f'�V���抾�S�]9 �A����� XG�T��A]�t�x��r�o��\�������h�r�Py�".��f�ﱥ����єr��)�G<Od n�}v8���R3�=�c���"��k�/O�@��ޡ���" ����A|C�yWF˨ّk$�����2R��T#4���_��o+��n}|�N{R&�(*�*D��k�-S�i8�������0%_�YHd#$��Q�ޜ�����w�]��L8��5?�k�&���������AƏ�B&��O��f��'g�U��t�x�^J@_����y��UA��U�'�ˆa��mEJ'L�"�������,L]��B��i�뇖4Ǥ��Z��K�B�h�����4Ai�v���"{j�I��4��G�� 5��1�V�u�6��:�>�3�_�)�.Bz��{�4�QHq(��Yg|ujDA'��Gn����K�|j�Uj����������]��Z)U(�hm�1L���p�i>t2Q��s�i�IE��rq����ꝟ�Y�6�I�;�C]���1�s�.>˪��/��� ��:I��#�WR��ٙ&76Z����Ԥ)9����~?{A��w������c�}o��cf�Mk���\�c߱%�lR��!E����3A2嫩��{Z� �'&6=�O%�����M�Y_�{:F�}݉�E�4���0�^i ��"c����M��?�"�ifq��g�F�!����'ٟ��z[>������T��3��?A$z��M��]r�ve��i��:���b|���M@��Y�E,
л�t���]ن�6�����C�?Ec�R�!��}}y��x.��̇�]7��ޤ�l�y��JW�+��+����&ߕ@v�ݝ{�W�FB�;�sv�:V7"!N�I	�)qV�h����|WXX ���YE�W�tr�Pr��K�p~4j��CY�b�z���[�Z��l:�T��Vr |L>�� �&��v���W4������ �NP�����SxH���7���� �0K��Ϙ*��v03-7^������L�*"N�b�"�<��	�3�:c3P?@���ޚ������V%\���X[UY6f��R�]O��u��������Ϥ���_�㗒~rO�R�Ӳ 3�頬F�B_SdGi�?�k%5�4ww�ƿ�S�r�P���I��9�}�P3��LP�t�K!�RZ{,K�iQG�=Z���çe��wE�Oy���Q�_4�o��k�RR��&n`;��a����>���nTB�Z���+���p�I�.>z��� �����-8�� %ZdCf���4lcs]����<FNDX ԏ�
}�@�&��9��3���&��P�\c`������~"���<�|d���"8Pb�f�Չ�Xhc�z�֙*�~����U*�	 {/�lI���=eo7��&H���	@v�f�>F�i��T��GҐٮJv�i+�u����*��,�l:�����Ep9\de�p�� ��g����	L$��X��������;-8��ԡ��9��M��` [�;P��y�|7y܉����o��E� .N
2��C[Q���x[F
����]��[w�3�nw�c���-X����͉%�1���1�F�m��9�����t(�$F5������̅���ʿh/N�w�vm�R%p� ��0�mk�Le��j�T)'�i����qуl�Sշ�,�h��G��W�_=�N���FTt����tA�@�,k}�!������ivT���bi�$��/&u���aI�m�Tu�����(��y���6J���gNu��۬��@����'�*�D�?����.��6��[N�B+yT�/u�\nռ:a¨N��YodKI�H,����N�����E!.[�o9Z��ݳ�b�<`+`[Wp��*{O:l���B�9��Ƚ,�{��kiv�g�jc��K�\�2�Yi!&\e��~M�i���~ߡ��pgf���.%]XE�n����l1kOL7{,V3J^�~l9�b�1�S�|���u�ʼ~��Ҭ�c��>���58���11+�. @M���nq`id���5I��ń��?�.v��J����\�V�w��6L�r���A7"�v����L�Z;�I�.�u��>pI���f��d���$��SB �=~��x�Fh��47��$رe��&�/��x� ���&��	�HUy��(�q���FV����L�_���7U.k�nmʶyQB�%�Eu�E��Q��Y&y�Kx3$�U+�6@}~QH��Ywf[�nbN:��W���5�"����+#N8S�r+��s�h�1w�{�xZ�� ����>T�GZ۩\*|-pOE��;��<�ʲ��:�m{��o9Q�	E�&�m�:P���t��[�'�T�f�5<JT�����%5q*z���uU2�H�Κl�$ԙ2��1,-@�\i�^�q�\�U��q��Sb�-��m�:����w�w��ip��V��#�,��m���(]#�4�\m(�es1x�uD(w�[����t&��y|��W��`�ks!t,�jE���KYشj��h )��9�a�0��՗������?����Z�'롑��7��3l�q�$��_��5]�� 3Ÿ�h> @���O.~��+m�tS%:@z#����]�.:��	��yM��tX|I&)��RÄ@]���LP�;��@�5�������&�^h�ZN��v`���i{�ՕY5�8bo�+p�Z��MW��ᙞAޛY�h�D�GO��~+���槵��{n(�Z��Oӗ/Hs��=D���l S.˘�~��� ���7���k�>^�3}��M0kvZ.W%�g%^�K+�b8:m
���)��*�s���D���^o}���������X7�2�tq��qz���-~��J��)t>��"���ޓ)��s��AR�&bmBe���zA[��t��{�"s��{	1������U�b��c)&$Fwy����t��n��zխ�>�(N��ͤT85�c��zSSޕ6�i=�=G��h����/P
(ߴ��Ӧ� ����	ܑi�����#y�ƂK��
���zʎ��T�5���,���-�"IBl��Jġ."e�jȩdw��6I�O����(�}�7�;BM�(�;Q~>�� �b#9���{b
�6_#+RE͙hA!~Uy���{7;�X;v~����` N�sKY+}ٹ�֌"�3�-�@�z�޽ė[� S}H�2�\4�B��Z�4=gL�3_�Wv�Y[��M�L�ta���/F�:��ʻ�&u.Ĉ/��ZC�R�G�JŜ�P���.:>x=Q��-�S�蠮iyP��A��`�U��<4��c�є�/��� tמVq�*X��χ��DAM��[6�Q��~��&�0=��s�V~�2R��P��{�8���'����fk��Ê(��\���Q�B�7.RJQ�c���E��x֡��fK��9ϒ�0DѸ���Ϋx� ,ɦ���J�/c���Iō�hW7��P�W� � pcꂀwm�2��q��z ��Bu��!uێ���s��ݮ�͖�c��٭���۶ Z��U�|^g���չ�Ns�Gg��v߭��eH����I�>W�.�G�+��EcL����c��mo{�^�� \
4�1!614?�\f�	�����5b�� ��������_g}�N~h�?��Q�]����S{�H�c-�<yR�����b;�c\�����nl�nK���w�LE$��	���| �}_��.�Lx:)����6�^��͈F�gc��.{,)Nk�׫$�4D�YA�ŭpyY�"!D&�'�#�%�����]�$���������vՐ��C�<y� H�#^���B��05��e��N�M�ɇIaK�
���<��g}�0�민!3��m��
�n˹Q�6�s�nC�BEʚƭ�~X��Ou�u�O�G�o��;��jѤ�̬3b��:��H2>�v���Θv
�[���{�rC��T���X��t1�`��Qz�L��S<��������ka���G���1K� ������+�����`&���ef�:��6��,+�� ��O��a��(wEy��3s��F.7T�C�GH:����8r�n�:�8�H%'8HΌT�K)g��>�;���nQSX����^\��԰9|�̢�b� �@.�5�:��%ߏK�޹�C��7���	C��>�����+R��bPX,�۝�,#�2�����v�����A�>4��|��nBlW���h�c�-B*U��?�L80�����F��w�
X>s��k(+~�-^�� @!gA��I(<y8J�X���'�S�T��CUf����=�/�+��t�>9�_yβ�O�jW�|^���'\����ұ��b���]��u�$OML��9�!�̭���h�Op8y��R̿l�0����UqU��D�,*�UH~{�� ��Yb|5�E?�a���[H��=<,�f�q,s����t>�u��K�æ��c��G���c�L��l
��g��6f!�2�b$.Մ8�qLJ���~3y7�,�\��f,"���8`v��"S�@�ҚY�÷41x�o�a�c�w�C[&�=9FU��ZӞTF�}ؙ�� �9<�����I�)i����\�������t���u�oA	��'�*���{1v$^/�B�Ђsq�V�P��������$�$ы@Z���u�!�Gj�sy_�{���FI�O�������� ��"��M2Q<�a����c�?O/&�2OA�u�p�/��	ݣ<Sà����^'<�iN���!���/�䟁i-X��j��\c�����Rѱ�+�@\}����Q o����[�HA�*=>Mɀ� ����<	����ꌮ�wP�R��pW7�.��@���f"�\��o��-VʠAJ,G�����OQ�)�\��"�IY?���:�R�mnq]�� ���|����
�ۻ �!B��^��i�\�a;N�~�L(n�^b7�#�}06������7�ԭ�[�&z�Az�r+jY���f��tS��L5֘E����Znrf����.�FB'��\��=���T�>D�y��݅��p�R#�a�߉�?�K�Svl�
�%�\[<��hB���ז%}ŒhK�8'	�Q��/C��[]�
~���ja���a>���i�#�T�)����=�h�D��l+�b:�� �y�3�\�|U��*���r���҄�������(������~wD�[+�R�dS��c�\k�9[i�-�0�������h��E�x�l���q>��+}|�Y(rS��g�j�,�*v %ei�jgn��xq�B�����~����隮P�}`���
�9�1NF�!�	���!�0����T���jR�:G9��`>+q���PO��=N����>>�&�V?��{0�V���/�ŝ<���}��AM��]W�yEZ�"�����>�Kf�Ē]u��C ���s�["_ّ�-)�X�r���Y�d�`����4�4��M�σ��P�ⓓ�Q���AB��`/w��I���q��'\���b���c߷�s��n�1+�1��v]U�7MJ�A�bx��?�,H����0=���uq>A��q����n"T���2!�ǔ���L�.��i�D�7@�j�4��ѯ>�<��;��mI:����2��= '���������h�,X���
�~��K�6L�p�~eu�K��E�@<��"�RQIֆ�_N+Ғ��ʩ�	@"��z�^�ԭ�_å*!O�"�M��r2�J�rq�c���*g&Ga5�0bd�"�n{��>����zK���r�{q_�g���VS@љ5��hQ���Н�*�`X�g;k�Hg'<�(�e�I(�1�q�e��ZU�ȶzݎTi�Kv
 ��w Y�O�䅖��l���Cm��Mȍ�:��S��\_�N.�f~S�վ4�b��A�/����F+ot�����8{3C�D7��Q�:�6�D�jM<����PL���g�YWK��-#:f.�\�Y>�s�g�l��y�}���,=�,f�+9�:)��_�E�8@V��U�G�s���=��>{b�8�Vt��Θ�z��O.���o��}���A�Á{,[�.+����;��ؓ��ZG�hp]I%P簨Zr4�l�r}�{sr<��eJ��S�Iq6�F�氁㟗�>{�c���2���;?m�*\�t���E���/��mOj#��+}i-���������0�]S�ozOuч}��O%��D�iKi��留���v���t�]�$��xIN�cnO��h�QO갑�p��K6����nKYEd�ڈ�l�O��L�Џi�جuk@Y���C)�����kpn�PXȾ[�qK$zs�����>��ѧ�ުCcUj΋	>_Q1�����;Q�Y�qS-湲&~����Mv�ә����,�X����%=�g�Zc1}�
�d-��R��`T�f�W����H�,���+&w��&�&�Sݬ=���lZ�_1VJsj�#�����X�<��Yψ(���%���3m(e�'���d�@,:�+�c��Q�>��	�p�hh�>�j��B����=�Br�bfc���	2y�E`?�N��H�q���-��ԃ��ŷl{s$�]�{��|�*��h�����+<���Q'3�}C�lSa�*Q��r˟����Q���N G�pp�-��� <.���^���}�h|/?\�i[���Eg��zyӮqV���ZsR͏"�C�Aش���x;V�oȬ)����
�;��{8��m��2��TC��r��o\V����#��G?���2�A24�/hrkf(�V����&/f������TL#_��7R����&Rޙ [�_�,�)n9�9!f��ui�&��L� ����"�a����fnkA��2/_K��qZ^цj��. �r���V,��h��N��ύ����p�p �a�iς�`�ʃ�$3�<�&�/[�o��<-�҇A'8�?�m/� �י@B��gm˔O)}6��\�/Y�J�*8m=~ZI�t/z�T��*k�~~B_2^CQP��9I��Ϯ~��������	t6��p�U%KW]�1x�>�(�2�NWȲt�Ip �G#Kq�!�M�G�Z���x���eN�F7�~o�)�p���S�=+��d�-���jÀQ�(G��ƫ�w��a����y	�
���z�!|�j��l���h���Ŗ���z���x��`T�����F��q�dݍ����TB"3���?�&�'z����u�]�ѝ�`�5�����^�
&EZ]�p�[�j�-����:����Z�K�cP�5�jd�Y�'u;�و�ܱd�?���d���8L�3L<9B�Yg~���><��{�������f؜�Vb�����*)�3����d<��֘ix��r�-$M��j�2��H�I����M�x�C���69��H�n���b�Y����Kd�B(u�Rb�3�٥������=�6b[h���Z5�1$�)EQ:�m髣00��TɁ��ٗ��p����s��bt�@������"g�<<QDx��+K��C��Q5�Ln�:�涺U���kU��Fs�s/��dN8C'��E���Z����A��$t���� �o/��a�]<1jl��?Ǵ�p�?����6����������{|Ln)�}��cl�|ke�31�KbM��s��6g���o�B�F��������~Y�j���5 )�ߛ7Q��S̗�R����PL�6"皾�&{qg��A�s�L@.Ȩ�z��FMlD����.Q���V�_�ɦt�c*�!���ӫA�$��� �>��N�u�ʑ<��.��)�,%�����U�I#����i/��Ҍppzw������X�ę��"�vbh��xFg����pj"L���~��d�rS7�L�C����w�Z��hՆ�V;p$Js�EȒ��ز��tS��ع�Y���^F��� �e�U���U��֎V۝���,M�4�� �T�rj9��V�vl�zz=��t��k#�eȂ3fN���Д@�B��+:cB�6N�9��)F+�u�[d�p��
WE.�D@����1��>��q�q�ϊ��T����ݸ!Xu�I�r��_�K筻�޻����{�`��'Q�r���!�ԗx;�@��Q�\�:�&�}Z=�X]�MS��Y�к�k�z96�b-��s��������H	�uQ����xs�0a��|��t�P�d2�R����Qz�۬SZ"���\|Nv_G��.��r�>��C�[���Q+�T=�#�^�r�]��X�˓�,���{w�f<߅'�ʺ��7���P�tJ�vɽ$�pA��)Nd�0@���w�l7��Z+,\�H�L�3�ڿ(��s�s���f�cg�Qu�|~�YWH��;��)����a�0u?��P�a�hfTG)�7��I�:�2z�D+Y;$f�����o�=>;���������X����=�f�fiF���Cii~)����;5s�Ҙ	������G:?Jx}�_�ׂ�O���������a�ҥ��e�5U��.w������L����\ϕ���!���1�(���y'o�[$��[�6�"�a-|����<�"�a�%d�)���N*es~*�ֶZ+���@�q�mL�:=}��{��*��##�r.�<�y���W	���'�q�,���s��;@|l4���Υ�\�͖�z�E�u��+ "��՝1�3�I��J�
��!cܚ�������f�v���nbsV�"q�;��v.�]��x���Lh��F(�� ���K����!ߐ�7�\������t%���{Ғ��4�b�5���8/��T���j���ז�*5}h�C�	i�Պ�;�/���j:�<����m7�ְI^|K��q`h7�M��!ȱs��2����>T���Z���=^
�'������`� �/�y�����Nń^�������@+R~WR
�H�n�sY�lv{��H���l�����'�E����d���.K��(��=�]���Fl�a��9s� ~l.D��=<���uӘ=��l�ԯf��\DHHe�G�&�M�jڮ�Yco=�a��OLݺ}JHFW�mq�'ϰ�%Ս�oT�Hii���2:!�ߖO��X{}�7Xbd�\��~���A �K��@?l��蛱��!�&�D�	���,��Ǔ䥵9��>ԃ+�o��2?[���ݼ�(��:���$�2�<o-;�81qM��~�����ӗ���k��H\9��^�c��pU�J�Η�X��[��T�^�ؗ�}��=��L�����0 1�_��*�T6����)��`	����+K��u�Ar���������A�1����A,E��F
�^��x̳ȷ�Ȳ'���D��N�Ϗ%����(��4P��aV:����3�����Q�f ��Ta�t9Ao��t"GYO�\���%Ũ7�3�<�.��A/�7@6��ZS@t���0�X8��ڇ�bH��)���zۂ�Ř;ؗ����+��t�-lS�`9q�yiI+��o�&\�*��9d!�gx8�\B�΍�����(�~5���<>^��P���-v_9�����9�w�^g&��S{i�|�G͎��V���kk:č#�7���3%�W�iyQ�|�f��7�x�����SQ<��&��A���ͬ04mu��I����U��y�%g��e^<�')��m���IP7_�t`���"�?
����!]�[�h�/z�'H���9�k�*�+�R�N}��ΙРh��z���C�m�?U��1�pJ�|��Ψ&���y<�O 搘�W�C��*��Ԣ��R�
�[�9Luf��f5Ѻ�g�A�����cB�(B9f��/���Y%����FL��tP����I�Sd'`zb�F�)�ѽ��x��e-s��^]��֫�a㲡'��R��AS�s�$��o��o��U^ZǴo%����h2�%:�7�}��|�eټ�N!��v0�����+�Q�7 �}�zٸ�[��'q��"]��۾Nk��^����F�uX�>�Zo�3-����f;_f�d�/�K�.��=hf���,�!Bh��tW�]�PW]�p�C���u-�_`�s����x�0]c�����ގ��s�&C�zBp��(�Ȧ�4�4�M����x 
M(U�r[����֊��?5���t���l"OO���_��%��k�����~�h��v)�2$��\*!���,��Ŷ!{��sH{3㤎�������j�'�{�<��@Aũ� ��>`�lȽV"`"ޘ�����?F��A����P ��)6�ئ�FN�(�JM
�ӎ�3W� [x|�iegv����.nw�$�=$!TH����1�P���̛t9z���Z�{$�?5sӀ��Z{�Rm�k9c��f>Q�_��I��`�� �U	Չx�H�=fH�,���kFJt�G()%ڟ�Y|#-҆M�1�.�I PQ"h%G��H���OSA	%5(�L���w����ؓc�2II,��d�)(�,�c�-�me���d���_b�(T6�ED�Ȍ>�T	�i�B��D4�d�������B�j��X&��C[F���xs����&�ߖ����a?�T�������	�H����3x����&��5ؓ�1�
��b]����"汻���o��w�t���#C�^d%�N��bl�9Y�@���:T釫o�FC3P�+�J��9e_�=QT(�$Զ�:­_��5x�t:Ƶ*��YN�[��EH�*MPI����k�g��}m؅�[w*(޻4[���T셕���\��n3 �u\��y[~b"5ɘW�N�/���oP��6�'ŢH�$0�j8b�����T����UW
)�%�z�d�h�\�G�uC�Rv�����
�$�@L��E���\1#�n�侐'��dǓ�ș/xRz�S��<�u7�ܫ&��.u	#ʾc} )F/g����O��7�;��V�=3>�p'�:4������퇠�����q�)�ۊ�?��I�l�_�jv����4Ȯ�Щ��t���nؖ��6g )�7=��B��*џ�k�TܨP��eMS���£~r��=��k~�=�jM���3�Wj��G�9�uos �������/��Թ3���:c�_>>Q���Oh |��\�Jq��8æ魎wn���Z���L��e���{@��=��M����5���ie�,@�D�oc~Q��W��\���vU]Yh��gF�	V�|�m��X�i��%.�ee�OE�3Xp���~Dc��n�@����i}~�z)��J�_��{Y$��)�R_�{-��q碌O�RDP:�l�������?287+��~K�
'h�DV��X�X� U���>e�1ڌy��N�T?F**�q[�d�1l�=�rzj!J�P0�Sib��?�0�e�0RF��y���g ������5��x��u���
7}
�yդ�,���$&uB��Y��*��Z��Z�p"-�I�u��^�T�G�ϰ>��ޑ��vڣ(r��E�h]�N�����t�o|gú�<k7
^��f	w�w'e��� :�����W.T���,�fʝ�3�Y+m��M9��Zzj��*�G�,E��+��A�D!����FZ�����<��7�ϋ�86`��)dA��\?0���I�fS
t�.�ed.�y%t����݃>_�sp��|$'����lAK����]�1#<�g��ϸ�bGY��U�^)hT�I��Y���=R�.�C�$)vM7���vu!�f��H��">�&
�KІ>}A�	� 4�Z�*̱����o��5��	Эl���� ��y��^�S:�+=D?w��eTAí���ڎ�t�2D2iL�%>����� ��4~ƣZ���I3J�0(�C`:���j[�dJ��_�S����8�b�������_���.��_1T�0���~l���a�7�G��1f��M�@�-c:2-!��uJ+��]y�;Aj��a��̅�ưB�'V���6�N_�C�u�A:ɥ[�b�X�B�9-z� z� W���.qO�d��*^��<�S�O�t�F8���
�6y��;�]�ۏM�j�_#t�������O��k-����j��'W'�ܟ��(&Չ�����9w�0E��cѴ4\j��|����~U.��&�9<}l%��F"�,��J�K48ܶ���6�~�sG0�~i.�p�)	izX�tQ��y��_�;A	q
���e� &zê+V�C�<��߷b�����-�GA(���W��-6���s�H���e���� ��	���+��,8� Ź���%P���/_�l�{A����������:(y��1v.�B+=�Hm�'C�z2��(m��e;��"+ e���ȭ�94�,w���4�۲�0	-����-�{X.s>���_��]U��&�l\�\�5�us�&�Ι����C��E�`�I��=���e��"l���I��Ѐ9�n�X		l���.�4�I�-ഽ��j'�U��ڗ�_��YB�fH _/,X�|�P�P����Yͳ�[��/'rN���#����|iD�	�q&��a\��l{����H��8������>(d0��3�~�K�Vo��=%��n��N���� T��`~-���osZ`$��ҥ�h�/�����'ku��<�����`-+�G��P5�	��]�LM�Μi�3z4ː���/I�o�N��J|w��=];[j�����p�M���K[�;m�J@���*��,�����Ct�R�R����:e�Ƌ�i\۶r����ZE�C�|��ѳ���[��h�]�/10�i�qiC֨�v���j��jAӒ~s:O��+x}�)���T7�v�a��y���	�p}��Ѷk6�ę�N��ņQ��M�L9,^]r�b������.	`�^���q�#��6ND�����i[�9�n����ȤP2�<�;��VH�@Z'>R#}4L�+l��N�!������q����yqD�� ÏyN}dkY��"b@���ͅ��e|�p�ږ��U�w��#�0�%��������v	{�"~��̶3�n�j�M�����[��R�H4��p�A7Q�9@&���i����"���A�O�P�}���x8��=���N<�*�6/PdѸȵ�i����V	�V��.��bK�"�ȑ9znN�l���hvnb�6ށW�J�3��������UI�[�F��>Iu�=Y`��F�H�J5�>v.���ˊKO�g��'�����5��u��Ayޱ�W��r~��oMᚼcv���,���� �^n�:? /т5���HE�W�\AA��)Ќ�o4PO���#�Dil�d��k�5j;��1��챺ʬ���.p��״��}���:m����p�7�p��{�o���;����Ҝ�jN&\sHh��K���\HgK�X�R�鲈M�H��d�E��$5S�����=�!k�NOn�H���䅾pp�A*O�o�KHUN��2�bE:�hm���]�fv���_�s����j�C-EM�k�#	���Ȼ�o����];h<����3m�,v}�1�/m�A������z����T��ϸ}�3c50�R\k8mb� ��T�H7��P�#�l�Ʊ#��n������-�XDa�(o�$�~�����ى;�uK�0#%,�k���A���cʐĜ�[ ���}/j}��T���R �	j{rc��M��$�&TL���5 �m�G@����yqT���e%��GmO<�GqN�����;RN"�@P�6Ǌ�� ������Z���B�2o�
u��[�|]:'�j͑���2|�̞%9��P�-�С"��Q���e�4���f�%?j����J�$`)�n�NI1������􃰅�:J�S=wκp.joE�e.v��8��ӊ�̂��+���05�,�}-��H�s݇��+�b+�ϳ�8�?�#����xӺ\<�^�FrT�y
]T�����I���Ze�
q����K4F�K�32��*�zp�͂���+���*���^��_�K_u5������nC�OI�rCLjB�L�b�V�M`{�x�h����A�-�H+d�0��E���K#P��Y}�\�,y����a$��u�������P��;E/�@��
s9$}�v�d�HBv��)�n��n�F�i����A��o�J��_&)zE�������bbj�zabf(��)~m�UR��ޣ���:����� c�
�e ��`ha�^���e�pכ�R��~���Ԅ�a�Hm�s�}��	�����I_G�I��|t��܇6|�:���PK��j���~�!�>l|%�~9�TsqR�ঝ�i�Qo�A��b��.x_��VB}��n�5.6�ڌ�M��٭b�]�����5X.��ܠ;(/N�S�N�l������1�J����:G0�il��3�YY��(B2�ȷ��*=
惃\j#��oQ "vU�֡�j�my�R�B��|�ޝ�	�Pm�8�;�DƊ�Y 9�+H4Ayf��¨8gx13��MS���%+��k�	�8�^�D8��ժ�I>�x-j��>��>�?��`���oɀY+��mC%�G�\S���_d +#82�~��-���vc T#.}�����Q���c
9q���)���<t�=\�׫���F�@/�� ͨO��#�欆�A#��ɭ5w4�,�Q�ۭ�U��	N����^ �b]gJ����˾ѵ�� 9bm���&��*3�B�������]p�o�T�����<<}��-�E��_�5�U�`u�����.wQ
6)��=��l4z��'_�������D�W�œ��}�����@�`{�cb��༿«{d6��8(y��y:��/`kh�͝Q�S���$��U���E�Ɏ%UV�h�n�|-�O�ȳa�s4>�r��*�]fa����"M2c�f�\������-�ʵ�M���g[�%"hgZuW=@���?��������	QV�)��N	��0,r���D �mņ߂p�L2���H�<[Q�p�w�j�n9�+	�Rٗ\�4y���_���;���.lGc8�K,1��Zđ���_lM���apjj�Y(o������:]\�:�E@�+d�W�HX-L=/x��"jk�q�n1�><��(=E0|�f���0=������'��y�ˌ��Z<j21��*�k!�ǟ�r���wt�MA��ڊ� �?g @\BkTqĹg�KV�O>]=TU������Yq,�3O0E�@U��j\w�E�8	:ǐ8tt��0�SS��sd��#�`������[��ߐ|�I����lŝVgjI8ї=@���y�r�+�ē�0�F-S/�L|@���u�u:y.����I@&g��+˜g l������irwI'�5	��D��q�3�.�i?����.�n���p_k�3�ېh��oӱ|��:�W<C�x8�?��hT���/-�J�.��;"����Ħ��ab18	*!�x�.�7�#��5���l��b��s>X��>#��F�l��|C��"0�߱��2��I��G
~i������2׍�đ����{>̑| ���b��Ei���B�=���v	��cPק�!M��A��΋N3�jE����,`�|�NUB?#�[\���=��e
��5XaQ1_�ER�Yޚx�z�eЫ?��oG՜���56�J�T�����ri���jomVa�\#�-�s;@tD�Z�"�S�1����P
I��J�C�o�oC����STQ���.��q��r�J�i��aL�+�&��:�k�K�vj;���P6>y1n�nC��ܾE(62<������y�V7�{%��AĜ$H(`��B�O�����A�L�fO��p���4�N�70��\��)��]g@�%7��S��B�����vJ��b�6ѓ��G�Aݒn�*�8�p��S_%�p�k�&���t�k�N�*P$ h(��~W�EO�������p���Y�/��3uy��G[B��	 ��"qG�}KY����E��-=�P�4��k/�wґK�0k9�f��$�]&/�/o�&�*����0���y�HO��;��{�8k^������1� ���X���S��6v���sK���{�O��@��7]�p���t������`�}�(�AKp������iQT��e�e�Q�uҽ�P8�<������'�X�b,�%��H�O��jp_e���0�����!�{��������������_�,t��7^��|՟m��q�_/h;՚d),�QF��)钦;>ϯW����@��'��Ö����9ڳ����r�ʪR�8�hK���5Y��K��C��a�۪�񗂝g�z1rs�̻�q���`�?W3�V��r^�v��,ld8�=�<�\���6�&��r��}���^+�����,��r)('��z�D�����2<�5����AAE<���mԩsПr�i�UU{[���m��K�9f��$"[׏�l)�4Y�7ZV�?K*3�<ֶ((�|(f��C2��,Yw��VT�r�Һz<u��Q��d~Qdb�\�-��/T6�={1uGH�#b�h���jԌ�(QW�w	o@��Ke3��M��=@ڀc�-)�8��<���G����A�f�<��W��=�e�ܺ��������ѽ�F��?��,�U{�ػ��)�(�^ֳL~�F�u	Ĳ�E�p�U|��bY��c]��z�q�Fm��l,�~�7������
[���UCN����P��� �;�_@�qՔ�O�'���.�6g{�U�Ǎ�lcfm�u=+�͘F����B�꽐 �`ʗ���{��ւ}��
.�ᩊh�Ƙ��hQ񫐖67gg�$dʲfrqؒL�cл�ʸ{C�C�����MmS|p�%��UDt{I?�Y'�3WQ���{�\�~f9j�C%�RY7�c4Y=pT���A �[7�g%g��MS��q��EU��^D���5Z���.�D��SJ���g��L �H�q!n$?�H�G��Y|�Ө�}Si�X?x�()��K�{���^��H�H�\( �l����w��f�(E~��|	s�-�3A�_�W\7���v{>ur�0�z�_�����Z$�i\ڎJ�n�j��	Z��YR��q�w����xQ�Ӗ[��6���Y��0��ݜ��J1�P:��V�ˋv$__^I�r5(�=��� ג�B`:�nu$~��{���x]�ʾ|�n��L{X� 7�{)Gp	O!.C�ߖB�5��?$�qS�V��1� ��\�~,��� �"�=�ֹ�S��jy���Ӫ��_<߈p	����$Ѻa�2:���>���ɶ�� S�u�l�>��V��Oϫ��u��9治|�ߺ�wMĥ��I�K��|���E�~d�7�3\؂���]�����ׅV�Y���W��w�mh��`�F�$��Yˏ�Ҁ6`�������A[��r|�&9�����-�E�\�m)rk���@ �XV���ĲzA��"}��m�q�G��V� ���L��N�ȃd���oh�jG;=����1��T�ڄI,�?�߈���𝂐�^�I^�t���9k�w��^�4��K�f��b�,���^<ٞ�����z��ׂ>���cMQ��W���h�yS���e5�Q-�c�y���=�&.֨Ic~��E��V�n])�&ö�����D֟<ߵ��u�pH�Q`iT�q���U�}��P��5��'E�o
Ŋ6�z,�s�(To��=��ϖ&��J�Ʌ���j���'u