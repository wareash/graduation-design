��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]t���cJ���{t"a���~�������l݋"X����,�~�� A�ɀ��B'�"� g���Q'9Sq���G�u�O��a���>�f/��7��6!Pۈ��b=q@2�J��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��/��Q�w���a5P��B�~�/�'̙���S{���^�qѝz��'�hřD~dVr�F�!5�=��[�\�bYzy��d�(5���*���D#����=�6�c�p�GCE�N��+�xh�Eaa�Ƭ�z�5>��>s(�oƤx]C��F�i�TϚo�2���E���W�۠N	Rw��#fa�E����ǁ'�iM�$r����?�W���aݒ�3��L��'�ފ�q��p��FU����vJ�k�~���l���wFpe [�29��Zq���)Rq�� �CPu�)�;��/�V�2��'cu�*�Q��펊(�Ľ��N��������PDEL��DK�/9pD�P!;��V�P?t�;��ww�3��Ib�`G;��g����� ~�zӋ;��p#/Ǒ%c��U�����% #X���]w���x�Ͷ�׎呮�Pj�������O�*�p�ܝ��@jrQ|B���T(�?������!�묅��2E/��)�@#�O���.�"���E]	O��m!�����Zԟ�'�0��2�-��n�d�E����H.�х@�O�k�V�-�q7�^`��w���lr:Ry�VǞK�#�H�oC]��ǻ���Iu��4��oYЭ����+D_�ټ߃v/hR N�
���8B�ҧy�?50�JTn-U�q�5G��s�4���֙N��(q�B7qH1h� '���� ������k����3C��ݴ�.t�ͱ7F��|d&n�Ñڳ��;��p�]}�+�������z.�);芴�63�,(�gS�vZ+�e�λ@�0����U.�8[�2
����Ԗ���ٹJ\G�G����w^ɒ�×��6gVA��2�)�S���V~�Y��A��<B��/Gy�&�NA�X+�&PB��L��Jd�V�C�5P �]���Y��9�����Q<�f�BU=�1�x�Fc�\��Kp�&8S\l6�H���5~լ}bՏ�,�$u��-����}․\�z�l&�0&FD��縳�Mm��P�&��5s��X�h���l+Ǌ�b�������M�g�)>&�!��2��>X�0�M}������id����	�	D��E36_�/d�8弳�Y�^��iF~��� ?�xv�)����1�T�Vl�8�JkRq.���PR˛����_�%P��n'|w,�$�q�qw#	�{���[���O���pxG�;����-+������+NkA��6yP��V
���3U����H'��k����Ƨ���I8��J�8Fl��Vr.��L������\-��q��IԆ#�� o��72��Z�ݸ.��cG�n�bn�j S�A��AC���5a3��NP<"����ǹ��ؙ��nd����/�G��+_�|;m��ҬE|ҟ�oe��|�F V�\���������'���ΦM��a1�{���n"`���A���ךa�Uy���a	N��7k��J�p6��>�W���&넧I�ن zo'�����2(�Z��u�c9��&���71*P{�tA;��s�H7m)��qY��	��;4�N����v�"^�HT���'S���~��G->�4�L/��V�y?ڍZ��A��Ă��1)@1�4����#�qk��5� ҧ�{]v��P��wS�
�7���\'"��	�S��F�JW}�x��Q8%��39������-�R�
�S���=h��2= �^�ɴ��#k��T�"�|P	6�v	F� d-'���mC,`H}��y��<�jrU���给�e/��r� BM�-rЌ��:�wS2���ٟs����Ԭ0�k��߹���eÊD��dw���/U�N[�̍���ޅ�{<�OTYQ�%Q|7�)�c�M���ѵ��9(|��c�Q��3�Z]�a�σ� z>1e%[�45J��匿
��C��m��~>nT=1���g��r��^�%�;�VVd�?W'��f���?�C��3ު�t���} ��q��گ}{O�8i6y�A�y���1>:q��R�D�Mbs"�c��zh�
���)bJ}���_4��Œ���)�,�Yk���*Ǹ|3/(�A
�a��9�m�WwZ���-�L���u��������~l����L�4D�PɱF���K߂���ʫI~��Y���������J
��ީ}q*,��
!�׭K�5�e��F����8��:�b_�ߊ�rH����fA2�6��H�T �g|�&r�2_5_~Ha�8ܥ��QW\��V)���s�z�:�Jt���pbseFQ-�Fw�s㝤��h�<w�JQ���~)�s��*S�Q!tA�v��4�HD�4l_��O7��k'%�c��nG�60�-���s��0�Z8�6�i���8�(�+@�S��U��+	����vM	�t����JaƩ��#vlw�&wބ�\����	l��xX7K)8C�{])�(�]Q\I����ZޚX\��=XZ�^n�#��5�y��@/����UFL'2����.t��I�cΖ���]T�XR�{�����f�\�����2�+	�G͒2,T�s�O�`�����P�o� �?soyW�9��H7��&��.{vX�jˉi��3P�j,ní{
ԸW̞F�k��kc�
�% ���R!�G�z�]Ʊ��x�:���7ld��`��*�@3y`��g����x�6r�М�l�J��Zp�걦�b��=�g�+�|ˈ��tr�Ζ�L�Ww��B�7	QH;�ۄ�/%��#&KI�z���fpc�;�DP���0��T=ecp�mլ�"-�$�d��4�w����~����/�N��&I3���#籍*?�jʪ���~Bni[Nyp|��4WcV�U�ݱ���ej0���2����Y:�D�u�}|D���oPU�ʘ��s�]ұOD&~�d���rA���5	!��,*��[�j�I�b{�W���P�`�7gE�9�Y>KHa�
>[���=o�)��C�K��E��	��~�p̪W�~�0N�޾9ƶU+U���J�gŜ����KU�a�.E&Q�[�E�����;uu�j��Q�hU�{Kl=�3�y�(QvD���}��0�0�!J:f���<�+p��_��f��W��^��x(���p��`����u�i�J�ud%}E(�&�VK~��f#ߏ�Ӫ��0�F%0���kV��DJ�D��nP[�K�>-q��� ���8-y��|+#�*P�^[��;hK1��*>^�o�Z��[]X,|��᳥xP�C,����� �~#�δ��5yg�v���~#��Pt7����̈́����U�C�Ei�h�T����W��˝����Z��k���9%g�Z��	6��WS9�ݟWB�C6��2Mo=�ٵ^/��5*	����1��u�(2��ֳ
�/�'V�h�}H�o9�Of�j�E�/zV��mm�ދ�X"���z�~I��wuYw�M!Ӌ
dk��jr�沿��2�˪��u�M�
�Po��?,� ��v � �j�ywMM���^�73�~�s��;�u6���`�F�`{v,�.��u���V��L{>���T����� _gF�H|�
�˪|�yOk(�j^�{"2Sq��|�!^�0G|u��(�ȝz$���}�~���o����P��v�nP��9r1��}�7��	ɢ���Dtp�|$�Ӧ��ٹ\���naHȡKS���BgvZ"y#[	R?9���+Y�r�ʦ�����D���eX���]�'6�t���V����N�&���n::�B�1��2��f	,��3�Ws����<���ؑ�mwZ�8{R�ș�av{x��9)+�����4�ټ��B����*s���&A]��*�wK�}~�9��r%V��{X�ɤ�M�s 9�VzD��`^�y/�_thV�(D
�\��Ԏ�F<���ܕH�]g�:�y4��� ����o�������\,���B	k�R��L�QE5�%����M��=�����S���m���Å��)㵹�v3��ӱ�4�oOrս��?�n9h���V>��r*<I��� F�		]���'N�e�)1��X0��e�)���Q��ƹ~�� �(/�y3�ּg]L�m������3���Vp���$
�H�<�qFdY��B��\�	ځ��{�.��4F�8��Okr"��0A�Ҁ!SEĸkwXr�N0U]˙��/�����K��

�0�N:�[Px��VWw����8X���5�8X(2(:��J&-f-�]Oद~���9X#y�g�U���k:��}�+�ͬ�z���)�#͸�J!e�./���Ǥl(�?���6;��p,d�7�X�Ed�N�c&i��^��V(j�v����p�O��q�k22��g�y�k1�}�-����X.�*�z�
{Ź�T���<)��-�dR)=����Ed�d�-�d-��|����$c�l�e���Q����̐����h]}hiE�W3ؘ 9�A*Y�6b��8���]��^/L<����/��\WYks�k"���A���x�rX;hvڃ��]i�T�;M?ϣ��+�˫K)���BT�!L)��#5 Dy���$ �6ڐ$ޡ*��d�T,"�@+���/ &PkQ��ՂMx�x����b�1NiA�\�c�U��R߻'j�rD7,�a�P�*��}����R�maaCw�c��'H���-w��3M+��ј-�D��>�*0PU!��nֲ�Ԍ�NqhSj]M�/J[@/�ԑ����}<Y���fȗq�뉪li���z�r�Ac����d�r�\m�G����?�0(������Ҧ���6j���E,�t��������oɥ$��o�TҀO��Q�|� �w���G:ʫk���ȓ8'a�*mVP���k�gRpK�tt�9�ݐYb0,5sƚ$�x�ʊ��c�SQ�,���G���

�d�ޤIHo�<_��9U��N>����$bl8����5 X/-q�{���^˖l��\+�[N道��#��C�"�㒵T �sQh
�E��t��b��������#�߽	�XP�-���st�M�eȢw~�?�����h7�Hۯ^�Q}�������$�8�|j�%r��@�C�e�T�&��l�+ΝX�8�h���oCmJ};�딿06��e�|�b�ed��C=�	��g��p̔��JV@/gA�"��:�-M0�r������9�Y,���/Ȝ�b5t��k�(�N!�2��k�$�L~p;_^����Hܻ,��Za=,����|������{fv�|i�n�V�yp§h��9+є��dȲ���NL*hs,S�w��0�qk:��D2t�ї�v��i�O�x�|��L<9�:?c�ғ<+Z
CY�5��(�I�đ��y�8�m�k�Y�Ѓ�f��=b�2N�!Z(P�=�SjZKe,�=�x��R�-Gҏ�����~���U���|K�Z��Դ� ���b�L<��=֦�|\�dL_�����o���a���#d܇������)����:V���d��'�JN߫L�F�%��CV�us՞����0;^����&�m�13�V�M�=�L� �:M���9[��H}�Z>c}.���+oeV��ĩN��4*���@��~7u��Q�n`�Q��|x�pu]��2�[xb�65D&W��Z�����4�;Y�>ʄ�d��w`��6�X�z1�O�J�d�?���.��c��_��ۧL��]Q4�4D�ཏ��:Jx�x���E�B��oux�}����xY�����Ձ.b�W$���F���M�؛�-�����	�7���^� �g�^q�4R��� �?���b}9>pEv"G_��������B#Q�-�K��O�y�w�������D��0J����N>��;����1�GvA�kv��ĉ���`��f���`U�S+���������Q�2���kRK^P�������"|��-]���U��ԋM8KH<�U���Ѡ����T���h�����uTʝ���ྛ>�8����r��M$tT��F�p�b���P6�js��_|-��F����ھ���AAŵ�����;�t�x�2���"T��jٴ[�����@��8����p;	�@�D��/V��5c��P�����5�1��vt��8i\�-����R�
��"��Q>���4������Ҿ�7-/W��;$<Sƾv���>��B�����F�t��l��䦸;,3��MD�zGAy�i�9�c#_"�p��\�"���L�s��m��#�4�
����좬G����������4��,F�{�����a�Yt�x>���O�1b,ҹR����)#��э"k�w�tUsG�먮��/�41��1�c��JqξG�2/�B.�z��b�Wl�����l�K^�H>��yZ�
{����9�2y�vm�Kg�����4�x.Dld
��I;���up�����^�]u�$/�ф?�3�g�H�|+w��n�?:H]����C
B0���	��_�!4᜚��$:ʿ�j�g(>����wW/�#��{���d�x)_s�9���<hh�g踈s�|R����70Ux6�8�\/L�
q)X�
0����%���a\凲�'}60$�уx+�����|Ih��i�u����/�hӚ�;O���wLjX �n"ؚ���gq��'ū�s��>�XR+˼2�����;�|O)�e#�j��45�Y��]�Y}ń��PV�9a���W�:m��5�r*�-"�.����{�-vA�Y�.�N�y�Q:Tٶ%�Zl46d7R��b6$P�1Ŕ�VZH�!1d��B+�V�"���],
��=�(�
�Q)}+J��~o�D-�v��0ft�U���uY���&.���w��ck\!����ß�
������1�x�9��N��@�kJ��Qw�R�Vf�B�`��{��¯ ~u�!�t��P^���DZ�i|���K���*�d�k(�?��2S��=1I;ҏ^y�;dB>b~�+,Ä�h";����� ts���c��kc��v>is�S�S��F����Ꮑ�a��r�bGN�Z�+��L�!��`5?T�D���t��p�ky��D_�O`�d�5_���s��,�������/!����ڔQPH�Y��Xt}e����/�{eخf'e(M��w&��)�o����B��!He���[-V��opz��Q6N�z�~�^�R$o�s����GC �DFR&����L�ɇ��t��@�ǃK�}���<8 r���`�'V�f�gҭ@�q��&�1ZWZh�9b"�	�O�.h!+ /&B>ZQb�� 9=i���~�\��$��Z]�Z��>|a��h�M۳<���{5Bl���dN?h^w�2̪�����0���
|� �<P��{s�(�i�~U+6��߹�8g�V��f2,���\�Q��6��';���4�C(ؽG�kl'ޖ�wP�_��W�w#��9J�0��4�+�)J�!a�>�ԅ	�g�����0b��RT/?Mfe��iJ���n7X,]������K��ş؋>��D)��D�zK�?L����2Kx��J!ef�i��ޜyVi{��J+�%7����0�S;��3b�&ǪhoŐ�����V���%��?��#��E�a��|aّ�n`+���7�^_�S$��"�f�T�>[y`�bqWH�'ro$�Pq�8T���ASa���!<��D�y�& �h���q����`�/�(��� �u�	&P5�=m���^�=,ADk�+N��0�uL���j\����A�{�������Mz���"?%Q���݋�q�qy]�%dWu�n��(|{b�/gY+����'�~�>Da��p�<�y�#GM�X�n����� ���p�<���P��Ԟ��a}z17�{��*��3a�eVE���ϼ�>G���P�"�Lךހ�t[�I)l it��#h��U©E��$?Y-���X$Nf0��#���Ll��lAS�(R}c�Tvxw��Vr$^���������ЫQ�M>��P��O��+��wy��G�@O)5e�����4-��!>�x����SW�(�